module matrix_mul_10_comb(
  input wire [31:0] TestBlock__A_op0,
  input wire [31:0] TestBlock__A_op1,
  input wire [31:0] TestBlock__A_op2,
  input wire [31:0] TestBlock__A_op3,
  input wire [31:0] TestBlock__A_op4,
  input wire [31:0] TestBlock__A_op5,
  input wire [31:0] TestBlock__A_op6,
  input wire [31:0] TestBlock__A_op7,
  input wire [31:0] TestBlock__A_op8,
  input wire [31:0] TestBlock__A_op9,
  input wire [31:0] TestBlock__A_op10,
  input wire [31:0] TestBlock__A_op11,
  input wire [31:0] TestBlock__A_op12,
  input wire [31:0] TestBlock__A_op13,
  input wire [31:0] TestBlock__A_op14,
  input wire [31:0] TestBlock__A_op15,
  input wire [31:0] TestBlock__A_op16,
  input wire [31:0] TestBlock__A_op17,
  input wire [31:0] TestBlock__A_op18,
  input wire [31:0] TestBlock__A_op19,
  input wire [31:0] TestBlock__A_op20,
  input wire [31:0] TestBlock__A_op21,
  input wire [31:0] TestBlock__A_op22,
  input wire [31:0] TestBlock__A_op23,
  input wire [31:0] TestBlock__A_op24,
  input wire [31:0] TestBlock__A_op25,
  input wire [31:0] TestBlock__A_op26,
  input wire [31:0] TestBlock__A_op27,
  input wire [31:0] TestBlock__A_op28,
  input wire [31:0] TestBlock__A_op29,
  input wire [31:0] TestBlock__A_op30,
  input wire [31:0] TestBlock__A_op31,
  input wire [31:0] TestBlock__A_op32,
  input wire [31:0] TestBlock__A_op33,
  input wire [31:0] TestBlock__A_op34,
  input wire [31:0] TestBlock__A_op35,
  input wire [31:0] TestBlock__A_op36,
  input wire [31:0] TestBlock__A_op37,
  input wire [31:0] TestBlock__A_op38,
  input wire [31:0] TestBlock__A_op39,
  input wire [31:0] TestBlock__A_op40,
  input wire [31:0] TestBlock__A_op41,
  input wire [31:0] TestBlock__A_op42,
  input wire [31:0] TestBlock__A_op43,
  input wire [31:0] TestBlock__A_op44,
  input wire [31:0] TestBlock__A_op45,
  input wire [31:0] TestBlock__A_op46,
  input wire [31:0] TestBlock__A_op47,
  input wire [31:0] TestBlock__A_op48,
  input wire [31:0] TestBlock__A_op49,
  input wire [31:0] TestBlock__A_op50,
  input wire [31:0] TestBlock__A_op51,
  input wire [31:0] TestBlock__A_op52,
  input wire [31:0] TestBlock__A_op53,
  input wire [31:0] TestBlock__A_op54,
  input wire [31:0] TestBlock__A_op55,
  input wire [31:0] TestBlock__A_op56,
  input wire [31:0] TestBlock__A_op57,
  input wire [31:0] TestBlock__A_op58,
  input wire [31:0] TestBlock__A_op59,
  input wire [31:0] TestBlock__A_op60,
  input wire [31:0] TestBlock__A_op61,
  input wire [31:0] TestBlock__A_op62,
  input wire [31:0] TestBlock__A_op63,
  input wire [31:0] TestBlock__A_op64,
  input wire [31:0] TestBlock__A_op65,
  input wire [31:0] TestBlock__A_op66,
  input wire [31:0] TestBlock__A_op67,
  input wire [31:0] TestBlock__A_op68,
  input wire [31:0] TestBlock__A_op69,
  input wire [31:0] TestBlock__A_op70,
  input wire [31:0] TestBlock__A_op71,
  input wire [31:0] TestBlock__A_op72,
  input wire [31:0] TestBlock__A_op73,
  input wire [31:0] TestBlock__A_op74,
  input wire [31:0] TestBlock__A_op75,
  input wire [31:0] TestBlock__A_op76,
  input wire [31:0] TestBlock__A_op77,
  input wire [31:0] TestBlock__A_op78,
  input wire [31:0] TestBlock__A_op79,
  input wire [31:0] TestBlock__A_op80,
  input wire [31:0] TestBlock__A_op81,
  input wire [31:0] TestBlock__A_op82,
  input wire [31:0] TestBlock__A_op83,
  input wire [31:0] TestBlock__A_op84,
  input wire [31:0] TestBlock__A_op85,
  input wire [31:0] TestBlock__A_op86,
  input wire [31:0] TestBlock__A_op87,
  input wire [31:0] TestBlock__A_op88,
  input wire [31:0] TestBlock__A_op89,
  input wire [31:0] TestBlock__A_op90,
  input wire [31:0] TestBlock__A_op91,
  input wire [31:0] TestBlock__A_op92,
  input wire [31:0] TestBlock__A_op93,
  input wire [31:0] TestBlock__A_op94,
  input wire [31:0] TestBlock__A_op95,
  input wire [31:0] TestBlock__A_op96,
  input wire [31:0] TestBlock__A_op97,
  input wire [31:0] TestBlock__A_op98,
  input wire [31:0] TestBlock__A_op99,
  input wire [31:0] TestBlock__B_op0,
  input wire [31:0] TestBlock__B_op1,
  input wire [31:0] TestBlock__B_op2,
  input wire [31:0] TestBlock__B_op3,
  input wire [31:0] TestBlock__B_op4,
  input wire [31:0] TestBlock__B_op5,
  input wire [31:0] TestBlock__B_op6,
  input wire [31:0] TestBlock__B_op7,
  input wire [31:0] TestBlock__B_op8,
  input wire [31:0] TestBlock__B_op9,
  input wire [31:0] TestBlock__B_op10,
  input wire [31:0] TestBlock__B_op11,
  input wire [31:0] TestBlock__B_op12,
  input wire [31:0] TestBlock__B_op13,
  input wire [31:0] TestBlock__B_op14,
  input wire [31:0] TestBlock__B_op15,
  input wire [31:0] TestBlock__B_op16,
  input wire [31:0] TestBlock__B_op17,
  input wire [31:0] TestBlock__B_op18,
  input wire [31:0] TestBlock__B_op19,
  input wire [31:0] TestBlock__B_op20,
  input wire [31:0] TestBlock__B_op21,
  input wire [31:0] TestBlock__B_op22,
  input wire [31:0] TestBlock__B_op23,
  input wire [31:0] TestBlock__B_op24,
  input wire [31:0] TestBlock__B_op25,
  input wire [31:0] TestBlock__B_op26,
  input wire [31:0] TestBlock__B_op27,
  input wire [31:0] TestBlock__B_op28,
  input wire [31:0] TestBlock__B_op29,
  input wire [31:0] TestBlock__B_op30,
  input wire [31:0] TestBlock__B_op31,
  input wire [31:0] TestBlock__B_op32,
  input wire [31:0] TestBlock__B_op33,
  input wire [31:0] TestBlock__B_op34,
  input wire [31:0] TestBlock__B_op35,
  input wire [31:0] TestBlock__B_op36,
  input wire [31:0] TestBlock__B_op37,
  input wire [31:0] TestBlock__B_op38,
  input wire [31:0] TestBlock__B_op39,
  input wire [31:0] TestBlock__B_op40,
  input wire [31:0] TestBlock__B_op41,
  input wire [31:0] TestBlock__B_op42,
  input wire [31:0] TestBlock__B_op43,
  input wire [31:0] TestBlock__B_op44,
  input wire [31:0] TestBlock__B_op45,
  input wire [31:0] TestBlock__B_op46,
  input wire [31:0] TestBlock__B_op47,
  input wire [31:0] TestBlock__B_op48,
  input wire [31:0] TestBlock__B_op49,
  input wire [31:0] TestBlock__B_op50,
  input wire [31:0] TestBlock__B_op51,
  input wire [31:0] TestBlock__B_op52,
  input wire [31:0] TestBlock__B_op53,
  input wire [31:0] TestBlock__B_op54,
  input wire [31:0] TestBlock__B_op55,
  input wire [31:0] TestBlock__B_op56,
  input wire [31:0] TestBlock__B_op57,
  input wire [31:0] TestBlock__B_op58,
  input wire [31:0] TestBlock__B_op59,
  input wire [31:0] TestBlock__B_op60,
  input wire [31:0] TestBlock__B_op61,
  input wire [31:0] TestBlock__B_op62,
  input wire [31:0] TestBlock__B_op63,
  input wire [31:0] TestBlock__B_op64,
  input wire [31:0] TestBlock__B_op65,
  input wire [31:0] TestBlock__B_op66,
  input wire [31:0] TestBlock__B_op67,
  input wire [31:0] TestBlock__B_op68,
  input wire [31:0] TestBlock__B_op69,
  input wire [31:0] TestBlock__B_op70,
  input wire [31:0] TestBlock__B_op71,
  input wire [31:0] TestBlock__B_op72,
  input wire [31:0] TestBlock__B_op73,
  input wire [31:0] TestBlock__B_op74,
  input wire [31:0] TestBlock__B_op75,
  input wire [31:0] TestBlock__B_op76,
  input wire [31:0] TestBlock__B_op77,
  input wire [31:0] TestBlock__B_op78,
  input wire [31:0] TestBlock__B_op79,
  input wire [31:0] TestBlock__B_op80,
  input wire [31:0] TestBlock__B_op81,
  input wire [31:0] TestBlock__B_op82,
  input wire [31:0] TestBlock__B_op83,
  input wire [31:0] TestBlock__B_op84,
  input wire [31:0] TestBlock__B_op85,
  input wire [31:0] TestBlock__B_op86,
  input wire [31:0] TestBlock__B_op87,
  input wire [31:0] TestBlock__B_op88,
  input wire [31:0] TestBlock__B_op89,
  input wire [31:0] TestBlock__B_op90,
  input wire [31:0] TestBlock__B_op91,
  input wire [31:0] TestBlock__B_op92,
  input wire [31:0] TestBlock__B_op93,
  input wire [31:0] TestBlock__B_op94,
  input wire [31:0] TestBlock__B_op95,
  input wire [31:0] TestBlock__B_op96,
  input wire [31:0] TestBlock__B_op97,
  input wire [31:0] TestBlock__B_op98,
  input wire [31:0] TestBlock__B_op99,
  output wire [3499:0] out
);
  // lint_off SIGNED_TYPE
  // lint_off MULTIPLY
  function automatic [31:0] smul32b_32b_x_32b (input reg [31:0] lhs, input reg [31:0] rhs);
    reg signed [31:0] signed_lhs;
    reg signed [31:0] signed_rhs;
    reg signed [31:0] signed_result;
    begin
      signed_lhs = $signed(lhs);
      signed_rhs = $signed(rhs);
      signed_result = signed_lhs * signed_rhs;
      smul32b_32b_x_32b = $unsigned(signed_result);
    end
  endfunction
  // lint_on MULTIPLY
  // lint_on SIGNED_TYPE
  wire [31:0] literal_70996[10][10];
  assign literal_70996 = '{'{32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000}, '{32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000}, '{32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000}, '{32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000}, '{32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000}, '{32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000}, '{32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000}, '{32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000}, '{32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000}, '{32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000}};
  wire [31:0] literal_70998[10][10];
  assign literal_70998 = '{'{32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000}, '{32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000}, '{32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000}, '{32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000}, '{32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000}, '{32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000}, '{32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000}, '{32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000}, '{32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000}, '{32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000}};
  wire [31:0] literal_72008[10][10];
  assign literal_72008 = '{'{32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000}, '{32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000}, '{32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000}, '{32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000}, '{32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000}, '{32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000}, '{32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000}, '{32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000}, '{32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000}, '{32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000}};
  wire [31:0] literal_70997;
  wire [31:0] literal_70999;
  wire [31:0] array_index_71000[10];
  wire [31:0] literal_71001;
  wire [31:0] array_index_71002[10];
  wire [31:0] literal_71003;
  wire [31:0] array_update_71004[10];
  wire [31:0] array_update_71005[10];
  wire [31:0] array_update_71006[10][10];
  wire [31:0] array_update_71008[10][10];
  wire [31:0] array_index_71010[10];
  wire [31:0] add_71011;
  wire [31:0] array_index_71012[10];
  wire [31:0] add_71013;
  wire [31:0] array_update_71014[10];
  wire [31:0] array_update_71015[10];
  wire [31:0] array_update_71016[10][10];
  wire [31:0] array_update_71018[10][10];
  wire [31:0] array_index_71020[10];
  wire [31:0] add_71021;
  wire [31:0] array_index_71022[10];
  wire [31:0] add_71023;
  wire [31:0] array_update_71024[10];
  wire [31:0] array_update_71025[10];
  wire [31:0] array_update_71026[10][10];
  wire [31:0] array_update_71028[10][10];
  wire [31:0] array_index_71030[10];
  wire [31:0] add_71031;
  wire [31:0] array_index_71032[10];
  wire [31:0] add_71033;
  wire [31:0] array_update_71034[10];
  wire [31:0] array_update_71035[10];
  wire [31:0] array_update_71036[10][10];
  wire [31:0] array_update_71038[10][10];
  wire [31:0] array_index_71040[10];
  wire [31:0] add_71041;
  wire [31:0] array_index_71042[10];
  wire [31:0] add_71043;
  wire [31:0] array_update_71044[10];
  wire [31:0] array_update_71045[10];
  wire [31:0] array_update_71046[10][10];
  wire [31:0] array_update_71048[10][10];
  wire [31:0] array_index_71050[10];
  wire [31:0] add_71051;
  wire [31:0] array_index_71052[10];
  wire [31:0] add_71053;
  wire [31:0] array_update_71054[10];
  wire [31:0] array_update_71055[10];
  wire [31:0] array_update_71056[10][10];
  wire [31:0] array_update_71058[10][10];
  wire [31:0] array_index_71060[10];
  wire [31:0] add_71061;
  wire [31:0] array_index_71062[10];
  wire [31:0] add_71063;
  wire [31:0] array_update_71064[10];
  wire [31:0] array_update_71065[10];
  wire [31:0] array_update_71066[10][10];
  wire [31:0] array_update_71068[10][10];
  wire [31:0] array_index_71070[10];
  wire [31:0] add_71071;
  wire [31:0] array_index_71072[10];
  wire [31:0] add_71073;
  wire [31:0] array_update_71074[10];
  wire [31:0] array_update_71075[10];
  wire [31:0] array_update_71076[10][10];
  wire [31:0] array_update_71078[10][10];
  wire [31:0] array_index_71080[10];
  wire [31:0] add_71081;
  wire [31:0] array_index_71082[10];
  wire [31:0] add_71083;
  wire [31:0] array_update_71084[10];
  wire [31:0] array_update_71085[10];
  wire [31:0] array_update_71086[10][10];
  wire [31:0] array_update_71088[10][10];
  wire [31:0] array_index_71090[10];
  wire [31:0] add_71091;
  wire [31:0] array_index_71092[10];
  wire [31:0] add_71093;
  wire [31:0] array_update_71094[10];
  wire [31:0] array_update_71096[10];
  wire [31:0] array_update_71098[10][10];
  wire [31:0] add_71099;
  wire [31:0] array_update_71100[10][10];
  wire [31:0] add_71101;
  wire [31:0] array_index_71102[10];
  wire [31:0] literal_71103;
  wire [31:0] array_index_71104[10];
  wire [31:0] literal_71105;
  wire [31:0] array_update_71106[10];
  wire [31:0] array_update_71107[10];
  wire [31:0] array_update_71108[10][10];
  wire [31:0] array_update_71110[10][10];
  wire [31:0] array_index_71112[10];
  wire [31:0] add_71113;
  wire [31:0] array_index_71114[10];
  wire [31:0] add_71115;
  wire [31:0] array_update_71116[10];
  wire [31:0] array_update_71117[10];
  wire [31:0] array_update_71118[10][10];
  wire [31:0] array_update_71120[10][10];
  wire [31:0] array_index_71122[10];
  wire [31:0] add_71123;
  wire [31:0] array_index_71124[10];
  wire [31:0] add_71125;
  wire [31:0] array_update_71126[10];
  wire [31:0] array_update_71127[10];
  wire [31:0] array_update_71128[10][10];
  wire [31:0] array_update_71130[10][10];
  wire [31:0] array_index_71132[10];
  wire [31:0] add_71133;
  wire [31:0] array_index_71134[10];
  wire [31:0] add_71135;
  wire [31:0] array_update_71136[10];
  wire [31:0] array_update_71137[10];
  wire [31:0] array_update_71138[10][10];
  wire [31:0] array_update_71140[10][10];
  wire [31:0] array_index_71142[10];
  wire [31:0] add_71143;
  wire [31:0] array_index_71144[10];
  wire [31:0] add_71145;
  wire [31:0] array_update_71146[10];
  wire [31:0] array_update_71147[10];
  wire [31:0] array_update_71148[10][10];
  wire [31:0] array_update_71150[10][10];
  wire [31:0] array_index_71152[10];
  wire [31:0] add_71153;
  wire [31:0] array_index_71154[10];
  wire [31:0] add_71155;
  wire [31:0] array_update_71156[10];
  wire [31:0] array_update_71157[10];
  wire [31:0] array_update_71158[10][10];
  wire [31:0] array_update_71160[10][10];
  wire [31:0] array_index_71162[10];
  wire [31:0] add_71163;
  wire [31:0] array_index_71164[10];
  wire [31:0] add_71165;
  wire [31:0] array_update_71166[10];
  wire [31:0] array_update_71167[10];
  wire [31:0] array_update_71168[10][10];
  wire [31:0] array_update_71170[10][10];
  wire [31:0] array_index_71172[10];
  wire [31:0] add_71173;
  wire [31:0] array_index_71174[10];
  wire [31:0] add_71175;
  wire [31:0] array_update_71176[10];
  wire [31:0] array_update_71177[10];
  wire [31:0] array_update_71178[10][10];
  wire [31:0] array_update_71180[10][10];
  wire [31:0] array_index_71182[10];
  wire [31:0] add_71183;
  wire [31:0] array_index_71184[10];
  wire [31:0] add_71185;
  wire [31:0] array_update_71186[10];
  wire [31:0] array_update_71187[10];
  wire [31:0] array_update_71188[10][10];
  wire [31:0] array_update_71190[10][10];
  wire [31:0] array_index_71192[10];
  wire [31:0] add_71193;
  wire [31:0] array_index_71194[10];
  wire [31:0] add_71195;
  wire [31:0] array_update_71196[10];
  wire [31:0] array_update_71198[10];
  wire [31:0] array_update_71200[10][10];
  wire [31:0] add_71201;
  wire [31:0] array_update_71202[10][10];
  wire [31:0] add_71203;
  wire [31:0] array_index_71204[10];
  wire [31:0] literal_71205;
  wire [31:0] array_index_71206[10];
  wire [31:0] literal_71207;
  wire [31:0] array_update_71208[10];
  wire [31:0] array_update_71209[10];
  wire [31:0] array_update_71210[10][10];
  wire [31:0] array_update_71212[10][10];
  wire [31:0] array_index_71214[10];
  wire [31:0] add_71215;
  wire [31:0] array_index_71216[10];
  wire [31:0] add_71217;
  wire [31:0] array_update_71218[10];
  wire [31:0] array_update_71219[10];
  wire [31:0] array_update_71220[10][10];
  wire [31:0] array_update_71222[10][10];
  wire [31:0] array_index_71224[10];
  wire [31:0] add_71225;
  wire [31:0] array_index_71226[10];
  wire [31:0] add_71227;
  wire [31:0] array_update_71228[10];
  wire [31:0] array_update_71229[10];
  wire [31:0] array_update_71230[10][10];
  wire [31:0] array_update_71232[10][10];
  wire [31:0] array_index_71234[10];
  wire [31:0] add_71235;
  wire [31:0] array_index_71236[10];
  wire [31:0] add_71237;
  wire [31:0] array_update_71238[10];
  wire [31:0] array_update_71239[10];
  wire [31:0] array_update_71240[10][10];
  wire [31:0] array_update_71242[10][10];
  wire [31:0] array_index_71244[10];
  wire [31:0] add_71245;
  wire [31:0] array_index_71246[10];
  wire [31:0] add_71247;
  wire [31:0] array_update_71248[10];
  wire [31:0] array_update_71249[10];
  wire [31:0] array_update_71250[10][10];
  wire [31:0] array_update_71252[10][10];
  wire [31:0] array_index_71254[10];
  wire [31:0] add_71255;
  wire [31:0] array_index_71256[10];
  wire [31:0] add_71257;
  wire [31:0] array_update_71258[10];
  wire [31:0] array_update_71259[10];
  wire [31:0] array_update_71260[10][10];
  wire [31:0] array_update_71262[10][10];
  wire [31:0] array_index_71264[10];
  wire [31:0] add_71265;
  wire [31:0] array_index_71266[10];
  wire [31:0] add_71267;
  wire [31:0] array_update_71268[10];
  wire [31:0] array_update_71269[10];
  wire [31:0] array_update_71270[10][10];
  wire [31:0] array_update_71272[10][10];
  wire [31:0] array_index_71274[10];
  wire [31:0] add_71275;
  wire [31:0] array_index_71276[10];
  wire [31:0] add_71277;
  wire [31:0] array_update_71278[10];
  wire [31:0] array_update_71279[10];
  wire [31:0] array_update_71280[10][10];
  wire [31:0] array_update_71282[10][10];
  wire [31:0] array_index_71284[10];
  wire [31:0] add_71285;
  wire [31:0] array_index_71286[10];
  wire [31:0] add_71287;
  wire [31:0] array_update_71288[10];
  wire [31:0] array_update_71289[10];
  wire [31:0] array_update_71290[10][10];
  wire [31:0] array_update_71292[10][10];
  wire [31:0] array_index_71294[10];
  wire [31:0] add_71295;
  wire [31:0] array_index_71296[10];
  wire [31:0] add_71297;
  wire [31:0] array_update_71298[10];
  wire [31:0] array_update_71300[10];
  wire [31:0] array_update_71302[10][10];
  wire [31:0] add_71303;
  wire [31:0] array_update_71304[10][10];
  wire [31:0] add_71305;
  wire [31:0] array_index_71306[10];
  wire [31:0] literal_71307;
  wire [31:0] array_index_71308[10];
  wire [31:0] literal_71309;
  wire [31:0] array_update_71310[10];
  wire [31:0] array_update_71311[10];
  wire [31:0] array_update_71312[10][10];
  wire [31:0] array_update_71314[10][10];
  wire [31:0] array_index_71316[10];
  wire [31:0] add_71317;
  wire [31:0] array_index_71318[10];
  wire [31:0] add_71319;
  wire [31:0] array_update_71320[10];
  wire [31:0] array_update_71321[10];
  wire [31:0] array_update_71322[10][10];
  wire [31:0] array_update_71324[10][10];
  wire [31:0] array_index_71326[10];
  wire [31:0] add_71327;
  wire [31:0] array_index_71328[10];
  wire [31:0] add_71329;
  wire [31:0] array_update_71330[10];
  wire [31:0] array_update_71331[10];
  wire [31:0] array_update_71332[10][10];
  wire [31:0] array_update_71334[10][10];
  wire [31:0] array_index_71336[10];
  wire [31:0] add_71337;
  wire [31:0] array_index_71338[10];
  wire [31:0] add_71339;
  wire [31:0] array_update_71340[10];
  wire [31:0] array_update_71341[10];
  wire [31:0] array_update_71342[10][10];
  wire [31:0] array_update_71344[10][10];
  wire [31:0] array_index_71346[10];
  wire [31:0] add_71347;
  wire [31:0] array_index_71348[10];
  wire [31:0] add_71349;
  wire [31:0] array_update_71350[10];
  wire [31:0] array_update_71351[10];
  wire [31:0] array_update_71352[10][10];
  wire [31:0] array_update_71354[10][10];
  wire [31:0] array_index_71356[10];
  wire [31:0] add_71357;
  wire [31:0] array_index_71358[10];
  wire [31:0] add_71359;
  wire [31:0] array_update_71360[10];
  wire [31:0] array_update_71361[10];
  wire [31:0] array_update_71362[10][10];
  wire [31:0] array_update_71364[10][10];
  wire [31:0] array_index_71366[10];
  wire [31:0] add_71367;
  wire [31:0] array_index_71368[10];
  wire [31:0] add_71369;
  wire [31:0] array_update_71370[10];
  wire [31:0] array_update_71371[10];
  wire [31:0] array_update_71372[10][10];
  wire [31:0] array_update_71374[10][10];
  wire [31:0] array_index_71376[10];
  wire [31:0] add_71377;
  wire [31:0] array_index_71378[10];
  wire [31:0] add_71379;
  wire [31:0] array_update_71380[10];
  wire [31:0] array_update_71381[10];
  wire [31:0] array_update_71382[10][10];
  wire [31:0] array_update_71384[10][10];
  wire [31:0] array_index_71386[10];
  wire [31:0] add_71387;
  wire [31:0] array_index_71388[10];
  wire [31:0] add_71389;
  wire [31:0] array_update_71390[10];
  wire [31:0] array_update_71391[10];
  wire [31:0] array_update_71392[10][10];
  wire [31:0] array_update_71394[10][10];
  wire [31:0] array_index_71396[10];
  wire [31:0] add_71397;
  wire [31:0] array_index_71398[10];
  wire [31:0] add_71399;
  wire [31:0] array_update_71400[10];
  wire [31:0] array_update_71402[10];
  wire [31:0] array_update_71404[10][10];
  wire [31:0] add_71405;
  wire [31:0] array_update_71406[10][10];
  wire [31:0] add_71407;
  wire [31:0] array_index_71408[10];
  wire [31:0] literal_71409;
  wire [31:0] array_index_71410[10];
  wire [31:0] literal_71411;
  wire [31:0] array_update_71412[10];
  wire [31:0] array_update_71413[10];
  wire [31:0] array_update_71414[10][10];
  wire [31:0] array_update_71416[10][10];
  wire [31:0] array_index_71418[10];
  wire [31:0] add_71419;
  wire [31:0] array_index_71420[10];
  wire [31:0] add_71421;
  wire [31:0] array_update_71422[10];
  wire [31:0] array_update_71423[10];
  wire [31:0] array_update_71424[10][10];
  wire [31:0] array_update_71426[10][10];
  wire [31:0] array_index_71428[10];
  wire [31:0] add_71429;
  wire [31:0] array_index_71430[10];
  wire [31:0] add_71431;
  wire [31:0] array_update_71432[10];
  wire [31:0] array_update_71433[10];
  wire [31:0] array_update_71434[10][10];
  wire [31:0] array_update_71436[10][10];
  wire [31:0] array_index_71438[10];
  wire [31:0] add_71439;
  wire [31:0] array_index_71440[10];
  wire [31:0] add_71441;
  wire [31:0] array_update_71442[10];
  wire [31:0] array_update_71443[10];
  wire [31:0] array_update_71444[10][10];
  wire [31:0] array_update_71446[10][10];
  wire [31:0] array_index_71448[10];
  wire [31:0] add_71449;
  wire [31:0] array_index_71450[10];
  wire [31:0] add_71451;
  wire [31:0] array_update_71452[10];
  wire [31:0] array_update_71453[10];
  wire [31:0] array_update_71454[10][10];
  wire [31:0] array_update_71456[10][10];
  wire [31:0] array_index_71458[10];
  wire [31:0] add_71459;
  wire [31:0] array_index_71460[10];
  wire [31:0] add_71461;
  wire [31:0] array_update_71462[10];
  wire [31:0] array_update_71463[10];
  wire [31:0] array_update_71464[10][10];
  wire [31:0] array_update_71466[10][10];
  wire [31:0] array_index_71468[10];
  wire [31:0] add_71469;
  wire [31:0] array_index_71470[10];
  wire [31:0] add_71471;
  wire [31:0] array_update_71472[10];
  wire [31:0] array_update_71473[10];
  wire [31:0] array_update_71474[10][10];
  wire [31:0] array_update_71476[10][10];
  wire [31:0] array_index_71478[10];
  wire [31:0] add_71479;
  wire [31:0] array_index_71480[10];
  wire [31:0] add_71481;
  wire [31:0] array_update_71482[10];
  wire [31:0] array_update_71483[10];
  wire [31:0] array_update_71484[10][10];
  wire [31:0] array_update_71486[10][10];
  wire [31:0] array_index_71488[10];
  wire [31:0] add_71489;
  wire [31:0] array_index_71490[10];
  wire [31:0] add_71491;
  wire [31:0] array_update_71492[10];
  wire [31:0] array_update_71493[10];
  wire [31:0] array_update_71494[10][10];
  wire [31:0] array_update_71496[10][10];
  wire [31:0] array_index_71498[10];
  wire [31:0] add_71499;
  wire [31:0] array_index_71500[10];
  wire [31:0] add_71501;
  wire [31:0] array_update_71502[10];
  wire [31:0] array_update_71504[10];
  wire [31:0] array_update_71506[10][10];
  wire [31:0] add_71507;
  wire [31:0] array_update_71508[10][10];
  wire [31:0] add_71509;
  wire [31:0] array_index_71510[10];
  wire [31:0] literal_71511;
  wire [31:0] array_index_71512[10];
  wire [31:0] literal_71513;
  wire [31:0] array_update_71514[10];
  wire [31:0] array_update_71515[10];
  wire [31:0] array_update_71516[10][10];
  wire [31:0] array_update_71518[10][10];
  wire [31:0] array_index_71520[10];
  wire [31:0] add_71521;
  wire [31:0] array_index_71522[10];
  wire [31:0] add_71523;
  wire [31:0] array_update_71524[10];
  wire [31:0] array_update_71525[10];
  wire [31:0] array_update_71526[10][10];
  wire [31:0] array_update_71528[10][10];
  wire [31:0] array_index_71530[10];
  wire [31:0] add_71531;
  wire [31:0] array_index_71532[10];
  wire [31:0] add_71533;
  wire [31:0] array_update_71534[10];
  wire [31:0] array_update_71535[10];
  wire [31:0] array_update_71536[10][10];
  wire [31:0] array_update_71538[10][10];
  wire [31:0] array_index_71540[10];
  wire [31:0] add_71541;
  wire [31:0] array_index_71542[10];
  wire [31:0] add_71543;
  wire [31:0] array_update_71544[10];
  wire [31:0] array_update_71545[10];
  wire [31:0] array_update_71546[10][10];
  wire [31:0] array_update_71548[10][10];
  wire [31:0] array_index_71550[10];
  wire [31:0] add_71551;
  wire [31:0] array_index_71552[10];
  wire [31:0] add_71553;
  wire [31:0] array_update_71554[10];
  wire [31:0] array_update_71555[10];
  wire [31:0] array_update_71556[10][10];
  wire [31:0] array_update_71558[10][10];
  wire [31:0] array_index_71560[10];
  wire [31:0] add_71561;
  wire [31:0] array_index_71562[10];
  wire [31:0] add_71563;
  wire [31:0] array_update_71564[10];
  wire [31:0] array_update_71565[10];
  wire [31:0] array_update_71566[10][10];
  wire [31:0] array_update_71568[10][10];
  wire [31:0] array_index_71570[10];
  wire [31:0] add_71571;
  wire [31:0] array_index_71572[10];
  wire [31:0] add_71573;
  wire [31:0] array_update_71574[10];
  wire [31:0] array_update_71575[10];
  wire [31:0] array_update_71576[10][10];
  wire [31:0] array_update_71578[10][10];
  wire [31:0] array_index_71580[10];
  wire [31:0] add_71581;
  wire [31:0] array_index_71582[10];
  wire [31:0] add_71583;
  wire [31:0] array_update_71584[10];
  wire [31:0] array_update_71585[10];
  wire [31:0] array_update_71586[10][10];
  wire [31:0] array_update_71588[10][10];
  wire [31:0] array_index_71590[10];
  wire [31:0] add_71591;
  wire [31:0] array_index_71592[10];
  wire [31:0] add_71593;
  wire [31:0] array_update_71594[10];
  wire [31:0] array_update_71595[10];
  wire [31:0] array_update_71596[10][10];
  wire [31:0] array_update_71598[10][10];
  wire [31:0] array_index_71600[10];
  wire [31:0] add_71601;
  wire [31:0] array_index_71602[10];
  wire [31:0] add_71603;
  wire [31:0] array_update_71604[10];
  wire [31:0] array_update_71606[10];
  wire [31:0] array_update_71608[10][10];
  wire [31:0] add_71609;
  wire [31:0] array_update_71610[10][10];
  wire [31:0] add_71611;
  wire [31:0] array_index_71612[10];
  wire [31:0] literal_71613;
  wire [31:0] array_index_71614[10];
  wire [31:0] literal_71615;
  wire [31:0] array_update_71616[10];
  wire [31:0] array_update_71617[10];
  wire [31:0] array_update_71618[10][10];
  wire [31:0] array_update_71620[10][10];
  wire [31:0] array_index_71622[10];
  wire [31:0] add_71623;
  wire [31:0] array_index_71624[10];
  wire [31:0] add_71625;
  wire [31:0] array_update_71626[10];
  wire [31:0] array_update_71627[10];
  wire [31:0] array_update_71628[10][10];
  wire [31:0] array_update_71630[10][10];
  wire [31:0] array_index_71632[10];
  wire [31:0] add_71633;
  wire [31:0] array_index_71634[10];
  wire [31:0] add_71635;
  wire [31:0] array_update_71636[10];
  wire [31:0] array_update_71637[10];
  wire [31:0] array_update_71638[10][10];
  wire [31:0] array_update_71640[10][10];
  wire [31:0] array_index_71642[10];
  wire [31:0] add_71643;
  wire [31:0] array_index_71644[10];
  wire [31:0] add_71645;
  wire [31:0] array_update_71646[10];
  wire [31:0] array_update_71647[10];
  wire [31:0] array_update_71648[10][10];
  wire [31:0] array_update_71650[10][10];
  wire [31:0] array_index_71652[10];
  wire [31:0] add_71653;
  wire [31:0] array_index_71654[10];
  wire [31:0] add_71655;
  wire [31:0] array_update_71656[10];
  wire [31:0] array_update_71657[10];
  wire [31:0] array_update_71658[10][10];
  wire [31:0] array_update_71660[10][10];
  wire [31:0] array_index_71662[10];
  wire [31:0] add_71663;
  wire [31:0] array_index_71664[10];
  wire [31:0] add_71665;
  wire [31:0] array_update_71666[10];
  wire [31:0] array_update_71667[10];
  wire [31:0] array_update_71668[10][10];
  wire [31:0] array_update_71670[10][10];
  wire [31:0] array_index_71672[10];
  wire [31:0] add_71673;
  wire [31:0] array_index_71674[10];
  wire [31:0] add_71675;
  wire [31:0] array_update_71676[10];
  wire [31:0] array_update_71677[10];
  wire [31:0] array_update_71678[10][10];
  wire [31:0] array_update_71680[10][10];
  wire [31:0] array_index_71682[10];
  wire [31:0] add_71683;
  wire [31:0] array_index_71684[10];
  wire [31:0] add_71685;
  wire [31:0] array_update_71686[10];
  wire [31:0] array_update_71687[10];
  wire [31:0] array_update_71688[10][10];
  wire [31:0] array_update_71690[10][10];
  wire [31:0] array_index_71692[10];
  wire [31:0] add_71693;
  wire [31:0] array_index_71694[10];
  wire [31:0] add_71695;
  wire [31:0] array_update_71696[10];
  wire [31:0] array_update_71697[10];
  wire [31:0] array_update_71698[10][10];
  wire [31:0] array_update_71700[10][10];
  wire [31:0] array_index_71702[10];
  wire [31:0] add_71703;
  wire [31:0] array_index_71704[10];
  wire [31:0] add_71705;
  wire [31:0] array_update_71706[10];
  wire [31:0] array_update_71708[10];
  wire [31:0] array_update_71710[10][10];
  wire [31:0] add_71711;
  wire [31:0] array_update_71712[10][10];
  wire [31:0] add_71713;
  wire [31:0] array_index_71714[10];
  wire [31:0] literal_71715;
  wire [31:0] array_index_71716[10];
  wire [31:0] literal_71717;
  wire [31:0] array_update_71718[10];
  wire [31:0] array_update_71719[10];
  wire [31:0] array_update_71720[10][10];
  wire [31:0] array_update_71722[10][10];
  wire [31:0] array_index_71724[10];
  wire [31:0] add_71725;
  wire [31:0] array_index_71726[10];
  wire [31:0] add_71727;
  wire [31:0] array_update_71728[10];
  wire [31:0] array_update_71729[10];
  wire [31:0] array_update_71730[10][10];
  wire [31:0] array_update_71732[10][10];
  wire [31:0] array_index_71734[10];
  wire [31:0] add_71735;
  wire [31:0] array_index_71736[10];
  wire [31:0] add_71737;
  wire [31:0] array_update_71738[10];
  wire [31:0] array_update_71739[10];
  wire [31:0] array_update_71740[10][10];
  wire [31:0] array_update_71742[10][10];
  wire [31:0] array_index_71744[10];
  wire [31:0] add_71745;
  wire [31:0] array_index_71746[10];
  wire [31:0] add_71747;
  wire [31:0] array_update_71748[10];
  wire [31:0] array_update_71749[10];
  wire [31:0] array_update_71750[10][10];
  wire [31:0] array_update_71752[10][10];
  wire [31:0] array_index_71754[10];
  wire [31:0] add_71755;
  wire [31:0] array_index_71756[10];
  wire [31:0] add_71757;
  wire [31:0] array_update_71758[10];
  wire [31:0] array_update_71759[10];
  wire [31:0] array_update_71760[10][10];
  wire [31:0] array_update_71762[10][10];
  wire [31:0] array_index_71764[10];
  wire [31:0] add_71765;
  wire [31:0] array_index_71766[10];
  wire [31:0] add_71767;
  wire [31:0] array_update_71768[10];
  wire [31:0] array_update_71769[10];
  wire [31:0] array_update_71770[10][10];
  wire [31:0] array_update_71772[10][10];
  wire [31:0] array_index_71774[10];
  wire [31:0] add_71775;
  wire [31:0] array_index_71776[10];
  wire [31:0] add_71777;
  wire [31:0] array_update_71778[10];
  wire [31:0] array_update_71779[10];
  wire [31:0] array_update_71780[10][10];
  wire [31:0] array_update_71782[10][10];
  wire [31:0] array_index_71784[10];
  wire [31:0] add_71785;
  wire [31:0] array_index_71786[10];
  wire [31:0] add_71787;
  wire [31:0] array_update_71788[10];
  wire [31:0] array_update_71789[10];
  wire [31:0] array_update_71790[10][10];
  wire [31:0] array_update_71792[10][10];
  wire [31:0] array_index_71794[10];
  wire [31:0] add_71795;
  wire [31:0] array_index_71796[10];
  wire [31:0] add_71797;
  wire [31:0] array_update_71798[10];
  wire [31:0] array_update_71799[10];
  wire [31:0] array_update_71800[10][10];
  wire [31:0] array_update_71802[10][10];
  wire [31:0] array_index_71804[10];
  wire [31:0] add_71805;
  wire [31:0] array_index_71806[10];
  wire [31:0] add_71807;
  wire [31:0] array_update_71808[10];
  wire [31:0] array_update_71810[10];
  wire [31:0] array_update_71812[10][10];
  wire [31:0] add_71813;
  wire [31:0] array_update_71814[10][10];
  wire [31:0] add_71815;
  wire [31:0] array_index_71816[10];
  wire [31:0] literal_71817;
  wire [31:0] array_index_71818[10];
  wire [31:0] literal_71819;
  wire [31:0] array_update_71820[10];
  wire [31:0] array_update_71821[10];
  wire [31:0] array_update_71822[10][10];
  wire [31:0] array_update_71824[10][10];
  wire [31:0] array_index_71826[10];
  wire [31:0] add_71827;
  wire [31:0] array_index_71828[10];
  wire [31:0] add_71829;
  wire [31:0] array_update_71830[10];
  wire [31:0] array_update_71831[10];
  wire [31:0] array_update_71832[10][10];
  wire [31:0] array_update_71834[10][10];
  wire [31:0] array_index_71836[10];
  wire [31:0] add_71837;
  wire [31:0] array_index_71838[10];
  wire [31:0] add_71839;
  wire [31:0] array_update_71840[10];
  wire [31:0] array_update_71841[10];
  wire [31:0] array_update_71842[10][10];
  wire [31:0] array_update_71844[10][10];
  wire [31:0] array_index_71846[10];
  wire [31:0] add_71847;
  wire [31:0] array_index_71848[10];
  wire [31:0] add_71849;
  wire [31:0] array_update_71850[10];
  wire [31:0] array_update_71851[10];
  wire [31:0] array_update_71852[10][10];
  wire [31:0] array_update_71854[10][10];
  wire [31:0] array_index_71856[10];
  wire [31:0] add_71857;
  wire [31:0] array_index_71858[10];
  wire [31:0] add_71859;
  wire [31:0] array_update_71860[10];
  wire [31:0] array_update_71861[10];
  wire [31:0] array_update_71862[10][10];
  wire [31:0] array_update_71864[10][10];
  wire [31:0] array_index_71866[10];
  wire [31:0] add_71867;
  wire [31:0] array_index_71868[10];
  wire [31:0] add_71869;
  wire [31:0] array_update_71870[10];
  wire [31:0] array_update_71871[10];
  wire [31:0] array_update_71872[10][10];
  wire [31:0] array_update_71874[10][10];
  wire [31:0] array_index_71876[10];
  wire [31:0] add_71877;
  wire [31:0] array_index_71878[10];
  wire [31:0] add_71879;
  wire [31:0] array_update_71880[10];
  wire [31:0] array_update_71881[10];
  wire [31:0] array_update_71882[10][10];
  wire [31:0] array_update_71884[10][10];
  wire [31:0] array_index_71886[10];
  wire [31:0] add_71887;
  wire [31:0] array_index_71888[10];
  wire [31:0] add_71889;
  wire [31:0] array_update_71890[10];
  wire [31:0] array_update_71891[10];
  wire [31:0] array_update_71892[10][10];
  wire [31:0] array_update_71894[10][10];
  wire [31:0] array_index_71896[10];
  wire [31:0] add_71897;
  wire [31:0] array_index_71898[10];
  wire [31:0] add_71899;
  wire [31:0] array_update_71900[10];
  wire [31:0] array_update_71901[10];
  wire [31:0] array_update_71902[10][10];
  wire [31:0] array_update_71904[10][10];
  wire [31:0] array_index_71906[10];
  wire [31:0] add_71907;
  wire [31:0] array_index_71908[10];
  wire [31:0] add_71909;
  wire [31:0] array_update_71910[10];
  wire [31:0] array_update_71912[10];
  wire [31:0] array_update_71914[10][10];
  wire [31:0] add_71915;
  wire [31:0] array_update_71916[10][10];
  wire [31:0] add_71917;
  wire [31:0] array_index_71918[10];
  wire [31:0] literal_71919;
  wire [31:0] array_index_71920[10];
  wire [31:0] literal_71921;
  wire [31:0] array_update_71922[10];
  wire [31:0] array_update_71923[10];
  wire [31:0] array_update_71924[10][10];
  wire [31:0] array_update_71926[10][10];
  wire [31:0] array_index_71928[10];
  wire [31:0] add_71929;
  wire [31:0] array_index_71930[10];
  wire [31:0] add_71931;
  wire [31:0] array_update_71932[10];
  wire [31:0] array_update_71933[10];
  wire [31:0] array_update_71934[10][10];
  wire [31:0] array_update_71936[10][10];
  wire [31:0] array_index_71938[10];
  wire [31:0] add_71939;
  wire [31:0] array_index_71940[10];
  wire [31:0] add_71941;
  wire [31:0] array_update_71942[10];
  wire [31:0] array_update_71943[10];
  wire [31:0] array_update_71944[10][10];
  wire [31:0] array_update_71946[10][10];
  wire [31:0] array_index_71948[10];
  wire [31:0] add_71949;
  wire [31:0] array_index_71950[10];
  wire [31:0] add_71951;
  wire [31:0] array_update_71952[10];
  wire [31:0] array_update_71953[10];
  wire [31:0] array_update_71954[10][10];
  wire [31:0] array_update_71956[10][10];
  wire [31:0] array_index_71958[10];
  wire [31:0] add_71959;
  wire [31:0] array_index_71960[10];
  wire [31:0] add_71961;
  wire [31:0] array_update_71962[10];
  wire [31:0] array_update_71963[10];
  wire [31:0] array_update_71964[10][10];
  wire [31:0] array_update_71966[10][10];
  wire [31:0] array_index_71968[10];
  wire [31:0] add_71969;
  wire [31:0] array_index_71970[10];
  wire [31:0] add_71971;
  wire [31:0] array_update_71972[10];
  wire [31:0] array_update_71973[10];
  wire [31:0] array_update_71974[10][10];
  wire [31:0] array_update_71976[10][10];
  wire [31:0] array_index_71978[10];
  wire [31:0] add_71979;
  wire [31:0] array_index_71980[10];
  wire [31:0] add_71981;
  wire [31:0] array_update_71982[10];
  wire [31:0] array_update_71983[10];
  wire [31:0] array_update_71984[10][10];
  wire [31:0] array_update_71986[10][10];
  wire [31:0] array_index_71988[10];
  wire [31:0] add_71989;
  wire [31:0] array_index_71990[10];
  wire [31:0] add_71991;
  wire [31:0] array_update_71992[10];
  wire [31:0] array_update_71993[10];
  wire [31:0] array_update_71994[10][10];
  wire [31:0] array_update_71996[10][10];
  wire [31:0] array_index_71998[10];
  wire [31:0] add_71999;
  wire [31:0] array_index_72000[10];
  wire [31:0] add_72001;
  wire [31:0] array_update_72002[10];
  wire [31:0] array_update_72003[10];
  wire [31:0] array_update_72004[10][10];
  wire [31:0] array_update_72006[10][10];
  wire [31:0] literal_72009;
  wire [31:0] array_index_72010[10];
  wire [31:0] add_72011;
  wire [31:0] array_index_72012[10];
  wire [31:0] add_72013;
  wire [31:0] array_index_72014[10];
  wire [31:0] literal_72016;
  wire [31:0] array_update_72017[10];
  wire [31:0] array_update_72018[10];
  wire [31:0] array_update_72019[10];
  wire [31:0] array_update_72020[10][10];
  wire [31:0] array_update_72021[10][10];
  wire [31:0] literal_72022;
  wire [31:0] array_update_72023[10][10];
  wire [31:0] array_index_72024[10];
  wire [31:0] array_index_72025[10];
  wire [31:0] array_index_72026[10];
  wire [31:0] smul_72030;
  wire [31:0] add_72032;
  wire [31:0] array_update_72034[10];
  wire [31:0] add_72035;
  wire [31:0] array_update_72036[10][10];
  wire [31:0] array_index_72038[10];
  wire [31:0] array_index_72039[10];
  wire [31:0] smul_72043;
  wire [31:0] add_72045;
  wire [31:0] array_update_72047[10];
  wire [31:0] add_72048;
  wire [31:0] array_update_72049[10][10];
  wire [31:0] array_index_72051[10];
  wire [31:0] array_index_72052[10];
  wire [31:0] smul_72056;
  wire [31:0] add_72058;
  wire [31:0] array_update_72060[10];
  wire [31:0] add_72061;
  wire [31:0] array_update_72062[10][10];
  wire [31:0] array_index_72064[10];
  wire [31:0] array_index_72065[10];
  wire [31:0] smul_72069;
  wire [31:0] add_72071;
  wire [31:0] array_update_72073[10];
  wire [31:0] add_72074;
  wire [31:0] array_update_72075[10][10];
  wire [31:0] array_index_72077[10];
  wire [31:0] array_index_72078[10];
  wire [31:0] smul_72082;
  wire [31:0] add_72084;
  wire [31:0] array_update_72086[10];
  wire [31:0] add_72087;
  wire [31:0] array_update_72088[10][10];
  wire [31:0] array_index_72090[10];
  wire [31:0] array_index_72091[10];
  wire [31:0] smul_72095;
  wire [31:0] add_72097;
  wire [31:0] array_update_72099[10];
  wire [31:0] add_72100;
  wire [31:0] array_update_72101[10][10];
  wire [31:0] array_index_72103[10];
  wire [31:0] array_index_72104[10];
  wire [31:0] smul_72108;
  wire [31:0] add_72110;
  wire [31:0] array_update_72112[10];
  wire [31:0] add_72113;
  wire [31:0] array_update_72114[10][10];
  wire [31:0] array_index_72116[10];
  wire [31:0] array_index_72117[10];
  wire [31:0] smul_72121;
  wire [31:0] add_72123;
  wire [31:0] array_update_72125[10];
  wire [31:0] add_72126;
  wire [31:0] array_update_72127[10][10];
  wire [31:0] array_index_72129[10];
  wire [31:0] array_index_72130[10];
  wire [31:0] smul_72134;
  wire [31:0] add_72136;
  wire [31:0] array_update_72138[10];
  wire [31:0] add_72139;
  wire [31:0] array_update_72140[10][10];
  wire [31:0] array_index_72142[10];
  wire [31:0] array_index_72143[10];
  wire [31:0] smul_72147;
  wire [31:0] add_72149;
  wire [31:0] array_update_72150[10];
  wire [31:0] array_update_72151[10][10];
  wire [31:0] array_index_72153[10];
  wire [31:0] add_72155;
  wire [31:0] array_update_72156[10];
  wire [31:0] literal_72157;
  wire [31:0] array_update_72158[10][10];
  wire [31:0] array_index_72160[10];
  wire [31:0] array_index_72161[10];
  wire [31:0] smul_72165;
  wire [31:0] add_72167;
  wire [31:0] array_update_72169[10];
  wire [31:0] add_72170;
  wire [31:0] array_update_72171[10][10];
  wire [31:0] array_index_72173[10];
  wire [31:0] array_index_72174[10];
  wire [31:0] smul_72178;
  wire [31:0] add_72180;
  wire [31:0] array_update_72182[10];
  wire [31:0] add_72183;
  wire [31:0] array_update_72184[10][10];
  wire [31:0] array_index_72186[10];
  wire [31:0] array_index_72187[10];
  wire [31:0] smul_72191;
  wire [31:0] add_72193;
  wire [31:0] array_update_72195[10];
  wire [31:0] add_72196;
  wire [31:0] array_update_72197[10][10];
  wire [31:0] array_index_72199[10];
  wire [31:0] array_index_72200[10];
  wire [31:0] smul_72204;
  wire [31:0] add_72206;
  wire [31:0] array_update_72208[10];
  wire [31:0] add_72209;
  wire [31:0] array_update_72210[10][10];
  wire [31:0] array_index_72212[10];
  wire [31:0] array_index_72213[10];
  wire [31:0] smul_72217;
  wire [31:0] add_72219;
  wire [31:0] array_update_72221[10];
  wire [31:0] add_72222;
  wire [31:0] array_update_72223[10][10];
  wire [31:0] array_index_72225[10];
  wire [31:0] array_index_72226[10];
  wire [31:0] smul_72230;
  wire [31:0] add_72232;
  wire [31:0] array_update_72234[10];
  wire [31:0] add_72235;
  wire [31:0] array_update_72236[10][10];
  wire [31:0] array_index_72238[10];
  wire [31:0] array_index_72239[10];
  wire [31:0] smul_72243;
  wire [31:0] add_72245;
  wire [31:0] array_update_72247[10];
  wire [31:0] add_72248;
  wire [31:0] array_update_72249[10][10];
  wire [31:0] array_index_72251[10];
  wire [31:0] array_index_72252[10];
  wire [31:0] smul_72256;
  wire [31:0] add_72258;
  wire [31:0] array_update_72260[10];
  wire [31:0] add_72261;
  wire [31:0] array_update_72262[10][10];
  wire [31:0] array_index_72264[10];
  wire [31:0] array_index_72265[10];
  wire [31:0] smul_72269;
  wire [31:0] add_72271;
  wire [31:0] array_update_72273[10];
  wire [31:0] add_72274;
  wire [31:0] array_update_72275[10][10];
  wire [31:0] array_index_72277[10];
  wire [31:0] array_index_72278[10];
  wire [31:0] smul_72282;
  wire [31:0] add_72284;
  wire [31:0] array_update_72285[10];
  wire [31:0] array_update_72286[10][10];
  wire [31:0] array_index_72288[10];
  wire [31:0] add_72290;
  wire [31:0] array_update_72291[10];
  wire [31:0] literal_72292;
  wire [31:0] array_update_72293[10][10];
  wire [31:0] array_index_72295[10];
  wire [31:0] array_index_72296[10];
  wire [31:0] smul_72300;
  wire [31:0] add_72302;
  wire [31:0] array_update_72304[10];
  wire [31:0] add_72305;
  wire [31:0] array_update_72306[10][10];
  wire [31:0] array_index_72308[10];
  wire [31:0] array_index_72309[10];
  wire [31:0] smul_72313;
  wire [31:0] add_72315;
  wire [31:0] array_update_72317[10];
  wire [31:0] add_72318;
  wire [31:0] array_update_72319[10][10];
  wire [31:0] array_index_72321[10];
  wire [31:0] array_index_72322[10];
  wire [31:0] smul_72326;
  wire [31:0] add_72328;
  wire [31:0] array_update_72330[10];
  wire [31:0] add_72331;
  wire [31:0] array_update_72332[10][10];
  wire [31:0] array_index_72334[10];
  wire [31:0] array_index_72335[10];
  wire [31:0] smul_72339;
  wire [31:0] add_72341;
  wire [31:0] array_update_72343[10];
  wire [31:0] add_72344;
  wire [31:0] array_update_72345[10][10];
  wire [31:0] array_index_72347[10];
  wire [31:0] array_index_72348[10];
  wire [31:0] smul_72352;
  wire [31:0] add_72354;
  wire [31:0] array_update_72356[10];
  wire [31:0] add_72357;
  wire [31:0] array_update_72358[10][10];
  wire [31:0] array_index_72360[10];
  wire [31:0] array_index_72361[10];
  wire [31:0] smul_72365;
  wire [31:0] add_72367;
  wire [31:0] array_update_72369[10];
  wire [31:0] add_72370;
  wire [31:0] array_update_72371[10][10];
  wire [31:0] array_index_72373[10];
  wire [31:0] array_index_72374[10];
  wire [31:0] smul_72378;
  wire [31:0] add_72380;
  wire [31:0] array_update_72382[10];
  wire [31:0] add_72383;
  wire [31:0] array_update_72384[10][10];
  wire [31:0] array_index_72386[10];
  wire [31:0] array_index_72387[10];
  wire [31:0] smul_72391;
  wire [31:0] add_72393;
  wire [31:0] array_update_72395[10];
  wire [31:0] add_72396;
  wire [31:0] array_update_72397[10][10];
  wire [31:0] array_index_72399[10];
  wire [31:0] array_index_72400[10];
  wire [31:0] smul_72404;
  wire [31:0] add_72406;
  wire [31:0] array_update_72408[10];
  wire [31:0] add_72409;
  wire [31:0] array_update_72410[10][10];
  wire [31:0] array_index_72412[10];
  wire [31:0] array_index_72413[10];
  wire [31:0] smul_72417;
  wire [31:0] add_72419;
  wire [31:0] array_update_72420[10];
  wire [31:0] array_update_72421[10][10];
  wire [31:0] array_index_72423[10];
  wire [31:0] add_72425;
  wire [31:0] array_update_72426[10];
  wire [31:0] literal_72427;
  wire [31:0] array_update_72428[10][10];
  wire [31:0] array_index_72430[10];
  wire [31:0] array_index_72431[10];
  wire [31:0] smul_72435;
  wire [31:0] add_72437;
  wire [31:0] array_update_72439[10];
  wire [31:0] add_72440;
  wire [31:0] array_update_72441[10][10];
  wire [31:0] array_index_72443[10];
  wire [31:0] array_index_72444[10];
  wire [31:0] smul_72448;
  wire [31:0] add_72450;
  wire [31:0] array_update_72452[10];
  wire [31:0] add_72453;
  wire [31:0] array_update_72454[10][10];
  wire [31:0] array_index_72456[10];
  wire [31:0] array_index_72457[10];
  wire [31:0] smul_72461;
  wire [31:0] add_72463;
  wire [31:0] array_update_72465[10];
  wire [31:0] add_72466;
  wire [31:0] array_update_72467[10][10];
  wire [31:0] array_index_72469[10];
  wire [31:0] array_index_72470[10];
  wire [31:0] smul_72474;
  wire [31:0] add_72476;
  wire [31:0] array_update_72478[10];
  wire [31:0] add_72479;
  wire [31:0] array_update_72480[10][10];
  wire [31:0] array_index_72482[10];
  wire [31:0] array_index_72483[10];
  wire [31:0] smul_72487;
  wire [31:0] add_72489;
  wire [31:0] array_update_72491[10];
  wire [31:0] add_72492;
  wire [31:0] array_update_72493[10][10];
  wire [31:0] array_index_72495[10];
  wire [31:0] array_index_72496[10];
  wire [31:0] smul_72500;
  wire [31:0] add_72502;
  wire [31:0] array_update_72504[10];
  wire [31:0] add_72505;
  wire [31:0] array_update_72506[10][10];
  wire [31:0] array_index_72508[10];
  wire [31:0] array_index_72509[10];
  wire [31:0] smul_72513;
  wire [31:0] add_72515;
  wire [31:0] array_update_72517[10];
  wire [31:0] add_72518;
  wire [31:0] array_update_72519[10][10];
  wire [31:0] array_index_72521[10];
  wire [31:0] array_index_72522[10];
  wire [31:0] smul_72526;
  wire [31:0] add_72528;
  wire [31:0] array_update_72530[10];
  wire [31:0] add_72531;
  wire [31:0] array_update_72532[10][10];
  wire [31:0] array_index_72534[10];
  wire [31:0] array_index_72535[10];
  wire [31:0] smul_72539;
  wire [31:0] add_72541;
  wire [31:0] array_update_72543[10];
  wire [31:0] add_72544;
  wire [31:0] array_update_72545[10][10];
  wire [31:0] array_index_72547[10];
  wire [31:0] array_index_72548[10];
  wire [31:0] smul_72552;
  wire [31:0] add_72554;
  wire [31:0] array_update_72555[10];
  wire [31:0] array_update_72556[10][10];
  wire [31:0] array_index_72558[10];
  wire [31:0] add_72560;
  wire [31:0] array_update_72561[10];
  wire [31:0] literal_72562;
  wire [31:0] array_update_72563[10][10];
  wire [31:0] array_index_72565[10];
  wire [31:0] array_index_72566[10];
  wire [31:0] smul_72570;
  wire [31:0] add_72572;
  wire [31:0] array_update_72574[10];
  wire [31:0] add_72575;
  wire [31:0] array_update_72576[10][10];
  wire [31:0] array_index_72578[10];
  wire [31:0] array_index_72579[10];
  wire [31:0] smul_72583;
  wire [31:0] add_72585;
  wire [31:0] array_update_72587[10];
  wire [31:0] add_72588;
  wire [31:0] array_update_72589[10][10];
  wire [31:0] array_index_72591[10];
  wire [31:0] array_index_72592[10];
  wire [31:0] smul_72596;
  wire [31:0] add_72598;
  wire [31:0] array_update_72600[10];
  wire [31:0] add_72601;
  wire [31:0] array_update_72602[10][10];
  wire [31:0] array_index_72604[10];
  wire [31:0] array_index_72605[10];
  wire [31:0] smul_72609;
  wire [31:0] add_72611;
  wire [31:0] array_update_72613[10];
  wire [31:0] add_72614;
  wire [31:0] array_update_72615[10][10];
  wire [31:0] array_index_72617[10];
  wire [31:0] array_index_72618[10];
  wire [31:0] smul_72622;
  wire [31:0] add_72624;
  wire [31:0] array_update_72626[10];
  wire [31:0] add_72627;
  wire [31:0] array_update_72628[10][10];
  wire [31:0] array_index_72630[10];
  wire [31:0] array_index_72631[10];
  wire [31:0] smul_72635;
  wire [31:0] add_72637;
  wire [31:0] array_update_72639[10];
  wire [31:0] add_72640;
  wire [31:0] array_update_72641[10][10];
  wire [31:0] array_index_72643[10];
  wire [31:0] array_index_72644[10];
  wire [31:0] smul_72648;
  wire [31:0] add_72650;
  wire [31:0] array_update_72652[10];
  wire [31:0] add_72653;
  wire [31:0] array_update_72654[10][10];
  wire [31:0] array_index_72656[10];
  wire [31:0] array_index_72657[10];
  wire [31:0] smul_72661;
  wire [31:0] add_72663;
  wire [31:0] array_update_72665[10];
  wire [31:0] add_72666;
  wire [31:0] array_update_72667[10][10];
  wire [31:0] array_index_72669[10];
  wire [31:0] array_index_72670[10];
  wire [31:0] smul_72674;
  wire [31:0] add_72676;
  wire [31:0] array_update_72678[10];
  wire [31:0] add_72679;
  wire [31:0] array_update_72680[10][10];
  wire [31:0] array_index_72682[10];
  wire [31:0] array_index_72683[10];
  wire [31:0] smul_72687;
  wire [31:0] add_72689;
  wire [31:0] array_update_72690[10];
  wire [31:0] array_update_72691[10][10];
  wire [31:0] array_index_72693[10];
  wire [31:0] add_72695;
  wire [31:0] array_update_72696[10];
  wire [31:0] literal_72697;
  wire [31:0] array_update_72698[10][10];
  wire [31:0] array_index_72700[10];
  wire [31:0] array_index_72701[10];
  wire [31:0] smul_72705;
  wire [31:0] add_72707;
  wire [31:0] array_update_72709[10];
  wire [31:0] add_72710;
  wire [31:0] array_update_72711[10][10];
  wire [31:0] array_index_72713[10];
  wire [31:0] array_index_72714[10];
  wire [31:0] smul_72718;
  wire [31:0] add_72720;
  wire [31:0] array_update_72722[10];
  wire [31:0] add_72723;
  wire [31:0] array_update_72724[10][10];
  wire [31:0] array_index_72726[10];
  wire [31:0] array_index_72727[10];
  wire [31:0] smul_72731;
  wire [31:0] add_72733;
  wire [31:0] array_update_72735[10];
  wire [31:0] add_72736;
  wire [31:0] array_update_72737[10][10];
  wire [31:0] array_index_72739[10];
  wire [31:0] array_index_72740[10];
  wire [31:0] smul_72744;
  wire [31:0] add_72746;
  wire [31:0] array_update_72748[10];
  wire [31:0] add_72749;
  wire [31:0] array_update_72750[10][10];
  wire [31:0] array_index_72752[10];
  wire [31:0] array_index_72753[10];
  wire [31:0] smul_72757;
  wire [31:0] add_72759;
  wire [31:0] array_update_72761[10];
  wire [31:0] add_72762;
  wire [31:0] array_update_72763[10][10];
  wire [31:0] array_index_72765[10];
  wire [31:0] array_index_72766[10];
  wire [31:0] smul_72770;
  wire [31:0] add_72772;
  wire [31:0] array_update_72774[10];
  wire [31:0] add_72775;
  wire [31:0] array_update_72776[10][10];
  wire [31:0] array_index_72778[10];
  wire [31:0] array_index_72779[10];
  wire [31:0] smul_72783;
  wire [31:0] add_72785;
  wire [31:0] array_update_72787[10];
  wire [31:0] add_72788;
  wire [31:0] array_update_72789[10][10];
  wire [31:0] array_index_72791[10];
  wire [31:0] array_index_72792[10];
  wire [31:0] smul_72796;
  wire [31:0] add_72798;
  wire [31:0] array_update_72800[10];
  wire [31:0] add_72801;
  wire [31:0] array_update_72802[10][10];
  wire [31:0] array_index_72804[10];
  wire [31:0] array_index_72805[10];
  wire [31:0] smul_72809;
  wire [31:0] add_72811;
  wire [31:0] array_update_72813[10];
  wire [31:0] add_72814;
  wire [31:0] array_update_72815[10][10];
  wire [31:0] array_index_72817[10];
  wire [31:0] array_index_72818[10];
  wire [31:0] smul_72822;
  wire [31:0] add_72824;
  wire [31:0] array_update_72825[10];
  wire [31:0] array_update_72826[10][10];
  wire [31:0] array_index_72828[10];
  wire [31:0] add_72830;
  wire [31:0] array_update_72831[10];
  wire [31:0] literal_72832;
  wire [31:0] array_update_72833[10][10];
  wire [31:0] array_index_72835[10];
  wire [31:0] array_index_72836[10];
  wire [31:0] smul_72840;
  wire [31:0] add_72842;
  wire [31:0] array_update_72844[10];
  wire [31:0] add_72845;
  wire [31:0] array_update_72846[10][10];
  wire [31:0] array_index_72848[10];
  wire [31:0] array_index_72849[10];
  wire [31:0] smul_72853;
  wire [31:0] add_72855;
  wire [31:0] array_update_72857[10];
  wire [31:0] add_72858;
  wire [31:0] array_update_72859[10][10];
  wire [31:0] array_index_72861[10];
  wire [31:0] array_index_72862[10];
  wire [31:0] smul_72866;
  wire [31:0] add_72868;
  wire [31:0] array_update_72870[10];
  wire [31:0] add_72871;
  wire [31:0] array_update_72872[10][10];
  wire [31:0] array_index_72874[10];
  wire [31:0] array_index_72875[10];
  wire [31:0] smul_72879;
  wire [31:0] add_72881;
  wire [31:0] array_update_72883[10];
  wire [31:0] add_72884;
  wire [31:0] array_update_72885[10][10];
  wire [31:0] array_index_72887[10];
  wire [31:0] array_index_72888[10];
  wire [31:0] smul_72892;
  wire [31:0] add_72894;
  wire [31:0] array_update_72896[10];
  wire [31:0] add_72897;
  wire [31:0] array_update_72898[10][10];
  wire [31:0] array_index_72900[10];
  wire [31:0] array_index_72901[10];
  wire [31:0] smul_72905;
  wire [31:0] add_72907;
  wire [31:0] array_update_72909[10];
  wire [31:0] add_72910;
  wire [31:0] array_update_72911[10][10];
  wire [31:0] array_index_72913[10];
  wire [31:0] array_index_72914[10];
  wire [31:0] smul_72918;
  wire [31:0] add_72920;
  wire [31:0] array_update_72922[10];
  wire [31:0] add_72923;
  wire [31:0] array_update_72924[10][10];
  wire [31:0] array_index_72926[10];
  wire [31:0] array_index_72927[10];
  wire [31:0] smul_72931;
  wire [31:0] add_72933;
  wire [31:0] array_update_72935[10];
  wire [31:0] add_72936;
  wire [31:0] array_update_72937[10][10];
  wire [31:0] array_index_72939[10];
  wire [31:0] array_index_72940[10];
  wire [31:0] smul_72944;
  wire [31:0] add_72946;
  wire [31:0] array_update_72948[10];
  wire [31:0] add_72949;
  wire [31:0] array_update_72950[10][10];
  wire [31:0] array_index_72952[10];
  wire [31:0] array_index_72953[10];
  wire [31:0] smul_72957;
  wire [31:0] add_72959;
  wire [31:0] array_update_72960[10];
  wire [31:0] array_update_72961[10][10];
  wire [31:0] array_index_72963[10];
  wire [31:0] add_72965;
  wire [31:0] array_update_72966[10];
  wire [31:0] literal_72967;
  wire [31:0] array_update_72968[10][10];
  wire [31:0] array_index_72970[10];
  wire [31:0] array_index_72971[10];
  wire [31:0] smul_72975;
  wire [31:0] add_72977;
  wire [31:0] array_update_72979[10];
  wire [31:0] add_72980;
  wire [31:0] array_update_72981[10][10];
  wire [31:0] array_index_72983[10];
  wire [31:0] array_index_72984[10];
  wire [31:0] smul_72988;
  wire [31:0] add_72990;
  wire [31:0] array_update_72992[10];
  wire [31:0] add_72993;
  wire [31:0] array_update_72994[10][10];
  wire [31:0] array_index_72996[10];
  wire [31:0] array_index_72997[10];
  wire [31:0] smul_73001;
  wire [31:0] add_73003;
  wire [31:0] array_update_73005[10];
  wire [31:0] add_73006;
  wire [31:0] array_update_73007[10][10];
  wire [31:0] array_index_73009[10];
  wire [31:0] array_index_73010[10];
  wire [31:0] smul_73014;
  wire [31:0] add_73016;
  wire [31:0] array_update_73018[10];
  wire [31:0] add_73019;
  wire [31:0] array_update_73020[10][10];
  wire [31:0] array_index_73022[10];
  wire [31:0] array_index_73023[10];
  wire [31:0] smul_73027;
  wire [31:0] add_73029;
  wire [31:0] array_update_73031[10];
  wire [31:0] add_73032;
  wire [31:0] array_update_73033[10][10];
  wire [31:0] array_index_73035[10];
  wire [31:0] array_index_73036[10];
  wire [31:0] smul_73040;
  wire [31:0] add_73042;
  wire [31:0] array_update_73044[10];
  wire [31:0] add_73045;
  wire [31:0] array_update_73046[10][10];
  wire [31:0] array_index_73048[10];
  wire [31:0] array_index_73049[10];
  wire [31:0] smul_73053;
  wire [31:0] add_73055;
  wire [31:0] array_update_73057[10];
  wire [31:0] add_73058;
  wire [31:0] array_update_73059[10][10];
  wire [31:0] array_index_73061[10];
  wire [31:0] array_index_73062[10];
  wire [31:0] smul_73066;
  wire [31:0] add_73068;
  wire [31:0] array_update_73070[10];
  wire [31:0] add_73071;
  wire [31:0] array_update_73072[10][10];
  wire [31:0] array_index_73074[10];
  wire [31:0] array_index_73075[10];
  wire [31:0] smul_73079;
  wire [31:0] add_73081;
  wire [31:0] array_update_73083[10];
  wire [31:0] add_73084;
  wire [31:0] array_update_73085[10][10];
  wire [31:0] array_index_73087[10];
  wire [31:0] array_index_73088[10];
  wire [31:0] smul_73092;
  wire [31:0] add_73094;
  wire [31:0] array_update_73095[10];
  wire [31:0] array_update_73096[10][10];
  wire [31:0] array_index_73098[10];
  wire [31:0] add_73100;
  wire [31:0] array_update_73101[10];
  wire [31:0] literal_73102;
  wire [31:0] array_update_73103[10][10];
  wire [31:0] array_index_73105[10];
  wire [31:0] array_index_73106[10];
  wire [31:0] smul_73110;
  wire [31:0] add_73112;
  wire [31:0] array_update_73114[10];
  wire [31:0] add_73115;
  wire [31:0] array_update_73116[10][10];
  wire [31:0] array_index_73118[10];
  wire [31:0] array_index_73119[10];
  wire [31:0] smul_73123;
  wire [31:0] add_73125;
  wire [31:0] array_update_73127[10];
  wire [31:0] add_73128;
  wire [31:0] array_update_73129[10][10];
  wire [31:0] array_index_73131[10];
  wire [31:0] array_index_73132[10];
  wire [31:0] smul_73136;
  wire [31:0] add_73138;
  wire [31:0] array_update_73140[10];
  wire [31:0] add_73141;
  wire [31:0] array_update_73142[10][10];
  wire [31:0] array_index_73144[10];
  wire [31:0] array_index_73145[10];
  wire [31:0] smul_73149;
  wire [31:0] add_73151;
  wire [31:0] array_update_73153[10];
  wire [31:0] add_73154;
  wire [31:0] array_update_73155[10][10];
  wire [31:0] array_index_73157[10];
  wire [31:0] array_index_73158[10];
  wire [31:0] smul_73162;
  wire [31:0] add_73164;
  wire [31:0] array_update_73166[10];
  wire [31:0] add_73167;
  wire [31:0] array_update_73168[10][10];
  wire [31:0] array_index_73170[10];
  wire [31:0] array_index_73171[10];
  wire [31:0] smul_73175;
  wire [31:0] add_73177;
  wire [31:0] array_update_73179[10];
  wire [31:0] add_73180;
  wire [31:0] array_update_73181[10][10];
  wire [31:0] array_index_73183[10];
  wire [31:0] array_index_73184[10];
  wire [31:0] smul_73188;
  wire [31:0] add_73190;
  wire [31:0] array_update_73192[10];
  wire [31:0] add_73193;
  wire [31:0] array_update_73194[10][10];
  wire [31:0] array_index_73196[10];
  wire [31:0] array_index_73197[10];
  wire [31:0] smul_73201;
  wire [31:0] add_73203;
  wire [31:0] array_update_73205[10];
  wire [31:0] add_73206;
  wire [31:0] array_update_73207[10][10];
  wire [31:0] array_index_73209[10];
  wire [31:0] array_index_73210[10];
  wire [31:0] smul_73214;
  wire [31:0] add_73216;
  wire [31:0] array_update_73218[10];
  wire [31:0] add_73219;
  wire [31:0] array_update_73220[10][10];
  wire [31:0] array_index_73222[10];
  wire [31:0] array_index_73223[10];
  wire [31:0] smul_73227;
  wire [31:0] add_73229;
  wire [31:0] array_update_73230[10];
  wire [31:0] array_update_73231[10][10];
  wire [31:0] array_index_73233[10];
  wire [31:0] add_73235;
  wire [31:0] array_update_73236[10];
  wire [31:0] literal_73237;
  wire [31:0] array_update_73238[10][10];
  wire [31:0] array_index_73240[10];
  wire [31:0] array_index_73241[10];
  wire [31:0] smul_73245;
  wire [31:0] add_73247;
  wire [31:0] array_update_73249[10];
  wire [31:0] add_73250;
  wire [31:0] array_update_73251[10][10];
  wire [31:0] array_index_73253[10];
  wire [31:0] array_index_73254[10];
  wire [31:0] smul_73258;
  wire [31:0] add_73260;
  wire [31:0] array_update_73262[10];
  wire [31:0] add_73263;
  wire [31:0] array_update_73264[10][10];
  wire [31:0] array_index_73266[10];
  wire [31:0] array_index_73267[10];
  wire [31:0] smul_73271;
  wire [31:0] add_73273;
  wire [31:0] array_update_73275[10];
  wire [31:0] add_73276;
  wire [31:0] array_update_73277[10][10];
  wire [31:0] array_index_73279[10];
  wire [31:0] array_index_73280[10];
  wire [31:0] smul_73284;
  wire [31:0] add_73286;
  wire [31:0] array_update_73288[10];
  wire [31:0] add_73289;
  wire [31:0] array_update_73290[10][10];
  wire [31:0] array_index_73292[10];
  wire [31:0] array_index_73293[10];
  wire [31:0] smul_73297;
  wire [31:0] add_73299;
  wire [31:0] array_update_73301[10];
  wire [31:0] add_73302;
  wire [31:0] array_update_73303[10][10];
  wire [31:0] array_index_73305[10];
  wire [31:0] array_index_73306[10];
  wire [31:0] smul_73310;
  wire [31:0] add_73312;
  wire [31:0] array_update_73314[10];
  wire [31:0] add_73315;
  wire [31:0] array_update_73316[10][10];
  wire [31:0] array_index_73318[10];
  wire [31:0] array_index_73319[10];
  wire [31:0] smul_73323;
  wire [31:0] add_73325;
  wire [31:0] array_update_73327[10];
  wire [31:0] add_73328;
  wire [31:0] array_update_73329[10][10];
  wire [31:0] array_index_73331[10];
  wire [31:0] array_index_73332[10];
  wire [31:0] smul_73336;
  wire [31:0] add_73338;
  wire [31:0] array_update_73340[10];
  wire [31:0] add_73341;
  wire [31:0] array_update_73342[10][10];
  wire [31:0] array_index_73344[10];
  wire [31:0] array_index_73345[10];
  wire [31:0] smul_73349;
  wire [31:0] add_73351;
  wire [31:0] array_update_73353[10];
  wire [31:0] add_73354;
  wire [31:0] array_update_73355[10][10];
  wire [31:0] array_index_73357[10];
  wire [31:0] array_index_73358[10];
  wire [31:0] smul_73362;
  wire [31:0] add_73364;
  wire [31:0] array_update_73365[10];
  wire [31:0] array_update_73367[10][10];
  wire [31:0] add_73368;
  wire [31:0] array_index_73369[10];
  wire [31:0] literal_73371;
  wire [31:0] array_update_73372[10];
  wire [31:0] literal_73373;
  wire [31:0] array_update_73374[10][10];
  wire [31:0] array_index_73375[10];
  wire [31:0] array_index_73376[10];
  wire [31:0] array_index_73377[10];
  wire [31:0] smul_73381;
  wire [31:0] add_73383;
  wire [31:0] array_update_73385[10];
  wire [31:0] add_73386;
  wire [31:0] array_update_73387[10][10];
  wire [31:0] array_index_73389[10];
  wire [31:0] array_index_73390[10];
  wire [31:0] smul_73394;
  wire [31:0] add_73396;
  wire [31:0] array_update_73398[10];
  wire [31:0] add_73399;
  wire [31:0] array_update_73400[10][10];
  wire [31:0] array_index_73402[10];
  wire [31:0] array_index_73403[10];
  wire [31:0] smul_73407;
  wire [31:0] add_73409;
  wire [31:0] array_update_73411[10];
  wire [31:0] add_73412;
  wire [31:0] array_update_73413[10][10];
  wire [31:0] array_index_73415[10];
  wire [31:0] array_index_73416[10];
  wire [31:0] smul_73420;
  wire [31:0] add_73422;
  wire [31:0] array_update_73424[10];
  wire [31:0] add_73425;
  wire [31:0] array_update_73426[10][10];
  wire [31:0] array_index_73428[10];
  wire [31:0] array_index_73429[10];
  wire [31:0] smul_73433;
  wire [31:0] add_73435;
  wire [31:0] array_update_73437[10];
  wire [31:0] add_73438;
  wire [31:0] array_update_73439[10][10];
  wire [31:0] array_index_73441[10];
  wire [31:0] array_index_73442[10];
  wire [31:0] smul_73446;
  wire [31:0] add_73448;
  wire [31:0] array_update_73450[10];
  wire [31:0] add_73451;
  wire [31:0] array_update_73452[10][10];
  wire [31:0] array_index_73454[10];
  wire [31:0] array_index_73455[10];
  wire [31:0] smul_73459;
  wire [31:0] add_73461;
  wire [31:0] array_update_73463[10];
  wire [31:0] add_73464;
  wire [31:0] array_update_73465[10][10];
  wire [31:0] array_index_73467[10];
  wire [31:0] array_index_73468[10];
  wire [31:0] smul_73472;
  wire [31:0] add_73474;
  wire [31:0] array_update_73476[10];
  wire [31:0] add_73477;
  wire [31:0] array_update_73478[10][10];
  wire [31:0] array_index_73480[10];
  wire [31:0] array_index_73481[10];
  wire [31:0] smul_73485;
  wire [31:0] add_73487;
  wire [31:0] array_update_73489[10];
  wire [31:0] add_73490;
  wire [31:0] array_update_73491[10][10];
  wire [31:0] array_index_73493[10];
  wire [31:0] array_index_73494[10];
  wire [31:0] smul_73498;
  wire [31:0] add_73500;
  wire [31:0] array_update_73501[10];
  wire [31:0] array_update_73502[10][10];
  wire [31:0] array_index_73504[10];
  wire [31:0] add_73506;
  wire [31:0] array_update_73507[10];
  wire [31:0] literal_73508;
  wire [31:0] array_update_73509[10][10];
  wire [31:0] array_index_73511[10];
  wire [31:0] array_index_73512[10];
  wire [31:0] smul_73516;
  wire [31:0] add_73518;
  wire [31:0] array_update_73520[10];
  wire [31:0] add_73521;
  wire [31:0] array_update_73522[10][10];
  wire [31:0] array_index_73524[10];
  wire [31:0] array_index_73525[10];
  wire [31:0] smul_73529;
  wire [31:0] add_73531;
  wire [31:0] array_update_73533[10];
  wire [31:0] add_73534;
  wire [31:0] array_update_73535[10][10];
  wire [31:0] array_index_73537[10];
  wire [31:0] array_index_73538[10];
  wire [31:0] smul_73542;
  wire [31:0] add_73544;
  wire [31:0] array_update_73546[10];
  wire [31:0] add_73547;
  wire [31:0] array_update_73548[10][10];
  wire [31:0] array_index_73550[10];
  wire [31:0] array_index_73551[10];
  wire [31:0] smul_73555;
  wire [31:0] add_73557;
  wire [31:0] array_update_73559[10];
  wire [31:0] add_73560;
  wire [31:0] array_update_73561[10][10];
  wire [31:0] array_index_73563[10];
  wire [31:0] array_index_73564[10];
  wire [31:0] smul_73568;
  wire [31:0] add_73570;
  wire [31:0] array_update_73572[10];
  wire [31:0] add_73573;
  wire [31:0] array_update_73574[10][10];
  wire [31:0] array_index_73576[10];
  wire [31:0] array_index_73577[10];
  wire [31:0] smul_73581;
  wire [31:0] add_73583;
  wire [31:0] array_update_73585[10];
  wire [31:0] add_73586;
  wire [31:0] array_update_73587[10][10];
  wire [31:0] array_index_73589[10];
  wire [31:0] array_index_73590[10];
  wire [31:0] smul_73594;
  wire [31:0] add_73596;
  wire [31:0] array_update_73598[10];
  wire [31:0] add_73599;
  wire [31:0] array_update_73600[10][10];
  wire [31:0] array_index_73602[10];
  wire [31:0] array_index_73603[10];
  wire [31:0] smul_73607;
  wire [31:0] add_73609;
  wire [31:0] array_update_73611[10];
  wire [31:0] add_73612;
  wire [31:0] array_update_73613[10][10];
  wire [31:0] array_index_73615[10];
  wire [31:0] array_index_73616[10];
  wire [31:0] smul_73620;
  wire [31:0] add_73622;
  wire [31:0] array_update_73624[10];
  wire [31:0] add_73625;
  wire [31:0] array_update_73626[10][10];
  wire [31:0] array_index_73628[10];
  wire [31:0] array_index_73629[10];
  wire [31:0] smul_73633;
  wire [31:0] add_73635;
  wire [31:0] array_update_73636[10];
  wire [31:0] array_update_73637[10][10];
  wire [31:0] array_index_73639[10];
  wire [31:0] add_73641;
  wire [31:0] array_update_73642[10];
  wire [31:0] literal_73643;
  wire [31:0] array_update_73644[10][10];
  wire [31:0] array_index_73646[10];
  wire [31:0] array_index_73647[10];
  wire [31:0] smul_73651;
  wire [31:0] add_73653;
  wire [31:0] array_update_73655[10];
  wire [31:0] add_73656;
  wire [31:0] array_update_73657[10][10];
  wire [31:0] array_index_73659[10];
  wire [31:0] array_index_73660[10];
  wire [31:0] smul_73664;
  wire [31:0] add_73666;
  wire [31:0] array_update_73668[10];
  wire [31:0] add_73669;
  wire [31:0] array_update_73670[10][10];
  wire [31:0] array_index_73672[10];
  wire [31:0] array_index_73673[10];
  wire [31:0] smul_73677;
  wire [31:0] add_73679;
  wire [31:0] array_update_73681[10];
  wire [31:0] add_73682;
  wire [31:0] array_update_73683[10][10];
  wire [31:0] array_index_73685[10];
  wire [31:0] array_index_73686[10];
  wire [31:0] smul_73690;
  wire [31:0] add_73692;
  wire [31:0] array_update_73694[10];
  wire [31:0] add_73695;
  wire [31:0] array_update_73696[10][10];
  wire [31:0] array_index_73698[10];
  wire [31:0] array_index_73699[10];
  wire [31:0] smul_73703;
  wire [31:0] add_73705;
  wire [31:0] array_update_73707[10];
  wire [31:0] add_73708;
  wire [31:0] array_update_73709[10][10];
  wire [31:0] array_index_73711[10];
  wire [31:0] array_index_73712[10];
  wire [31:0] smul_73716;
  wire [31:0] add_73718;
  wire [31:0] array_update_73720[10];
  wire [31:0] add_73721;
  wire [31:0] array_update_73722[10][10];
  wire [31:0] array_index_73724[10];
  wire [31:0] array_index_73725[10];
  wire [31:0] smul_73729;
  wire [31:0] add_73731;
  wire [31:0] array_update_73733[10];
  wire [31:0] add_73734;
  wire [31:0] array_update_73735[10][10];
  wire [31:0] array_index_73737[10];
  wire [31:0] array_index_73738[10];
  wire [31:0] smul_73742;
  wire [31:0] add_73744;
  wire [31:0] array_update_73746[10];
  wire [31:0] add_73747;
  wire [31:0] array_update_73748[10][10];
  wire [31:0] array_index_73750[10];
  wire [31:0] array_index_73751[10];
  wire [31:0] smul_73755;
  wire [31:0] add_73757;
  wire [31:0] array_update_73759[10];
  wire [31:0] add_73760;
  wire [31:0] array_update_73761[10][10];
  wire [31:0] array_index_73763[10];
  wire [31:0] array_index_73764[10];
  wire [31:0] smul_73768;
  wire [31:0] add_73770;
  wire [31:0] array_update_73771[10];
  wire [31:0] array_update_73772[10][10];
  wire [31:0] array_index_73774[10];
  wire [31:0] add_73776;
  wire [31:0] array_update_73777[10];
  wire [31:0] literal_73778;
  wire [31:0] array_update_73779[10][10];
  wire [31:0] array_index_73781[10];
  wire [31:0] array_index_73782[10];
  wire [31:0] smul_73786;
  wire [31:0] add_73788;
  wire [31:0] array_update_73790[10];
  wire [31:0] add_73791;
  wire [31:0] array_update_73792[10][10];
  wire [31:0] array_index_73794[10];
  wire [31:0] array_index_73795[10];
  wire [31:0] smul_73799;
  wire [31:0] add_73801;
  wire [31:0] array_update_73803[10];
  wire [31:0] add_73804;
  wire [31:0] array_update_73805[10][10];
  wire [31:0] array_index_73807[10];
  wire [31:0] array_index_73808[10];
  wire [31:0] smul_73812;
  wire [31:0] add_73814;
  wire [31:0] array_update_73816[10];
  wire [31:0] add_73817;
  wire [31:0] array_update_73818[10][10];
  wire [31:0] array_index_73820[10];
  wire [31:0] array_index_73821[10];
  wire [31:0] smul_73825;
  wire [31:0] add_73827;
  wire [31:0] array_update_73829[10];
  wire [31:0] add_73830;
  wire [31:0] array_update_73831[10][10];
  wire [31:0] array_index_73833[10];
  wire [31:0] array_index_73834[10];
  wire [31:0] smul_73838;
  wire [31:0] add_73840;
  wire [31:0] array_update_73842[10];
  wire [31:0] add_73843;
  wire [31:0] array_update_73844[10][10];
  wire [31:0] array_index_73846[10];
  wire [31:0] array_index_73847[10];
  wire [31:0] smul_73851;
  wire [31:0] add_73853;
  wire [31:0] array_update_73855[10];
  wire [31:0] add_73856;
  wire [31:0] array_update_73857[10][10];
  wire [31:0] array_index_73859[10];
  wire [31:0] array_index_73860[10];
  wire [31:0] smul_73864;
  wire [31:0] add_73866;
  wire [31:0] array_update_73868[10];
  wire [31:0] add_73869;
  wire [31:0] array_update_73870[10][10];
  wire [31:0] array_index_73872[10];
  wire [31:0] array_index_73873[10];
  wire [31:0] smul_73877;
  wire [31:0] add_73879;
  wire [31:0] array_update_73881[10];
  wire [31:0] add_73882;
  wire [31:0] array_update_73883[10][10];
  wire [31:0] array_index_73885[10];
  wire [31:0] array_index_73886[10];
  wire [31:0] smul_73890;
  wire [31:0] add_73892;
  wire [31:0] array_update_73894[10];
  wire [31:0] add_73895;
  wire [31:0] array_update_73896[10][10];
  wire [31:0] array_index_73898[10];
  wire [31:0] array_index_73899[10];
  wire [31:0] smul_73903;
  wire [31:0] add_73905;
  wire [31:0] array_update_73906[10];
  wire [31:0] array_update_73907[10][10];
  wire [31:0] array_index_73909[10];
  wire [31:0] add_73911;
  wire [31:0] array_update_73912[10];
  wire [31:0] literal_73913;
  wire [31:0] array_update_73914[10][10];
  wire [31:0] array_index_73916[10];
  wire [31:0] array_index_73917[10];
  wire [31:0] smul_73921;
  wire [31:0] add_73923;
  wire [31:0] array_update_73925[10];
  wire [31:0] add_73926;
  wire [31:0] array_update_73927[10][10];
  wire [31:0] array_index_73929[10];
  wire [31:0] array_index_73930[10];
  wire [31:0] smul_73934;
  wire [31:0] add_73936;
  wire [31:0] array_update_73938[10];
  wire [31:0] add_73939;
  wire [31:0] array_update_73940[10][10];
  wire [31:0] array_index_73942[10];
  wire [31:0] array_index_73943[10];
  wire [31:0] smul_73947;
  wire [31:0] add_73949;
  wire [31:0] array_update_73951[10];
  wire [31:0] add_73952;
  wire [31:0] array_update_73953[10][10];
  wire [31:0] array_index_73955[10];
  wire [31:0] array_index_73956[10];
  wire [31:0] smul_73960;
  wire [31:0] add_73962;
  wire [31:0] array_update_73964[10];
  wire [31:0] add_73965;
  wire [31:0] array_update_73966[10][10];
  wire [31:0] array_index_73968[10];
  wire [31:0] array_index_73969[10];
  wire [31:0] smul_73973;
  wire [31:0] add_73975;
  wire [31:0] array_update_73977[10];
  wire [31:0] add_73978;
  wire [31:0] array_update_73979[10][10];
  wire [31:0] array_index_73981[10];
  wire [31:0] array_index_73982[10];
  wire [31:0] smul_73986;
  wire [31:0] add_73988;
  wire [31:0] array_update_73990[10];
  wire [31:0] add_73991;
  wire [31:0] array_update_73992[10][10];
  wire [31:0] array_index_73994[10];
  wire [31:0] array_index_73995[10];
  wire [31:0] smul_73999;
  wire [31:0] add_74001;
  wire [31:0] array_update_74003[10];
  wire [31:0] add_74004;
  wire [31:0] array_update_74005[10][10];
  wire [31:0] array_index_74007[10];
  wire [31:0] array_index_74008[10];
  wire [31:0] smul_74012;
  wire [31:0] add_74014;
  wire [31:0] array_update_74016[10];
  wire [31:0] add_74017;
  wire [31:0] array_update_74018[10][10];
  wire [31:0] array_index_74020[10];
  wire [31:0] array_index_74021[10];
  wire [31:0] smul_74025;
  wire [31:0] add_74027;
  wire [31:0] array_update_74029[10];
  wire [31:0] add_74030;
  wire [31:0] array_update_74031[10][10];
  wire [31:0] array_index_74033[10];
  wire [31:0] array_index_74034[10];
  wire [31:0] smul_74038;
  wire [31:0] add_74040;
  wire [31:0] array_update_74041[10];
  wire [31:0] array_update_74042[10][10];
  wire [31:0] array_index_74044[10];
  wire [31:0] add_74046;
  wire [31:0] array_update_74047[10];
  wire [31:0] literal_74048;
  wire [31:0] array_update_74049[10][10];
  wire [31:0] array_index_74051[10];
  wire [31:0] array_index_74052[10];
  wire [31:0] smul_74056;
  wire [31:0] add_74058;
  wire [31:0] array_update_74060[10];
  wire [31:0] add_74061;
  wire [31:0] array_update_74062[10][10];
  wire [31:0] array_index_74064[10];
  wire [31:0] array_index_74065[10];
  wire [31:0] smul_74069;
  wire [31:0] add_74071;
  wire [31:0] array_update_74073[10];
  wire [31:0] add_74074;
  wire [31:0] array_update_74075[10][10];
  wire [31:0] array_index_74077[10];
  wire [31:0] array_index_74078[10];
  wire [31:0] smul_74082;
  wire [31:0] add_74084;
  wire [31:0] array_update_74086[10];
  wire [31:0] add_74087;
  wire [31:0] array_update_74088[10][10];
  wire [31:0] array_index_74090[10];
  wire [31:0] array_index_74091[10];
  wire [31:0] smul_74095;
  wire [31:0] add_74097;
  wire [31:0] array_update_74099[10];
  wire [31:0] add_74100;
  wire [31:0] array_update_74101[10][10];
  wire [31:0] array_index_74103[10];
  wire [31:0] array_index_74104[10];
  wire [31:0] smul_74108;
  wire [31:0] add_74110;
  wire [31:0] array_update_74112[10];
  wire [31:0] add_74113;
  wire [31:0] array_update_74114[10][10];
  wire [31:0] array_index_74116[10];
  wire [31:0] array_index_74117[10];
  wire [31:0] smul_74121;
  wire [31:0] add_74123;
  wire [31:0] array_update_74125[10];
  wire [31:0] add_74126;
  wire [31:0] array_update_74127[10][10];
  wire [31:0] array_index_74129[10];
  wire [31:0] array_index_74130[10];
  wire [31:0] smul_74134;
  wire [31:0] add_74136;
  wire [31:0] array_update_74138[10];
  wire [31:0] add_74139;
  wire [31:0] array_update_74140[10][10];
  wire [31:0] array_index_74142[10];
  wire [31:0] array_index_74143[10];
  wire [31:0] smul_74147;
  wire [31:0] add_74149;
  wire [31:0] array_update_74151[10];
  wire [31:0] add_74152;
  wire [31:0] array_update_74153[10][10];
  wire [31:0] array_index_74155[10];
  wire [31:0] array_index_74156[10];
  wire [31:0] smul_74160;
  wire [31:0] add_74162;
  wire [31:0] array_update_74164[10];
  wire [31:0] add_74165;
  wire [31:0] array_update_74166[10][10];
  wire [31:0] array_index_74168[10];
  wire [31:0] array_index_74169[10];
  wire [31:0] smul_74173;
  wire [31:0] add_74175;
  wire [31:0] array_update_74176[10];
  wire [31:0] array_update_74177[10][10];
  wire [31:0] array_index_74179[10];
  wire [31:0] add_74181;
  wire [31:0] array_update_74182[10];
  wire [31:0] literal_74183;
  wire [31:0] array_update_74184[10][10];
  wire [31:0] array_index_74186[10];
  wire [31:0] array_index_74187[10];
  wire [31:0] smul_74191;
  wire [31:0] add_74193;
  wire [31:0] array_update_74195[10];
  wire [31:0] add_74196;
  wire [31:0] array_update_74197[10][10];
  wire [31:0] array_index_74199[10];
  wire [31:0] array_index_74200[10];
  wire [31:0] smul_74204;
  wire [31:0] add_74206;
  wire [31:0] array_update_74208[10];
  wire [31:0] add_74209;
  wire [31:0] array_update_74210[10][10];
  wire [31:0] array_index_74212[10];
  wire [31:0] array_index_74213[10];
  wire [31:0] smul_74217;
  wire [31:0] add_74219;
  wire [31:0] array_update_74221[10];
  wire [31:0] add_74222;
  wire [31:0] array_update_74223[10][10];
  wire [31:0] array_index_74225[10];
  wire [31:0] array_index_74226[10];
  wire [31:0] smul_74230;
  wire [31:0] add_74232;
  wire [31:0] array_update_74234[10];
  wire [31:0] add_74235;
  wire [31:0] array_update_74236[10][10];
  wire [31:0] array_index_74238[10];
  wire [31:0] array_index_74239[10];
  wire [31:0] smul_74243;
  wire [31:0] add_74245;
  wire [31:0] array_update_74247[10];
  wire [31:0] add_74248;
  wire [31:0] array_update_74249[10][10];
  wire [31:0] array_index_74251[10];
  wire [31:0] array_index_74252[10];
  wire [31:0] smul_74256;
  wire [31:0] add_74258;
  wire [31:0] array_update_74260[10];
  wire [31:0] add_74261;
  wire [31:0] array_update_74262[10][10];
  wire [31:0] array_index_74264[10];
  wire [31:0] array_index_74265[10];
  wire [31:0] smul_74269;
  wire [31:0] add_74271;
  wire [31:0] array_update_74273[10];
  wire [31:0] add_74274;
  wire [31:0] array_update_74275[10][10];
  wire [31:0] array_index_74277[10];
  wire [31:0] array_index_74278[10];
  wire [31:0] smul_74282;
  wire [31:0] add_74284;
  wire [31:0] array_update_74286[10];
  wire [31:0] add_74287;
  wire [31:0] array_update_74288[10][10];
  wire [31:0] array_index_74290[10];
  wire [31:0] array_index_74291[10];
  wire [31:0] smul_74295;
  wire [31:0] add_74297;
  wire [31:0] array_update_74299[10];
  wire [31:0] add_74300;
  wire [31:0] array_update_74301[10][10];
  wire [31:0] array_index_74303[10];
  wire [31:0] array_index_74304[10];
  wire [31:0] smul_74308;
  wire [31:0] add_74310;
  wire [31:0] array_update_74311[10];
  wire [31:0] array_update_74312[10][10];
  wire [31:0] array_index_74314[10];
  wire [31:0] add_74316;
  wire [31:0] array_update_74317[10];
  wire [31:0] literal_74318;
  wire [31:0] array_update_74319[10][10];
  wire [31:0] array_index_74321[10];
  wire [31:0] array_index_74322[10];
  wire [31:0] smul_74326;
  wire [31:0] add_74328;
  wire [31:0] array_update_74330[10];
  wire [31:0] add_74331;
  wire [31:0] array_update_74332[10][10];
  wire [31:0] array_index_74334[10];
  wire [31:0] array_index_74335[10];
  wire [31:0] smul_74339;
  wire [31:0] add_74341;
  wire [31:0] array_update_74343[10];
  wire [31:0] add_74344;
  wire [31:0] array_update_74345[10][10];
  wire [31:0] array_index_74347[10];
  wire [31:0] array_index_74348[10];
  wire [31:0] smul_74352;
  wire [31:0] add_74354;
  wire [31:0] array_update_74356[10];
  wire [31:0] add_74357;
  wire [31:0] array_update_74358[10][10];
  wire [31:0] array_index_74360[10];
  wire [31:0] array_index_74361[10];
  wire [31:0] smul_74365;
  wire [31:0] add_74367;
  wire [31:0] array_update_74369[10];
  wire [31:0] add_74370;
  wire [31:0] array_update_74371[10][10];
  wire [31:0] array_index_74373[10];
  wire [31:0] array_index_74374[10];
  wire [31:0] smul_74378;
  wire [31:0] add_74380;
  wire [31:0] array_update_74382[10];
  wire [31:0] add_74383;
  wire [31:0] array_update_74384[10][10];
  wire [31:0] array_index_74386[10];
  wire [31:0] array_index_74387[10];
  wire [31:0] smul_74391;
  wire [31:0] add_74393;
  wire [31:0] array_update_74395[10];
  wire [31:0] add_74396;
  wire [31:0] array_update_74397[10][10];
  wire [31:0] array_index_74399[10];
  wire [31:0] array_index_74400[10];
  wire [31:0] smul_74404;
  wire [31:0] add_74406;
  wire [31:0] array_update_74408[10];
  wire [31:0] add_74409;
  wire [31:0] array_update_74410[10][10];
  wire [31:0] array_index_74412[10];
  wire [31:0] array_index_74413[10];
  wire [31:0] smul_74417;
  wire [31:0] add_74419;
  wire [31:0] array_update_74421[10];
  wire [31:0] add_74422;
  wire [31:0] array_update_74423[10][10];
  wire [31:0] array_index_74425[10];
  wire [31:0] array_index_74426[10];
  wire [31:0] smul_74430;
  wire [31:0] add_74432;
  wire [31:0] array_update_74434[10];
  wire [31:0] add_74435;
  wire [31:0] array_update_74436[10][10];
  wire [31:0] array_index_74438[10];
  wire [31:0] array_index_74439[10];
  wire [31:0] smul_74443;
  wire [31:0] add_74445;
  wire [31:0] array_update_74446[10];
  wire [31:0] array_update_74447[10][10];
  wire [31:0] array_index_74449[10];
  wire [31:0] add_74451;
  wire [31:0] array_update_74452[10];
  wire [31:0] literal_74453;
  wire [31:0] array_update_74454[10][10];
  wire [31:0] array_index_74456[10];
  wire [31:0] array_index_74457[10];
  wire [31:0] smul_74461;
  wire [31:0] add_74463;
  wire [31:0] array_update_74465[10];
  wire [31:0] add_74466;
  wire [31:0] array_update_74467[10][10];
  wire [31:0] array_index_74469[10];
  wire [31:0] array_index_74470[10];
  wire [31:0] smul_74474;
  wire [31:0] add_74476;
  wire [31:0] array_update_74478[10];
  wire [31:0] add_74479;
  wire [31:0] array_update_74480[10][10];
  wire [31:0] array_index_74482[10];
  wire [31:0] array_index_74483[10];
  wire [31:0] smul_74487;
  wire [31:0] add_74489;
  wire [31:0] array_update_74491[10];
  wire [31:0] add_74492;
  wire [31:0] array_update_74493[10][10];
  wire [31:0] array_index_74495[10];
  wire [31:0] array_index_74496[10];
  wire [31:0] smul_74500;
  wire [31:0] add_74502;
  wire [31:0] array_update_74504[10];
  wire [31:0] add_74505;
  wire [31:0] array_update_74506[10][10];
  wire [31:0] array_index_74508[10];
  wire [31:0] array_index_74509[10];
  wire [31:0] smul_74513;
  wire [31:0] add_74515;
  wire [31:0] array_update_74517[10];
  wire [31:0] add_74518;
  wire [31:0] array_update_74519[10][10];
  wire [31:0] array_index_74521[10];
  wire [31:0] array_index_74522[10];
  wire [31:0] smul_74526;
  wire [31:0] add_74528;
  wire [31:0] array_update_74530[10];
  wire [31:0] add_74531;
  wire [31:0] array_update_74532[10][10];
  wire [31:0] array_index_74534[10];
  wire [31:0] array_index_74535[10];
  wire [31:0] smul_74539;
  wire [31:0] add_74541;
  wire [31:0] array_update_74543[10];
  wire [31:0] add_74544;
  wire [31:0] array_update_74545[10][10];
  wire [31:0] array_index_74547[10];
  wire [31:0] array_index_74548[10];
  wire [31:0] smul_74552;
  wire [31:0] add_74554;
  wire [31:0] array_update_74556[10];
  wire [31:0] add_74557;
  wire [31:0] array_update_74558[10][10];
  wire [31:0] array_index_74560[10];
  wire [31:0] array_index_74561[10];
  wire [31:0] smul_74565;
  wire [31:0] add_74567;
  wire [31:0] array_update_74569[10];
  wire [31:0] add_74570;
  wire [31:0] array_update_74571[10][10];
  wire [31:0] array_index_74573[10];
  wire [31:0] array_index_74574[10];
  wire [31:0] smul_74578;
  wire [31:0] add_74580;
  wire [31:0] array_update_74581[10];
  wire [31:0] array_update_74582[10][10];
  wire [31:0] array_index_74584[10];
  wire [31:0] add_74586;
  wire [31:0] array_update_74587[10];
  wire [31:0] literal_74588;
  wire [31:0] array_update_74589[10][10];
  wire [31:0] array_index_74591[10];
  wire [31:0] array_index_74592[10];
  wire [31:0] smul_74596;
  wire [31:0] add_74598;
  wire [31:0] array_update_74600[10];
  wire [31:0] add_74601;
  wire [31:0] array_update_74602[10][10];
  wire [31:0] array_index_74604[10];
  wire [31:0] array_index_74605[10];
  wire [31:0] smul_74609;
  wire [31:0] add_74611;
  wire [31:0] array_update_74613[10];
  wire [31:0] add_74614;
  wire [31:0] array_update_74615[10][10];
  wire [31:0] array_index_74617[10];
  wire [31:0] array_index_74618[10];
  wire [31:0] smul_74622;
  wire [31:0] add_74624;
  wire [31:0] array_update_74626[10];
  wire [31:0] add_74627;
  wire [31:0] array_update_74628[10][10];
  wire [31:0] array_index_74630[10];
  wire [31:0] array_index_74631[10];
  wire [31:0] smul_74635;
  wire [31:0] add_74637;
  wire [31:0] array_update_74639[10];
  wire [31:0] add_74640;
  wire [31:0] array_update_74641[10][10];
  wire [31:0] array_index_74643[10];
  wire [31:0] array_index_74644[10];
  wire [31:0] smul_74648;
  wire [31:0] add_74650;
  wire [31:0] array_update_74652[10];
  wire [31:0] add_74653;
  wire [31:0] array_update_74654[10][10];
  wire [31:0] array_index_74656[10];
  wire [31:0] array_index_74657[10];
  wire [31:0] smul_74661;
  wire [31:0] add_74663;
  wire [31:0] array_update_74665[10];
  wire [31:0] add_74666;
  wire [31:0] array_update_74667[10][10];
  wire [31:0] array_index_74669[10];
  wire [31:0] array_index_74670[10];
  wire [31:0] smul_74674;
  wire [31:0] add_74676;
  wire [31:0] array_update_74678[10];
  wire [31:0] add_74679;
  wire [31:0] array_update_74680[10][10];
  wire [31:0] array_index_74682[10];
  wire [31:0] array_index_74683[10];
  wire [31:0] smul_74687;
  wire [31:0] add_74689;
  wire [31:0] array_update_74691[10];
  wire [31:0] add_74692;
  wire [31:0] array_update_74693[10][10];
  wire [31:0] array_index_74695[10];
  wire [31:0] array_index_74696[10];
  wire [31:0] smul_74700;
  wire [31:0] add_74702;
  wire [31:0] array_update_74704[10];
  wire [31:0] add_74705;
  wire [31:0] array_update_74706[10][10];
  wire [31:0] array_index_74708[10];
  wire [31:0] array_index_74709[10];
  wire [31:0] smul_74713;
  wire [31:0] add_74715;
  wire [31:0] array_update_74716[10];
  wire [31:0] array_update_74718[10][10];
  wire [31:0] add_74719;
  wire [31:0] array_index_74720[10];
  wire [31:0] literal_74722;
  wire [31:0] array_update_74723[10];
  wire [31:0] literal_74724;
  wire [31:0] array_update_74725[10][10];
  wire [31:0] array_index_74726[10];
  wire [31:0] array_index_74727[10];
  wire [31:0] array_index_74728[10];
  wire [31:0] smul_74732;
  wire [31:0] add_74734;
  wire [31:0] array_update_74736[10];
  wire [31:0] add_74737;
  wire [31:0] array_update_74738[10][10];
  wire [31:0] array_index_74740[10];
  wire [31:0] array_index_74741[10];
  wire [31:0] smul_74745;
  wire [31:0] add_74747;
  wire [31:0] array_update_74749[10];
  wire [31:0] add_74750;
  wire [31:0] array_update_74751[10][10];
  wire [31:0] array_index_74753[10];
  wire [31:0] array_index_74754[10];
  wire [31:0] smul_74758;
  wire [31:0] add_74760;
  wire [31:0] array_update_74762[10];
  wire [31:0] add_74763;
  wire [31:0] array_update_74764[10][10];
  wire [31:0] array_index_74766[10];
  wire [31:0] array_index_74767[10];
  wire [31:0] smul_74771;
  wire [31:0] add_74773;
  wire [31:0] array_update_74775[10];
  wire [31:0] add_74776;
  wire [31:0] array_update_74777[10][10];
  wire [31:0] array_index_74779[10];
  wire [31:0] array_index_74780[10];
  wire [31:0] smul_74784;
  wire [31:0] add_74786;
  wire [31:0] array_update_74788[10];
  wire [31:0] add_74789;
  wire [31:0] array_update_74790[10][10];
  wire [31:0] array_index_74792[10];
  wire [31:0] array_index_74793[10];
  wire [31:0] smul_74797;
  wire [31:0] add_74799;
  wire [31:0] array_update_74801[10];
  wire [31:0] add_74802;
  wire [31:0] array_update_74803[10][10];
  wire [31:0] array_index_74805[10];
  wire [31:0] array_index_74806[10];
  wire [31:0] smul_74810;
  wire [31:0] add_74812;
  wire [31:0] array_update_74814[10];
  wire [31:0] add_74815;
  wire [31:0] array_update_74816[10][10];
  wire [31:0] array_index_74818[10];
  wire [31:0] array_index_74819[10];
  wire [31:0] smul_74823;
  wire [31:0] add_74825;
  wire [31:0] array_update_74827[10];
  wire [31:0] add_74828;
  wire [31:0] array_update_74829[10][10];
  wire [31:0] array_index_74831[10];
  wire [31:0] array_index_74832[10];
  wire [31:0] smul_74836;
  wire [31:0] add_74838;
  wire [31:0] array_update_74840[10];
  wire [31:0] add_74841;
  wire [31:0] array_update_74842[10][10];
  wire [31:0] array_index_74844[10];
  wire [31:0] array_index_74845[10];
  wire [31:0] smul_74849;
  wire [31:0] add_74851;
  wire [31:0] array_update_74852[10];
  wire [31:0] array_update_74853[10][10];
  wire [31:0] array_index_74855[10];
  wire [31:0] add_74857;
  wire [31:0] array_update_74858[10];
  wire [31:0] literal_74859;
  wire [31:0] array_update_74860[10][10];
  wire [31:0] array_index_74862[10];
  wire [31:0] array_index_74863[10];
  wire [31:0] smul_74867;
  wire [31:0] add_74869;
  wire [31:0] array_update_74871[10];
  wire [31:0] add_74872;
  wire [31:0] array_update_74873[10][10];
  wire [31:0] array_index_74875[10];
  wire [31:0] array_index_74876[10];
  wire [31:0] smul_74880;
  wire [31:0] add_74882;
  wire [31:0] array_update_74884[10];
  wire [31:0] add_74885;
  wire [31:0] array_update_74886[10][10];
  wire [31:0] array_index_74888[10];
  wire [31:0] array_index_74889[10];
  wire [31:0] smul_74893;
  wire [31:0] add_74895;
  wire [31:0] array_update_74897[10];
  wire [31:0] add_74898;
  wire [31:0] array_update_74899[10][10];
  wire [31:0] array_index_74901[10];
  wire [31:0] array_index_74902[10];
  wire [31:0] smul_74906;
  wire [31:0] add_74908;
  wire [31:0] array_update_74910[10];
  wire [31:0] add_74911;
  wire [31:0] array_update_74912[10][10];
  wire [31:0] array_index_74914[10];
  wire [31:0] array_index_74915[10];
  wire [31:0] smul_74919;
  wire [31:0] add_74921;
  wire [31:0] array_update_74923[10];
  wire [31:0] add_74924;
  wire [31:0] array_update_74925[10][10];
  wire [31:0] array_index_74927[10];
  wire [31:0] array_index_74928[10];
  wire [31:0] smul_74932;
  wire [31:0] add_74934;
  wire [31:0] array_update_74936[10];
  wire [31:0] add_74937;
  wire [31:0] array_update_74938[10][10];
  wire [31:0] array_index_74940[10];
  wire [31:0] array_index_74941[10];
  wire [31:0] smul_74945;
  wire [31:0] add_74947;
  wire [31:0] array_update_74949[10];
  wire [31:0] add_74950;
  wire [31:0] array_update_74951[10][10];
  wire [31:0] array_index_74953[10];
  wire [31:0] array_index_74954[10];
  wire [31:0] smul_74958;
  wire [31:0] add_74960;
  wire [31:0] array_update_74962[10];
  wire [31:0] add_74963;
  wire [31:0] array_update_74964[10][10];
  wire [31:0] array_index_74966[10];
  wire [31:0] array_index_74967[10];
  wire [31:0] smul_74971;
  wire [31:0] add_74973;
  wire [31:0] array_update_74975[10];
  wire [31:0] add_74976;
  wire [31:0] array_update_74977[10][10];
  wire [31:0] array_index_74979[10];
  wire [31:0] array_index_74980[10];
  wire [31:0] smul_74984;
  wire [31:0] add_74986;
  wire [31:0] array_update_74987[10];
  wire [31:0] array_update_74988[10][10];
  wire [31:0] array_index_74990[10];
  wire [31:0] add_74992;
  wire [31:0] array_update_74993[10];
  wire [31:0] literal_74994;
  wire [31:0] array_update_74995[10][10];
  wire [31:0] array_index_74997[10];
  wire [31:0] array_index_74998[10];
  wire [31:0] smul_75002;
  wire [31:0] add_75004;
  wire [31:0] array_update_75006[10];
  wire [31:0] add_75007;
  wire [31:0] array_update_75008[10][10];
  wire [31:0] array_index_75010[10];
  wire [31:0] array_index_75011[10];
  wire [31:0] smul_75015;
  wire [31:0] add_75017;
  wire [31:0] array_update_75019[10];
  wire [31:0] add_75020;
  wire [31:0] array_update_75021[10][10];
  wire [31:0] array_index_75023[10];
  wire [31:0] array_index_75024[10];
  wire [31:0] smul_75028;
  wire [31:0] add_75030;
  wire [31:0] array_update_75032[10];
  wire [31:0] add_75033;
  wire [31:0] array_update_75034[10][10];
  wire [31:0] array_index_75036[10];
  wire [31:0] array_index_75037[10];
  wire [31:0] smul_75041;
  wire [31:0] add_75043;
  wire [31:0] array_update_75045[10];
  wire [31:0] add_75046;
  wire [31:0] array_update_75047[10][10];
  wire [31:0] array_index_75049[10];
  wire [31:0] array_index_75050[10];
  wire [31:0] smul_75054;
  wire [31:0] add_75056;
  wire [31:0] array_update_75058[10];
  wire [31:0] add_75059;
  wire [31:0] array_update_75060[10][10];
  wire [31:0] array_index_75062[10];
  wire [31:0] array_index_75063[10];
  wire [31:0] smul_75067;
  wire [31:0] add_75069;
  wire [31:0] array_update_75071[10];
  wire [31:0] add_75072;
  wire [31:0] array_update_75073[10][10];
  wire [31:0] array_index_75075[10];
  wire [31:0] array_index_75076[10];
  wire [31:0] smul_75080;
  wire [31:0] add_75082;
  wire [31:0] array_update_75084[10];
  wire [31:0] add_75085;
  wire [31:0] array_update_75086[10][10];
  wire [31:0] array_index_75088[10];
  wire [31:0] array_index_75089[10];
  wire [31:0] smul_75093;
  wire [31:0] add_75095;
  wire [31:0] array_update_75097[10];
  wire [31:0] add_75098;
  wire [31:0] array_update_75099[10][10];
  wire [31:0] array_index_75101[10];
  wire [31:0] array_index_75102[10];
  wire [31:0] smul_75106;
  wire [31:0] add_75108;
  wire [31:0] array_update_75110[10];
  wire [31:0] add_75111;
  wire [31:0] array_update_75112[10][10];
  wire [31:0] array_index_75114[10];
  wire [31:0] array_index_75115[10];
  wire [31:0] smul_75119;
  wire [31:0] add_75121;
  wire [31:0] array_update_75122[10];
  wire [31:0] array_update_75123[10][10];
  wire [31:0] array_index_75125[10];
  wire [31:0] add_75127;
  wire [31:0] array_update_75128[10];
  wire [31:0] literal_75129;
  wire [31:0] array_update_75130[10][10];
  wire [31:0] array_index_75132[10];
  wire [31:0] array_index_75133[10];
  wire [31:0] smul_75137;
  wire [31:0] add_75139;
  wire [31:0] array_update_75141[10];
  wire [31:0] add_75142;
  wire [31:0] array_update_75143[10][10];
  wire [31:0] array_index_75145[10];
  wire [31:0] array_index_75146[10];
  wire [31:0] smul_75150;
  wire [31:0] add_75152;
  wire [31:0] array_update_75154[10];
  wire [31:0] add_75155;
  wire [31:0] array_update_75156[10][10];
  wire [31:0] array_index_75158[10];
  wire [31:0] array_index_75159[10];
  wire [31:0] smul_75163;
  wire [31:0] add_75165;
  wire [31:0] array_update_75167[10];
  wire [31:0] add_75168;
  wire [31:0] array_update_75169[10][10];
  wire [31:0] array_index_75171[10];
  wire [31:0] array_index_75172[10];
  wire [31:0] smul_75176;
  wire [31:0] add_75178;
  wire [31:0] array_update_75180[10];
  wire [31:0] add_75181;
  wire [31:0] array_update_75182[10][10];
  wire [31:0] array_index_75184[10];
  wire [31:0] array_index_75185[10];
  wire [31:0] smul_75189;
  wire [31:0] add_75191;
  wire [31:0] array_update_75193[10];
  wire [31:0] add_75194;
  wire [31:0] array_update_75195[10][10];
  wire [31:0] array_index_75197[10];
  wire [31:0] array_index_75198[10];
  wire [31:0] smul_75202;
  wire [31:0] add_75204;
  wire [31:0] array_update_75206[10];
  wire [31:0] add_75207;
  wire [31:0] array_update_75208[10][10];
  wire [31:0] array_index_75210[10];
  wire [31:0] array_index_75211[10];
  wire [31:0] smul_75215;
  wire [31:0] add_75217;
  wire [31:0] array_update_75219[10];
  wire [31:0] add_75220;
  wire [31:0] array_update_75221[10][10];
  wire [31:0] array_index_75223[10];
  wire [31:0] array_index_75224[10];
  wire [31:0] smul_75228;
  wire [31:0] add_75230;
  wire [31:0] array_update_75232[10];
  wire [31:0] add_75233;
  wire [31:0] array_update_75234[10][10];
  wire [31:0] array_index_75236[10];
  wire [31:0] array_index_75237[10];
  wire [31:0] smul_75241;
  wire [31:0] add_75243;
  wire [31:0] array_update_75245[10];
  wire [31:0] add_75246;
  wire [31:0] array_update_75247[10][10];
  wire [31:0] array_index_75249[10];
  wire [31:0] array_index_75250[10];
  wire [31:0] smul_75254;
  wire [31:0] add_75256;
  wire [31:0] array_update_75257[10];
  wire [31:0] array_update_75258[10][10];
  wire [31:0] array_index_75260[10];
  wire [31:0] add_75262;
  wire [31:0] array_update_75263[10];
  wire [31:0] literal_75264;
  wire [31:0] array_update_75265[10][10];
  wire [31:0] array_index_75267[10];
  wire [31:0] array_index_75268[10];
  wire [31:0] smul_75272;
  wire [31:0] add_75274;
  wire [31:0] array_update_75276[10];
  wire [31:0] add_75277;
  wire [31:0] array_update_75278[10][10];
  wire [31:0] array_index_75280[10];
  wire [31:0] array_index_75281[10];
  wire [31:0] smul_75285;
  wire [31:0] add_75287;
  wire [31:0] array_update_75289[10];
  wire [31:0] add_75290;
  wire [31:0] array_update_75291[10][10];
  wire [31:0] array_index_75293[10];
  wire [31:0] array_index_75294[10];
  wire [31:0] smul_75298;
  wire [31:0] add_75300;
  wire [31:0] array_update_75302[10];
  wire [31:0] add_75303;
  wire [31:0] array_update_75304[10][10];
  wire [31:0] array_index_75306[10];
  wire [31:0] array_index_75307[10];
  wire [31:0] smul_75311;
  wire [31:0] add_75313;
  wire [31:0] array_update_75315[10];
  wire [31:0] add_75316;
  wire [31:0] array_update_75317[10][10];
  wire [31:0] array_index_75319[10];
  wire [31:0] array_index_75320[10];
  wire [31:0] smul_75324;
  wire [31:0] add_75326;
  wire [31:0] array_update_75328[10];
  wire [31:0] add_75329;
  wire [31:0] array_update_75330[10][10];
  wire [31:0] array_index_75332[10];
  wire [31:0] array_index_75333[10];
  wire [31:0] smul_75337;
  wire [31:0] add_75339;
  wire [31:0] array_update_75341[10];
  wire [31:0] add_75342;
  wire [31:0] array_update_75343[10][10];
  wire [31:0] array_index_75345[10];
  wire [31:0] array_index_75346[10];
  wire [31:0] smul_75350;
  wire [31:0] add_75352;
  wire [31:0] array_update_75354[10];
  wire [31:0] add_75355;
  wire [31:0] array_update_75356[10][10];
  wire [31:0] array_index_75358[10];
  wire [31:0] array_index_75359[10];
  wire [31:0] smul_75363;
  wire [31:0] add_75365;
  wire [31:0] array_update_75367[10];
  wire [31:0] add_75368;
  wire [31:0] array_update_75369[10][10];
  wire [31:0] array_index_75371[10];
  wire [31:0] array_index_75372[10];
  wire [31:0] smul_75376;
  wire [31:0] add_75378;
  wire [31:0] array_update_75380[10];
  wire [31:0] add_75381;
  wire [31:0] array_update_75382[10][10];
  wire [31:0] array_index_75384[10];
  wire [31:0] array_index_75385[10];
  wire [31:0] smul_75389;
  wire [31:0] add_75391;
  wire [31:0] array_update_75392[10];
  wire [31:0] array_update_75393[10][10];
  wire [31:0] array_index_75395[10];
  wire [31:0] add_75397;
  wire [31:0] array_update_75398[10];
  wire [31:0] literal_75399;
  wire [31:0] array_update_75400[10][10];
  wire [31:0] array_index_75402[10];
  wire [31:0] array_index_75403[10];
  wire [31:0] smul_75407;
  wire [31:0] add_75409;
  wire [31:0] array_update_75411[10];
  wire [31:0] add_75412;
  wire [31:0] array_update_75413[10][10];
  wire [31:0] array_index_75415[10];
  wire [31:0] array_index_75416[10];
  wire [31:0] smul_75420;
  wire [31:0] add_75422;
  wire [31:0] array_update_75424[10];
  wire [31:0] add_75425;
  wire [31:0] array_update_75426[10][10];
  wire [31:0] array_index_75428[10];
  wire [31:0] array_index_75429[10];
  wire [31:0] smul_75433;
  wire [31:0] add_75435;
  wire [31:0] array_update_75437[10];
  wire [31:0] add_75438;
  wire [31:0] array_update_75439[10][10];
  wire [31:0] array_index_75441[10];
  wire [31:0] array_index_75442[10];
  wire [31:0] smul_75446;
  wire [31:0] add_75448;
  wire [31:0] array_update_75450[10];
  wire [31:0] add_75451;
  wire [31:0] array_update_75452[10][10];
  wire [31:0] array_index_75454[10];
  wire [31:0] array_index_75455[10];
  wire [31:0] smul_75459;
  wire [31:0] add_75461;
  wire [31:0] array_update_75463[10];
  wire [31:0] add_75464;
  wire [31:0] array_update_75465[10][10];
  wire [31:0] array_index_75467[10];
  wire [31:0] array_index_75468[10];
  wire [31:0] smul_75472;
  wire [31:0] add_75474;
  wire [31:0] array_update_75476[10];
  wire [31:0] add_75477;
  wire [31:0] array_update_75478[10][10];
  wire [31:0] array_index_75480[10];
  wire [31:0] array_index_75481[10];
  wire [31:0] smul_75485;
  wire [31:0] add_75487;
  wire [31:0] array_update_75489[10];
  wire [31:0] add_75490;
  wire [31:0] array_update_75491[10][10];
  wire [31:0] array_index_75493[10];
  wire [31:0] array_index_75494[10];
  wire [31:0] smul_75498;
  wire [31:0] add_75500;
  wire [31:0] array_update_75502[10];
  wire [31:0] add_75503;
  wire [31:0] array_update_75504[10][10];
  wire [31:0] array_index_75506[10];
  wire [31:0] array_index_75507[10];
  wire [31:0] smul_75511;
  wire [31:0] add_75513;
  wire [31:0] array_update_75515[10];
  wire [31:0] add_75516;
  wire [31:0] array_update_75517[10][10];
  wire [31:0] array_index_75519[10];
  wire [31:0] array_index_75520[10];
  wire [31:0] smul_75524;
  wire [31:0] add_75526;
  wire [31:0] array_update_75527[10];
  wire [31:0] array_update_75528[10][10];
  wire [31:0] array_index_75530[10];
  wire [31:0] add_75532;
  wire [31:0] array_update_75533[10];
  wire [31:0] literal_75534;
  wire [31:0] array_update_75535[10][10];
  wire [31:0] array_index_75537[10];
  wire [31:0] array_index_75538[10];
  wire [31:0] smul_75542;
  wire [31:0] add_75544;
  wire [31:0] array_update_75546[10];
  wire [31:0] add_75547;
  wire [31:0] array_update_75548[10][10];
  wire [31:0] array_index_75550[10];
  wire [31:0] array_index_75551[10];
  wire [31:0] smul_75555;
  wire [31:0] add_75557;
  wire [31:0] array_update_75559[10];
  wire [31:0] add_75560;
  wire [31:0] array_update_75561[10][10];
  wire [31:0] array_index_75563[10];
  wire [31:0] array_index_75564[10];
  wire [31:0] smul_75568;
  wire [31:0] add_75570;
  wire [31:0] array_update_75572[10];
  wire [31:0] add_75573;
  wire [31:0] array_update_75574[10][10];
  wire [31:0] array_index_75576[10];
  wire [31:0] array_index_75577[10];
  wire [31:0] smul_75581;
  wire [31:0] add_75583;
  wire [31:0] array_update_75585[10];
  wire [31:0] add_75586;
  wire [31:0] array_update_75587[10][10];
  wire [31:0] array_index_75589[10];
  wire [31:0] array_index_75590[10];
  wire [31:0] smul_75594;
  wire [31:0] add_75596;
  wire [31:0] array_update_75598[10];
  wire [31:0] add_75599;
  wire [31:0] array_update_75600[10][10];
  wire [31:0] array_index_75602[10];
  wire [31:0] array_index_75603[10];
  wire [31:0] smul_75607;
  wire [31:0] add_75609;
  wire [31:0] array_update_75611[10];
  wire [31:0] add_75612;
  wire [31:0] array_update_75613[10][10];
  wire [31:0] array_index_75615[10];
  wire [31:0] array_index_75616[10];
  wire [31:0] smul_75620;
  wire [31:0] add_75622;
  wire [31:0] array_update_75624[10];
  wire [31:0] add_75625;
  wire [31:0] array_update_75626[10][10];
  wire [31:0] array_index_75628[10];
  wire [31:0] array_index_75629[10];
  wire [31:0] smul_75633;
  wire [31:0] add_75635;
  wire [31:0] array_update_75637[10];
  wire [31:0] add_75638;
  wire [31:0] array_update_75639[10][10];
  wire [31:0] array_index_75641[10];
  wire [31:0] array_index_75642[10];
  wire [31:0] smul_75646;
  wire [31:0] add_75648;
  wire [31:0] array_update_75650[10];
  wire [31:0] add_75651;
  wire [31:0] array_update_75652[10][10];
  wire [31:0] array_index_75654[10];
  wire [31:0] array_index_75655[10];
  wire [31:0] smul_75659;
  wire [31:0] add_75661;
  wire [31:0] array_update_75662[10];
  wire [31:0] array_update_75663[10][10];
  wire [31:0] array_index_75665[10];
  wire [31:0] add_75667;
  wire [31:0] array_update_75668[10];
  wire [31:0] literal_75669;
  wire [31:0] array_update_75670[10][10];
  wire [31:0] array_index_75672[10];
  wire [31:0] array_index_75673[10];
  wire [31:0] smul_75677;
  wire [31:0] add_75679;
  wire [31:0] array_update_75681[10];
  wire [31:0] add_75682;
  wire [31:0] array_update_75683[10][10];
  wire [31:0] array_index_75685[10];
  wire [31:0] array_index_75686[10];
  wire [31:0] smul_75690;
  wire [31:0] add_75692;
  wire [31:0] array_update_75694[10];
  wire [31:0] add_75695;
  wire [31:0] array_update_75696[10][10];
  wire [31:0] array_index_75698[10];
  wire [31:0] array_index_75699[10];
  wire [31:0] smul_75703;
  wire [31:0] add_75705;
  wire [31:0] array_update_75707[10];
  wire [31:0] add_75708;
  wire [31:0] array_update_75709[10][10];
  wire [31:0] array_index_75711[10];
  wire [31:0] array_index_75712[10];
  wire [31:0] smul_75716;
  wire [31:0] add_75718;
  wire [31:0] array_update_75720[10];
  wire [31:0] add_75721;
  wire [31:0] array_update_75722[10][10];
  wire [31:0] array_index_75724[10];
  wire [31:0] array_index_75725[10];
  wire [31:0] smul_75729;
  wire [31:0] add_75731;
  wire [31:0] array_update_75733[10];
  wire [31:0] add_75734;
  wire [31:0] array_update_75735[10][10];
  wire [31:0] array_index_75737[10];
  wire [31:0] array_index_75738[10];
  wire [31:0] smul_75742;
  wire [31:0] add_75744;
  wire [31:0] array_update_75746[10];
  wire [31:0] add_75747;
  wire [31:0] array_update_75748[10][10];
  wire [31:0] array_index_75750[10];
  wire [31:0] array_index_75751[10];
  wire [31:0] smul_75755;
  wire [31:0] add_75757;
  wire [31:0] array_update_75759[10];
  wire [31:0] add_75760;
  wire [31:0] array_update_75761[10][10];
  wire [31:0] array_index_75763[10];
  wire [31:0] array_index_75764[10];
  wire [31:0] smul_75768;
  wire [31:0] add_75770;
  wire [31:0] array_update_75772[10];
  wire [31:0] add_75773;
  wire [31:0] array_update_75774[10][10];
  wire [31:0] array_index_75776[10];
  wire [31:0] array_index_75777[10];
  wire [31:0] smul_75781;
  wire [31:0] add_75783;
  wire [31:0] array_update_75785[10];
  wire [31:0] add_75786;
  wire [31:0] array_update_75787[10][10];
  wire [31:0] array_index_75789[10];
  wire [31:0] array_index_75790[10];
  wire [31:0] smul_75794;
  wire [31:0] add_75796;
  wire [31:0] array_update_75797[10];
  wire [31:0] array_update_75798[10][10];
  wire [31:0] array_index_75800[10];
  wire [31:0] add_75802;
  wire [31:0] array_update_75803[10];
  wire [31:0] literal_75804;
  wire [31:0] array_update_75805[10][10];
  wire [31:0] array_index_75807[10];
  wire [31:0] array_index_75808[10];
  wire [31:0] smul_75812;
  wire [31:0] add_75814;
  wire [31:0] array_update_75816[10];
  wire [31:0] add_75817;
  wire [31:0] array_update_75818[10][10];
  wire [31:0] array_index_75820[10];
  wire [31:0] array_index_75821[10];
  wire [31:0] smul_75825;
  wire [31:0] add_75827;
  wire [31:0] array_update_75829[10];
  wire [31:0] add_75830;
  wire [31:0] array_update_75831[10][10];
  wire [31:0] array_index_75833[10];
  wire [31:0] array_index_75834[10];
  wire [31:0] smul_75838;
  wire [31:0] add_75840;
  wire [31:0] array_update_75842[10];
  wire [31:0] add_75843;
  wire [31:0] array_update_75844[10][10];
  wire [31:0] array_index_75846[10];
  wire [31:0] array_index_75847[10];
  wire [31:0] smul_75851;
  wire [31:0] add_75853;
  wire [31:0] array_update_75855[10];
  wire [31:0] add_75856;
  wire [31:0] array_update_75857[10][10];
  wire [31:0] array_index_75859[10];
  wire [31:0] array_index_75860[10];
  wire [31:0] smul_75864;
  wire [31:0] add_75866;
  wire [31:0] array_update_75868[10];
  wire [31:0] add_75869;
  wire [31:0] array_update_75870[10][10];
  wire [31:0] array_index_75872[10];
  wire [31:0] array_index_75873[10];
  wire [31:0] smul_75877;
  wire [31:0] add_75879;
  wire [31:0] array_update_75881[10];
  wire [31:0] add_75882;
  wire [31:0] array_update_75883[10][10];
  wire [31:0] array_index_75885[10];
  wire [31:0] array_index_75886[10];
  wire [31:0] smul_75890;
  wire [31:0] add_75892;
  wire [31:0] array_update_75894[10];
  wire [31:0] add_75895;
  wire [31:0] array_update_75896[10][10];
  wire [31:0] array_index_75898[10];
  wire [31:0] array_index_75899[10];
  wire [31:0] smul_75903;
  wire [31:0] add_75905;
  wire [31:0] array_update_75907[10];
  wire [31:0] add_75908;
  wire [31:0] array_update_75909[10][10];
  wire [31:0] array_index_75911[10];
  wire [31:0] array_index_75912[10];
  wire [31:0] smul_75916;
  wire [31:0] add_75918;
  wire [31:0] array_update_75920[10];
  wire [31:0] add_75921;
  wire [31:0] array_update_75922[10][10];
  wire [31:0] array_index_75924[10];
  wire [31:0] array_index_75925[10];
  wire [31:0] smul_75929;
  wire [31:0] add_75931;
  wire [31:0] array_update_75932[10];
  wire [31:0] array_update_75933[10][10];
  wire [31:0] array_index_75935[10];
  wire [31:0] add_75937;
  wire [31:0] array_update_75938[10];
  wire [31:0] literal_75939;
  wire [31:0] array_update_75940[10][10];
  wire [31:0] array_index_75942[10];
  wire [31:0] array_index_75943[10];
  wire [31:0] smul_75947;
  wire [31:0] add_75949;
  wire [31:0] array_update_75951[10];
  wire [31:0] add_75952;
  wire [31:0] array_update_75953[10][10];
  wire [31:0] array_index_75955[10];
  wire [31:0] array_index_75956[10];
  wire [31:0] smul_75960;
  wire [31:0] add_75962;
  wire [31:0] array_update_75964[10];
  wire [31:0] add_75965;
  wire [31:0] array_update_75966[10][10];
  wire [31:0] array_index_75968[10];
  wire [31:0] array_index_75969[10];
  wire [31:0] smul_75973;
  wire [31:0] add_75975;
  wire [31:0] array_update_75977[10];
  wire [31:0] add_75978;
  wire [31:0] array_update_75979[10][10];
  wire [31:0] array_index_75981[10];
  wire [31:0] array_index_75982[10];
  wire [31:0] smul_75986;
  wire [31:0] add_75988;
  wire [31:0] array_update_75990[10];
  wire [31:0] add_75991;
  wire [31:0] array_update_75992[10][10];
  wire [31:0] array_index_75994[10];
  wire [31:0] array_index_75995[10];
  wire [31:0] smul_75999;
  wire [31:0] add_76001;
  wire [31:0] array_update_76003[10];
  wire [31:0] add_76004;
  wire [31:0] array_update_76005[10][10];
  wire [31:0] array_index_76007[10];
  wire [31:0] array_index_76008[10];
  wire [31:0] smul_76012;
  wire [31:0] add_76014;
  wire [31:0] array_update_76016[10];
  wire [31:0] add_76017;
  wire [31:0] array_update_76018[10][10];
  wire [31:0] array_index_76020[10];
  wire [31:0] array_index_76021[10];
  wire [31:0] smul_76025;
  wire [31:0] add_76027;
  wire [31:0] array_update_76029[10];
  wire [31:0] add_76030;
  wire [31:0] array_update_76031[10][10];
  wire [31:0] array_index_76033[10];
  wire [31:0] array_index_76034[10];
  wire [31:0] smul_76038;
  wire [31:0] add_76040;
  wire [31:0] array_update_76042[10];
  wire [31:0] add_76043;
  wire [31:0] array_update_76044[10][10];
  wire [31:0] array_index_76046[10];
  wire [31:0] array_index_76047[10];
  wire [31:0] smul_76051;
  wire [31:0] add_76053;
  wire [31:0] array_update_76055[10];
  wire [31:0] add_76056;
  wire [31:0] array_update_76057[10][10];
  wire [31:0] array_index_76059[10];
  wire [31:0] array_index_76060[10];
  wire [31:0] smul_76064;
  wire [31:0] add_76066;
  wire [31:0] array_update_76067[10];
  wire [31:0] array_update_76069[10][10];
  wire [31:0] add_76070;
  wire [31:0] array_index_76071[10];
  wire [31:0] literal_76073;
  wire [31:0] array_update_76074[10];
  wire [31:0] literal_76075;
  wire [31:0] array_update_76076[10][10];
  wire [31:0] array_index_76077[10];
  wire [31:0] array_index_76078[10];
  wire [31:0] array_index_76079[10];
  wire [31:0] smul_76083;
  wire [31:0] add_76085;
  wire [31:0] array_update_76087[10];
  wire [31:0] add_76088;
  wire [31:0] array_update_76089[10][10];
  wire [31:0] array_index_76091[10];
  wire [31:0] array_index_76092[10];
  wire [31:0] smul_76096;
  wire [31:0] add_76098;
  wire [31:0] array_update_76100[10];
  wire [31:0] add_76101;
  wire [31:0] array_update_76102[10][10];
  wire [31:0] array_index_76104[10];
  wire [31:0] array_index_76105[10];
  wire [31:0] smul_76109;
  wire [31:0] add_76111;
  wire [31:0] array_update_76113[10];
  wire [31:0] add_76114;
  wire [31:0] array_update_76115[10][10];
  wire [31:0] array_index_76117[10];
  wire [31:0] array_index_76118[10];
  wire [31:0] smul_76122;
  wire [31:0] add_76124;
  wire [31:0] array_update_76126[10];
  wire [31:0] add_76127;
  wire [31:0] array_update_76128[10][10];
  wire [31:0] array_index_76130[10];
  wire [31:0] array_index_76131[10];
  wire [31:0] smul_76135;
  wire [31:0] add_76137;
  wire [31:0] array_update_76139[10];
  wire [31:0] add_76140;
  wire [31:0] array_update_76141[10][10];
  wire [31:0] array_index_76143[10];
  wire [31:0] array_index_76144[10];
  wire [31:0] smul_76148;
  wire [31:0] add_76150;
  wire [31:0] array_update_76152[10];
  wire [31:0] add_76153;
  wire [31:0] array_update_76154[10][10];
  wire [31:0] array_index_76156[10];
  wire [31:0] array_index_76157[10];
  wire [31:0] smul_76161;
  wire [31:0] add_76163;
  wire [31:0] array_update_76165[10];
  wire [31:0] add_76166;
  wire [31:0] array_update_76167[10][10];
  wire [31:0] array_index_76169[10];
  wire [31:0] array_index_76170[10];
  wire [31:0] smul_76174;
  wire [31:0] add_76176;
  wire [31:0] array_update_76178[10];
  wire [31:0] add_76179;
  wire [31:0] array_update_76180[10][10];
  wire [31:0] array_index_76182[10];
  wire [31:0] array_index_76183[10];
  wire [31:0] smul_76187;
  wire [31:0] add_76189;
  wire [31:0] array_update_76191[10];
  wire [31:0] add_76192;
  wire [31:0] array_update_76193[10][10];
  wire [31:0] array_index_76195[10];
  wire [31:0] array_index_76196[10];
  wire [31:0] smul_76200;
  wire [31:0] add_76202;
  wire [31:0] array_update_76203[10];
  wire [31:0] array_update_76204[10][10];
  wire [31:0] array_index_76206[10];
  wire [31:0] add_76208;
  wire [31:0] array_update_76209[10];
  wire [31:0] literal_76210;
  wire [31:0] array_update_76211[10][10];
  wire [31:0] array_index_76213[10];
  wire [31:0] array_index_76214[10];
  wire [31:0] smul_76218;
  wire [31:0] add_76220;
  wire [31:0] array_update_76222[10];
  wire [31:0] add_76223;
  wire [31:0] array_update_76224[10][10];
  wire [31:0] array_index_76226[10];
  wire [31:0] array_index_76227[10];
  wire [31:0] smul_76231;
  wire [31:0] add_76233;
  wire [31:0] array_update_76235[10];
  wire [31:0] add_76236;
  wire [31:0] array_update_76237[10][10];
  wire [31:0] array_index_76239[10];
  wire [31:0] array_index_76240[10];
  wire [31:0] smul_76244;
  wire [31:0] add_76246;
  wire [31:0] array_update_76248[10];
  wire [31:0] add_76249;
  wire [31:0] array_update_76250[10][10];
  wire [31:0] array_index_76252[10];
  wire [31:0] array_index_76253[10];
  wire [31:0] smul_76257;
  wire [31:0] add_76259;
  wire [31:0] array_update_76261[10];
  wire [31:0] add_76262;
  wire [31:0] array_update_76263[10][10];
  wire [31:0] array_index_76265[10];
  wire [31:0] array_index_76266[10];
  wire [31:0] smul_76270;
  wire [31:0] add_76272;
  wire [31:0] array_update_76274[10];
  wire [31:0] add_76275;
  wire [31:0] array_update_76276[10][10];
  wire [31:0] array_index_76278[10];
  wire [31:0] array_index_76279[10];
  wire [31:0] smul_76283;
  wire [31:0] add_76285;
  wire [31:0] array_update_76287[10];
  wire [31:0] add_76288;
  wire [31:0] array_update_76289[10][10];
  wire [31:0] array_index_76291[10];
  wire [31:0] array_index_76292[10];
  wire [31:0] smul_76296;
  wire [31:0] add_76298;
  wire [31:0] array_update_76300[10];
  wire [31:0] add_76301;
  wire [31:0] array_update_76302[10][10];
  wire [31:0] array_index_76304[10];
  wire [31:0] array_index_76305[10];
  wire [31:0] smul_76309;
  wire [31:0] add_76311;
  wire [31:0] array_update_76313[10];
  wire [31:0] add_76314;
  wire [31:0] array_update_76315[10][10];
  wire [31:0] array_index_76317[10];
  wire [31:0] array_index_76318[10];
  wire [31:0] smul_76322;
  wire [31:0] add_76324;
  wire [31:0] array_update_76326[10];
  wire [31:0] add_76327;
  wire [31:0] array_update_76328[10][10];
  wire [31:0] array_index_76330[10];
  wire [31:0] array_index_76331[10];
  wire [31:0] smul_76335;
  wire [31:0] add_76337;
  wire [31:0] array_update_76338[10];
  wire [31:0] array_update_76339[10][10];
  wire [31:0] array_index_76341[10];
  wire [31:0] add_76343;
  wire [31:0] array_update_76344[10];
  wire [31:0] literal_76345;
  wire [31:0] array_update_76346[10][10];
  wire [31:0] array_index_76348[10];
  wire [31:0] array_index_76349[10];
  wire [31:0] smul_76353;
  wire [31:0] add_76355;
  wire [31:0] array_update_76357[10];
  wire [31:0] add_76358;
  wire [31:0] array_update_76359[10][10];
  wire [31:0] array_index_76361[10];
  wire [31:0] array_index_76362[10];
  wire [31:0] smul_76366;
  wire [31:0] add_76368;
  wire [31:0] array_update_76370[10];
  wire [31:0] add_76371;
  wire [31:0] array_update_76372[10][10];
  wire [31:0] array_index_76374[10];
  wire [31:0] array_index_76375[10];
  wire [31:0] smul_76379;
  wire [31:0] add_76381;
  wire [31:0] array_update_76383[10];
  wire [31:0] add_76384;
  wire [31:0] array_update_76385[10][10];
  wire [31:0] array_index_76387[10];
  wire [31:0] array_index_76388[10];
  wire [31:0] smul_76392;
  wire [31:0] add_76394;
  wire [31:0] array_update_76396[10];
  wire [31:0] add_76397;
  wire [31:0] array_update_76398[10][10];
  wire [31:0] array_index_76400[10];
  wire [31:0] array_index_76401[10];
  wire [31:0] smul_76405;
  wire [31:0] add_76407;
  wire [31:0] array_update_76409[10];
  wire [31:0] add_76410;
  wire [31:0] array_update_76411[10][10];
  wire [31:0] array_index_76413[10];
  wire [31:0] array_index_76414[10];
  wire [31:0] smul_76418;
  wire [31:0] add_76420;
  wire [31:0] array_update_76422[10];
  wire [31:0] add_76423;
  wire [31:0] array_update_76424[10][10];
  wire [31:0] array_index_76426[10];
  wire [31:0] array_index_76427[10];
  wire [31:0] smul_76431;
  wire [31:0] add_76433;
  wire [31:0] array_update_76435[10];
  wire [31:0] add_76436;
  wire [31:0] array_update_76437[10][10];
  wire [31:0] array_index_76439[10];
  wire [31:0] array_index_76440[10];
  wire [31:0] smul_76444;
  wire [31:0] add_76446;
  wire [31:0] array_update_76448[10];
  wire [31:0] add_76449;
  wire [31:0] array_update_76450[10][10];
  wire [31:0] array_index_76452[10];
  wire [31:0] array_index_76453[10];
  wire [31:0] smul_76457;
  wire [31:0] add_76459;
  wire [31:0] array_update_76461[10];
  wire [31:0] add_76462;
  wire [31:0] array_update_76463[10][10];
  wire [31:0] array_index_76465[10];
  wire [31:0] array_index_76466[10];
  wire [31:0] smul_76470;
  wire [31:0] add_76472;
  wire [31:0] array_update_76473[10];
  wire [31:0] array_update_76474[10][10];
  wire [31:0] array_index_76476[10];
  wire [31:0] add_76478;
  wire [31:0] array_update_76479[10];
  wire [31:0] literal_76480;
  wire [31:0] array_update_76481[10][10];
  wire [31:0] array_index_76483[10];
  wire [31:0] array_index_76484[10];
  wire [31:0] smul_76488;
  wire [31:0] add_76490;
  wire [31:0] array_update_76492[10];
  wire [31:0] add_76493;
  wire [31:0] array_update_76494[10][10];
  wire [31:0] array_index_76496[10];
  wire [31:0] array_index_76497[10];
  wire [31:0] smul_76501;
  wire [31:0] add_76503;
  wire [31:0] array_update_76505[10];
  wire [31:0] add_76506;
  wire [31:0] array_update_76507[10][10];
  wire [31:0] array_index_76509[10];
  wire [31:0] array_index_76510[10];
  wire [31:0] smul_76514;
  wire [31:0] add_76516;
  wire [31:0] array_update_76518[10];
  wire [31:0] add_76519;
  wire [31:0] array_update_76520[10][10];
  wire [31:0] array_index_76522[10];
  wire [31:0] array_index_76523[10];
  wire [31:0] smul_76527;
  wire [31:0] add_76529;
  wire [31:0] array_update_76531[10];
  wire [31:0] add_76532;
  wire [31:0] array_update_76533[10][10];
  wire [31:0] array_index_76535[10];
  wire [31:0] array_index_76536[10];
  wire [31:0] smul_76540;
  wire [31:0] add_76542;
  wire [31:0] array_update_76544[10];
  wire [31:0] add_76545;
  wire [31:0] array_update_76546[10][10];
  wire [31:0] array_index_76548[10];
  wire [31:0] array_index_76549[10];
  wire [31:0] smul_76553;
  wire [31:0] add_76555;
  wire [31:0] array_update_76557[10];
  wire [31:0] add_76558;
  wire [31:0] array_update_76559[10][10];
  wire [31:0] array_index_76561[10];
  wire [31:0] array_index_76562[10];
  wire [31:0] smul_76566;
  wire [31:0] add_76568;
  wire [31:0] array_update_76570[10];
  wire [31:0] add_76571;
  wire [31:0] array_update_76572[10][10];
  wire [31:0] array_index_76574[10];
  wire [31:0] array_index_76575[10];
  wire [31:0] smul_76579;
  wire [31:0] add_76581;
  wire [31:0] array_update_76583[10];
  wire [31:0] add_76584;
  wire [31:0] array_update_76585[10][10];
  wire [31:0] array_index_76587[10];
  wire [31:0] array_index_76588[10];
  wire [31:0] smul_76592;
  wire [31:0] add_76594;
  wire [31:0] array_update_76596[10];
  wire [31:0] add_76597;
  wire [31:0] array_update_76598[10][10];
  wire [31:0] array_index_76600[10];
  wire [31:0] array_index_76601[10];
  wire [31:0] smul_76605;
  wire [31:0] add_76607;
  wire [31:0] array_update_76608[10];
  wire [31:0] array_update_76609[10][10];
  wire [31:0] array_index_76611[10];
  wire [31:0] add_76613;
  wire [31:0] array_update_76614[10];
  wire [31:0] literal_76615;
  wire [31:0] array_update_76616[10][10];
  wire [31:0] array_index_76618[10];
  wire [31:0] array_index_76619[10];
  wire [31:0] smul_76623;
  wire [31:0] add_76625;
  wire [31:0] array_update_76627[10];
  wire [31:0] add_76628;
  wire [31:0] array_update_76629[10][10];
  wire [31:0] array_index_76631[10];
  wire [31:0] array_index_76632[10];
  wire [31:0] smul_76636;
  wire [31:0] add_76638;
  wire [31:0] array_update_76640[10];
  wire [31:0] add_76641;
  wire [31:0] array_update_76642[10][10];
  wire [31:0] array_index_76644[10];
  wire [31:0] array_index_76645[10];
  wire [31:0] smul_76649;
  wire [31:0] add_76651;
  wire [31:0] array_update_76653[10];
  wire [31:0] add_76654;
  wire [31:0] array_update_76655[10][10];
  wire [31:0] array_index_76657[10];
  wire [31:0] array_index_76658[10];
  wire [31:0] smul_76662;
  wire [31:0] add_76664;
  wire [31:0] array_update_76666[10];
  wire [31:0] add_76667;
  wire [31:0] array_update_76668[10][10];
  wire [31:0] array_index_76670[10];
  wire [31:0] array_index_76671[10];
  wire [31:0] smul_76675;
  wire [31:0] add_76677;
  wire [31:0] array_update_76679[10];
  wire [31:0] add_76680;
  wire [31:0] array_update_76681[10][10];
  wire [31:0] array_index_76683[10];
  wire [31:0] array_index_76684[10];
  wire [31:0] smul_76688;
  wire [31:0] add_76690;
  wire [31:0] array_update_76692[10];
  wire [31:0] add_76693;
  wire [31:0] array_update_76694[10][10];
  wire [31:0] array_index_76696[10];
  wire [31:0] array_index_76697[10];
  wire [31:0] smul_76701;
  wire [31:0] add_76703;
  wire [31:0] array_update_76705[10];
  wire [31:0] add_76706;
  wire [31:0] array_update_76707[10][10];
  wire [31:0] array_index_76709[10];
  wire [31:0] array_index_76710[10];
  wire [31:0] smul_76714;
  wire [31:0] add_76716;
  wire [31:0] array_update_76718[10];
  wire [31:0] add_76719;
  wire [31:0] array_update_76720[10][10];
  wire [31:0] array_index_76722[10];
  wire [31:0] array_index_76723[10];
  wire [31:0] smul_76727;
  wire [31:0] add_76729;
  wire [31:0] array_update_76731[10];
  wire [31:0] add_76732;
  wire [31:0] array_update_76733[10][10];
  wire [31:0] array_index_76735[10];
  wire [31:0] array_index_76736[10];
  wire [31:0] smul_76740;
  wire [31:0] add_76742;
  wire [31:0] array_update_76743[10];
  wire [31:0] array_update_76744[10][10];
  wire [31:0] array_index_76746[10];
  wire [31:0] add_76748;
  wire [31:0] array_update_76749[10];
  wire [31:0] literal_76750;
  wire [31:0] array_update_76751[10][10];
  wire [31:0] array_index_76753[10];
  wire [31:0] array_index_76754[10];
  wire [31:0] smul_76758;
  wire [31:0] add_76760;
  wire [31:0] array_update_76762[10];
  wire [31:0] add_76763;
  wire [31:0] array_update_76764[10][10];
  wire [31:0] array_index_76766[10];
  wire [31:0] array_index_76767[10];
  wire [31:0] smul_76771;
  wire [31:0] add_76773;
  wire [31:0] array_update_76775[10];
  wire [31:0] add_76776;
  wire [31:0] array_update_76777[10][10];
  wire [31:0] array_index_76779[10];
  wire [31:0] array_index_76780[10];
  wire [31:0] smul_76784;
  wire [31:0] add_76786;
  wire [31:0] array_update_76788[10];
  wire [31:0] add_76789;
  wire [31:0] array_update_76790[10][10];
  wire [31:0] array_index_76792[10];
  wire [31:0] array_index_76793[10];
  wire [31:0] smul_76797;
  wire [31:0] add_76799;
  wire [31:0] array_update_76801[10];
  wire [31:0] add_76802;
  wire [31:0] array_update_76803[10][10];
  wire [31:0] array_index_76805[10];
  wire [31:0] array_index_76806[10];
  wire [31:0] smul_76810;
  wire [31:0] add_76812;
  wire [31:0] array_update_76814[10];
  wire [31:0] add_76815;
  wire [31:0] array_update_76816[10][10];
  wire [31:0] array_index_76818[10];
  wire [31:0] array_index_76819[10];
  wire [31:0] smul_76823;
  wire [31:0] add_76825;
  wire [31:0] array_update_76827[10];
  wire [31:0] add_76828;
  wire [31:0] array_update_76829[10][10];
  wire [31:0] array_index_76831[10];
  wire [31:0] array_index_76832[10];
  wire [31:0] smul_76836;
  wire [31:0] add_76838;
  wire [31:0] array_update_76840[10];
  wire [31:0] add_76841;
  wire [31:0] array_update_76842[10][10];
  wire [31:0] array_index_76844[10];
  wire [31:0] array_index_76845[10];
  wire [31:0] smul_76849;
  wire [31:0] add_76851;
  wire [31:0] array_update_76853[10];
  wire [31:0] add_76854;
  wire [31:0] array_update_76855[10][10];
  wire [31:0] array_index_76857[10];
  wire [31:0] array_index_76858[10];
  wire [31:0] smul_76862;
  wire [31:0] add_76864;
  wire [31:0] array_update_76866[10];
  wire [31:0] add_76867;
  wire [31:0] array_update_76868[10][10];
  wire [31:0] array_index_76870[10];
  wire [31:0] array_index_76871[10];
  wire [31:0] smul_76875;
  wire [31:0] add_76877;
  wire [31:0] array_update_76878[10];
  wire [31:0] array_update_76879[10][10];
  wire [31:0] array_index_76881[10];
  wire [31:0] add_76883;
  wire [31:0] array_update_76884[10];
  wire [31:0] literal_76885;
  wire [31:0] array_update_76886[10][10];
  wire [31:0] array_index_76888[10];
  wire [31:0] array_index_76889[10];
  wire [31:0] smul_76893;
  wire [31:0] add_76895;
  wire [31:0] array_update_76897[10];
  wire [31:0] add_76898;
  wire [31:0] array_update_76899[10][10];
  wire [31:0] array_index_76901[10];
  wire [31:0] array_index_76902[10];
  wire [31:0] smul_76906;
  wire [31:0] add_76908;
  wire [31:0] array_update_76910[10];
  wire [31:0] add_76911;
  wire [31:0] array_update_76912[10][10];
  wire [31:0] array_index_76914[10];
  wire [31:0] array_index_76915[10];
  wire [31:0] smul_76919;
  wire [31:0] add_76921;
  wire [31:0] array_update_76923[10];
  wire [31:0] add_76924;
  wire [31:0] array_update_76925[10][10];
  wire [31:0] array_index_76927[10];
  wire [31:0] array_index_76928[10];
  wire [31:0] smul_76932;
  wire [31:0] add_76934;
  wire [31:0] array_update_76936[10];
  wire [31:0] add_76937;
  wire [31:0] array_update_76938[10][10];
  wire [31:0] array_index_76940[10];
  wire [31:0] array_index_76941[10];
  wire [31:0] smul_76945;
  wire [31:0] add_76947;
  wire [31:0] array_update_76949[10];
  wire [31:0] add_76950;
  wire [31:0] array_update_76951[10][10];
  wire [31:0] array_index_76953[10];
  wire [31:0] array_index_76954[10];
  wire [31:0] smul_76958;
  wire [31:0] add_76960;
  wire [31:0] array_update_76962[10];
  wire [31:0] add_76963;
  wire [31:0] array_update_76964[10][10];
  wire [31:0] array_index_76966[10];
  wire [31:0] array_index_76967[10];
  wire [31:0] smul_76971;
  wire [31:0] add_76973;
  wire [31:0] array_update_76975[10];
  wire [31:0] add_76976;
  wire [31:0] array_update_76977[10][10];
  wire [31:0] array_index_76979[10];
  wire [31:0] array_index_76980[10];
  wire [31:0] smul_76984;
  wire [31:0] add_76986;
  wire [31:0] array_update_76988[10];
  wire [31:0] add_76989;
  wire [31:0] array_update_76990[10][10];
  wire [31:0] array_index_76992[10];
  wire [31:0] array_index_76993[10];
  wire [31:0] smul_76997;
  wire [31:0] add_76999;
  wire [31:0] array_update_77001[10];
  wire [31:0] add_77002;
  wire [31:0] array_update_77003[10][10];
  wire [31:0] array_index_77005[10];
  wire [31:0] array_index_77006[10];
  wire [31:0] smul_77010;
  wire [31:0] add_77012;
  wire [31:0] array_update_77013[10];
  wire [31:0] array_update_77014[10][10];
  wire [31:0] array_index_77016[10];
  wire [31:0] add_77018;
  wire [31:0] array_update_77019[10];
  wire [31:0] literal_77020;
  wire [31:0] array_update_77021[10][10];
  wire [31:0] array_index_77023[10];
  wire [31:0] array_index_77024[10];
  wire [31:0] smul_77028;
  wire [31:0] add_77030;
  wire [31:0] array_update_77032[10];
  wire [31:0] add_77033;
  wire [31:0] array_update_77034[10][10];
  wire [31:0] array_index_77036[10];
  wire [31:0] array_index_77037[10];
  wire [31:0] smul_77041;
  wire [31:0] add_77043;
  wire [31:0] array_update_77045[10];
  wire [31:0] add_77046;
  wire [31:0] array_update_77047[10][10];
  wire [31:0] array_index_77049[10];
  wire [31:0] array_index_77050[10];
  wire [31:0] smul_77054;
  wire [31:0] add_77056;
  wire [31:0] array_update_77058[10];
  wire [31:0] add_77059;
  wire [31:0] array_update_77060[10][10];
  wire [31:0] array_index_77062[10];
  wire [31:0] array_index_77063[10];
  wire [31:0] smul_77067;
  wire [31:0] add_77069;
  wire [31:0] array_update_77071[10];
  wire [31:0] add_77072;
  wire [31:0] array_update_77073[10][10];
  wire [31:0] array_index_77075[10];
  wire [31:0] array_index_77076[10];
  wire [31:0] smul_77080;
  wire [31:0] add_77082;
  wire [31:0] array_update_77084[10];
  wire [31:0] add_77085;
  wire [31:0] array_update_77086[10][10];
  wire [31:0] array_index_77088[10];
  wire [31:0] array_index_77089[10];
  wire [31:0] smul_77093;
  wire [31:0] add_77095;
  wire [31:0] array_update_77097[10];
  wire [31:0] add_77098;
  wire [31:0] array_update_77099[10][10];
  wire [31:0] array_index_77101[10];
  wire [31:0] array_index_77102[10];
  wire [31:0] smul_77106;
  wire [31:0] add_77108;
  wire [31:0] array_update_77110[10];
  wire [31:0] add_77111;
  wire [31:0] array_update_77112[10][10];
  wire [31:0] array_index_77114[10];
  wire [31:0] array_index_77115[10];
  wire [31:0] smul_77119;
  wire [31:0] add_77121;
  wire [31:0] array_update_77123[10];
  wire [31:0] add_77124;
  wire [31:0] array_update_77125[10][10];
  wire [31:0] array_index_77127[10];
  wire [31:0] array_index_77128[10];
  wire [31:0] smul_77132;
  wire [31:0] add_77134;
  wire [31:0] array_update_77136[10];
  wire [31:0] add_77137;
  wire [31:0] array_update_77138[10][10];
  wire [31:0] array_index_77140[10];
  wire [31:0] array_index_77141[10];
  wire [31:0] smul_77145;
  wire [31:0] add_77147;
  wire [31:0] array_update_77148[10];
  wire [31:0] array_update_77149[10][10];
  wire [31:0] array_index_77151[10];
  wire [31:0] add_77153;
  wire [31:0] array_update_77154[10];
  wire [31:0] literal_77155;
  wire [31:0] array_update_77156[10][10];
  wire [31:0] array_index_77158[10];
  wire [31:0] array_index_77159[10];
  wire [31:0] smul_77163;
  wire [31:0] add_77165;
  wire [31:0] array_update_77167[10];
  wire [31:0] add_77168;
  wire [31:0] array_update_77169[10][10];
  wire [31:0] array_index_77171[10];
  wire [31:0] array_index_77172[10];
  wire [31:0] smul_77176;
  wire [31:0] add_77178;
  wire [31:0] array_update_77180[10];
  wire [31:0] add_77181;
  wire [31:0] array_update_77182[10][10];
  wire [31:0] array_index_77184[10];
  wire [31:0] array_index_77185[10];
  wire [31:0] smul_77189;
  wire [31:0] add_77191;
  wire [31:0] array_update_77193[10];
  wire [31:0] add_77194;
  wire [31:0] array_update_77195[10][10];
  wire [31:0] array_index_77197[10];
  wire [31:0] array_index_77198[10];
  wire [31:0] smul_77202;
  wire [31:0] add_77204;
  wire [31:0] array_update_77206[10];
  wire [31:0] add_77207;
  wire [31:0] array_update_77208[10][10];
  wire [31:0] array_index_77210[10];
  wire [31:0] array_index_77211[10];
  wire [31:0] smul_77215;
  wire [31:0] add_77217;
  wire [31:0] array_update_77219[10];
  wire [31:0] add_77220;
  wire [31:0] array_update_77221[10][10];
  wire [31:0] array_index_77223[10];
  wire [31:0] array_index_77224[10];
  wire [31:0] smul_77228;
  wire [31:0] add_77230;
  wire [31:0] array_update_77232[10];
  wire [31:0] add_77233;
  wire [31:0] array_update_77234[10][10];
  wire [31:0] array_index_77236[10];
  wire [31:0] array_index_77237[10];
  wire [31:0] smul_77241;
  wire [31:0] add_77243;
  wire [31:0] array_update_77245[10];
  wire [31:0] add_77246;
  wire [31:0] array_update_77247[10][10];
  wire [31:0] array_index_77249[10];
  wire [31:0] array_index_77250[10];
  wire [31:0] smul_77254;
  wire [31:0] add_77256;
  wire [31:0] array_update_77258[10];
  wire [31:0] add_77259;
  wire [31:0] array_update_77260[10][10];
  wire [31:0] array_index_77262[10];
  wire [31:0] array_index_77263[10];
  wire [31:0] smul_77267;
  wire [31:0] add_77269;
  wire [31:0] array_update_77271[10];
  wire [31:0] add_77272;
  wire [31:0] array_update_77273[10][10];
  wire [31:0] array_index_77275[10];
  wire [31:0] array_index_77276[10];
  wire [31:0] smul_77280;
  wire [31:0] add_77282;
  wire [31:0] array_update_77283[10];
  wire [31:0] array_update_77284[10][10];
  wire [31:0] array_index_77286[10];
  wire [31:0] add_77288;
  wire [31:0] array_update_77289[10];
  wire [31:0] literal_77290;
  wire [31:0] array_update_77291[10][10];
  wire [31:0] array_index_77293[10];
  wire [31:0] array_index_77294[10];
  wire [31:0] smul_77298;
  wire [31:0] add_77300;
  wire [31:0] array_update_77302[10];
  wire [31:0] add_77303;
  wire [31:0] array_update_77304[10][10];
  wire [31:0] array_index_77306[10];
  wire [31:0] array_index_77307[10];
  wire [31:0] smul_77311;
  wire [31:0] add_77313;
  wire [31:0] array_update_77315[10];
  wire [31:0] add_77316;
  wire [31:0] array_update_77317[10][10];
  wire [31:0] array_index_77319[10];
  wire [31:0] array_index_77320[10];
  wire [31:0] smul_77324;
  wire [31:0] add_77326;
  wire [31:0] array_update_77328[10];
  wire [31:0] add_77329;
  wire [31:0] array_update_77330[10][10];
  wire [31:0] array_index_77332[10];
  wire [31:0] array_index_77333[10];
  wire [31:0] smul_77337;
  wire [31:0] add_77339;
  wire [31:0] array_update_77341[10];
  wire [31:0] add_77342;
  wire [31:0] array_update_77343[10][10];
  wire [31:0] array_index_77345[10];
  wire [31:0] array_index_77346[10];
  wire [31:0] smul_77350;
  wire [31:0] add_77352;
  wire [31:0] array_update_77354[10];
  wire [31:0] add_77355;
  wire [31:0] array_update_77356[10][10];
  wire [31:0] array_index_77358[10];
  wire [31:0] array_index_77359[10];
  wire [31:0] smul_77363;
  wire [31:0] add_77365;
  wire [31:0] array_update_77367[10];
  wire [31:0] add_77368;
  wire [31:0] array_update_77369[10][10];
  wire [31:0] array_index_77371[10];
  wire [31:0] array_index_77372[10];
  wire [31:0] smul_77376;
  wire [31:0] add_77378;
  wire [31:0] array_update_77380[10];
  wire [31:0] add_77381;
  wire [31:0] array_update_77382[10][10];
  wire [31:0] array_index_77384[10];
  wire [31:0] array_index_77385[10];
  wire [31:0] smul_77389;
  wire [31:0] add_77391;
  wire [31:0] array_update_77393[10];
  wire [31:0] add_77394;
  wire [31:0] array_update_77395[10][10];
  wire [31:0] array_index_77397[10];
  wire [31:0] array_index_77398[10];
  wire [31:0] smul_77402;
  wire [31:0] add_77404;
  wire [31:0] array_update_77406[10];
  wire [31:0] add_77407;
  wire [31:0] array_update_77408[10][10];
  wire [31:0] array_index_77410[10];
  wire [31:0] array_index_77411[10];
  wire [31:0] smul_77415;
  wire [31:0] add_77417;
  wire [31:0] array_update_77418[10];
  wire [31:0] array_update_77420[10][10];
  wire [31:0] add_77421;
  wire [31:0] array_index_77422[10];
  wire [31:0] literal_77424;
  wire [31:0] array_update_77425[10];
  wire [31:0] literal_77426;
  wire [31:0] array_update_77427[10][10];
  wire [31:0] array_index_77428[10];
  wire [31:0] array_index_77429[10];
  wire [31:0] array_index_77430[10];
  wire [31:0] smul_77434;
  wire [31:0] add_77436;
  wire [31:0] array_update_77438[10];
  wire [31:0] add_77439;
  wire [31:0] array_update_77440[10][10];
  wire [31:0] array_index_77442[10];
  wire [31:0] array_index_77443[10];
  wire [31:0] smul_77447;
  wire [31:0] add_77449;
  wire [31:0] array_update_77451[10];
  wire [31:0] add_77452;
  wire [31:0] array_update_77453[10][10];
  wire [31:0] array_index_77455[10];
  wire [31:0] array_index_77456[10];
  wire [31:0] smul_77460;
  wire [31:0] add_77462;
  wire [31:0] array_update_77464[10];
  wire [31:0] add_77465;
  wire [31:0] array_update_77466[10][10];
  wire [31:0] array_index_77468[10];
  wire [31:0] array_index_77469[10];
  wire [31:0] smul_77473;
  wire [31:0] add_77475;
  wire [31:0] array_update_77477[10];
  wire [31:0] add_77478;
  wire [31:0] array_update_77479[10][10];
  wire [31:0] array_index_77481[10];
  wire [31:0] array_index_77482[10];
  wire [31:0] smul_77486;
  wire [31:0] add_77488;
  wire [31:0] array_update_77490[10];
  wire [31:0] add_77491;
  wire [31:0] array_update_77492[10][10];
  wire [31:0] array_index_77494[10];
  wire [31:0] array_index_77495[10];
  wire [31:0] smul_77499;
  wire [31:0] add_77501;
  wire [31:0] array_update_77503[10];
  wire [31:0] add_77504;
  wire [31:0] array_update_77505[10][10];
  wire [31:0] array_index_77507[10];
  wire [31:0] array_index_77508[10];
  wire [31:0] smul_77512;
  wire [31:0] add_77514;
  wire [31:0] array_update_77516[10];
  wire [31:0] add_77517;
  wire [31:0] array_update_77518[10][10];
  wire [31:0] array_index_77520[10];
  wire [31:0] array_index_77521[10];
  wire [31:0] smul_77525;
  wire [31:0] add_77527;
  wire [31:0] array_update_77529[10];
  wire [31:0] add_77530;
  wire [31:0] array_update_77531[10][10];
  wire [31:0] array_index_77533[10];
  wire [31:0] array_index_77534[10];
  wire [31:0] smul_77538;
  wire [31:0] add_77540;
  wire [31:0] array_update_77542[10];
  wire [31:0] add_77543;
  wire [31:0] array_update_77544[10][10];
  wire [31:0] array_index_77546[10];
  wire [31:0] array_index_77547[10];
  wire [31:0] smul_77551;
  wire [31:0] add_77553;
  wire [31:0] array_update_77554[10];
  wire [31:0] array_update_77555[10][10];
  wire [31:0] array_index_77557[10];
  wire [31:0] add_77559;
  wire [31:0] array_update_77560[10];
  wire [31:0] literal_77561;
  wire [31:0] array_update_77562[10][10];
  wire [31:0] array_index_77564[10];
  wire [31:0] array_index_77565[10];
  wire [31:0] smul_77569;
  wire [31:0] add_77571;
  wire [31:0] array_update_77573[10];
  wire [31:0] add_77574;
  wire [31:0] array_update_77575[10][10];
  wire [31:0] array_index_77577[10];
  wire [31:0] array_index_77578[10];
  wire [31:0] smul_77582;
  wire [31:0] add_77584;
  wire [31:0] array_update_77586[10];
  wire [31:0] add_77587;
  wire [31:0] array_update_77588[10][10];
  wire [31:0] array_index_77590[10];
  wire [31:0] array_index_77591[10];
  wire [31:0] smul_77595;
  wire [31:0] add_77597;
  wire [31:0] array_update_77599[10];
  wire [31:0] add_77600;
  wire [31:0] array_update_77601[10][10];
  wire [31:0] array_index_77603[10];
  wire [31:0] array_index_77604[10];
  wire [31:0] smul_77608;
  wire [31:0] add_77610;
  wire [31:0] array_update_77612[10];
  wire [31:0] add_77613;
  wire [31:0] array_update_77614[10][10];
  wire [31:0] array_index_77616[10];
  wire [31:0] array_index_77617[10];
  wire [31:0] smul_77621;
  wire [31:0] add_77623;
  wire [31:0] array_update_77625[10];
  wire [31:0] add_77626;
  wire [31:0] array_update_77627[10][10];
  wire [31:0] array_index_77629[10];
  wire [31:0] array_index_77630[10];
  wire [31:0] smul_77634;
  wire [31:0] add_77636;
  wire [31:0] array_update_77638[10];
  wire [31:0] add_77639;
  wire [31:0] array_update_77640[10][10];
  wire [31:0] array_index_77642[10];
  wire [31:0] array_index_77643[10];
  wire [31:0] smul_77647;
  wire [31:0] add_77649;
  wire [31:0] array_update_77651[10];
  wire [31:0] add_77652;
  wire [31:0] array_update_77653[10][10];
  wire [31:0] array_index_77655[10];
  wire [31:0] array_index_77656[10];
  wire [31:0] smul_77660;
  wire [31:0] add_77662;
  wire [31:0] array_update_77664[10];
  wire [31:0] add_77665;
  wire [31:0] array_update_77666[10][10];
  wire [31:0] array_index_77668[10];
  wire [31:0] array_index_77669[10];
  wire [31:0] smul_77673;
  wire [31:0] add_77675;
  wire [31:0] array_update_77677[10];
  wire [31:0] add_77678;
  wire [31:0] array_update_77679[10][10];
  wire [31:0] array_index_77681[10];
  wire [31:0] array_index_77682[10];
  wire [31:0] smul_77686;
  wire [31:0] add_77688;
  wire [31:0] array_update_77689[10];
  wire [31:0] array_update_77690[10][10];
  wire [31:0] array_index_77692[10];
  wire [31:0] add_77694;
  wire [31:0] array_update_77695[10];
  wire [31:0] literal_77696;
  wire [31:0] array_update_77697[10][10];
  wire [31:0] array_index_77699[10];
  wire [31:0] array_index_77700[10];
  wire [31:0] smul_77704;
  wire [31:0] add_77706;
  wire [31:0] array_update_77708[10];
  wire [31:0] add_77709;
  wire [31:0] array_update_77710[10][10];
  wire [31:0] array_index_77712[10];
  wire [31:0] array_index_77713[10];
  wire [31:0] smul_77717;
  wire [31:0] add_77719;
  wire [31:0] array_update_77721[10];
  wire [31:0] add_77722;
  wire [31:0] array_update_77723[10][10];
  wire [31:0] array_index_77725[10];
  wire [31:0] array_index_77726[10];
  wire [31:0] smul_77730;
  wire [31:0] add_77732;
  wire [31:0] array_update_77734[10];
  wire [31:0] add_77735;
  wire [31:0] array_update_77736[10][10];
  wire [31:0] array_index_77738[10];
  wire [31:0] array_index_77739[10];
  wire [31:0] smul_77743;
  wire [31:0] add_77745;
  wire [31:0] array_update_77747[10];
  wire [31:0] add_77748;
  wire [31:0] array_update_77749[10][10];
  wire [31:0] array_index_77751[10];
  wire [31:0] array_index_77752[10];
  wire [31:0] smul_77756;
  wire [31:0] add_77758;
  wire [31:0] array_update_77760[10];
  wire [31:0] add_77761;
  wire [31:0] array_update_77762[10][10];
  wire [31:0] array_index_77764[10];
  wire [31:0] array_index_77765[10];
  wire [31:0] smul_77769;
  wire [31:0] add_77771;
  wire [31:0] array_update_77773[10];
  wire [31:0] add_77774;
  wire [31:0] array_update_77775[10][10];
  wire [31:0] array_index_77777[10];
  wire [31:0] array_index_77778[10];
  wire [31:0] smul_77782;
  wire [31:0] add_77784;
  wire [31:0] array_update_77786[10];
  wire [31:0] add_77787;
  wire [31:0] array_update_77788[10][10];
  wire [31:0] array_index_77790[10];
  wire [31:0] array_index_77791[10];
  wire [31:0] smul_77795;
  wire [31:0] add_77797;
  wire [31:0] array_update_77799[10];
  wire [31:0] add_77800;
  wire [31:0] array_update_77801[10][10];
  wire [31:0] array_index_77803[10];
  wire [31:0] array_index_77804[10];
  wire [31:0] smul_77808;
  wire [31:0] add_77810;
  wire [31:0] array_update_77812[10];
  wire [31:0] add_77813;
  wire [31:0] array_update_77814[10][10];
  wire [31:0] array_index_77816[10];
  wire [31:0] array_index_77817[10];
  wire [31:0] smul_77821;
  wire [31:0] add_77823;
  wire [31:0] array_update_77824[10];
  wire [31:0] array_update_77825[10][10];
  wire [31:0] array_index_77827[10];
  wire [31:0] add_77829;
  wire [31:0] array_update_77830[10];
  wire [31:0] literal_77831;
  wire [31:0] array_update_77832[10][10];
  wire [31:0] array_index_77834[10];
  wire [31:0] array_index_77835[10];
  wire [31:0] smul_77839;
  wire [31:0] add_77841;
  wire [31:0] array_update_77843[10];
  wire [31:0] add_77844;
  wire [31:0] array_update_77845[10][10];
  wire [31:0] array_index_77847[10];
  wire [31:0] array_index_77848[10];
  wire [31:0] smul_77852;
  wire [31:0] add_77854;
  wire [31:0] array_update_77856[10];
  wire [31:0] add_77857;
  wire [31:0] array_update_77858[10][10];
  wire [31:0] array_index_77860[10];
  wire [31:0] array_index_77861[10];
  wire [31:0] smul_77865;
  wire [31:0] add_77867;
  wire [31:0] array_update_77869[10];
  wire [31:0] add_77870;
  wire [31:0] array_update_77871[10][10];
  wire [31:0] array_index_77873[10];
  wire [31:0] array_index_77874[10];
  wire [31:0] smul_77878;
  wire [31:0] add_77880;
  wire [31:0] array_update_77882[10];
  wire [31:0] add_77883;
  wire [31:0] array_update_77884[10][10];
  wire [31:0] array_index_77886[10];
  wire [31:0] array_index_77887[10];
  wire [31:0] smul_77891;
  wire [31:0] add_77893;
  wire [31:0] array_update_77895[10];
  wire [31:0] add_77896;
  wire [31:0] array_update_77897[10][10];
  wire [31:0] array_index_77899[10];
  wire [31:0] array_index_77900[10];
  wire [31:0] smul_77904;
  wire [31:0] add_77906;
  wire [31:0] array_update_77908[10];
  wire [31:0] add_77909;
  wire [31:0] array_update_77910[10][10];
  wire [31:0] array_index_77912[10];
  wire [31:0] array_index_77913[10];
  wire [31:0] smul_77917;
  wire [31:0] add_77919;
  wire [31:0] array_update_77921[10];
  wire [31:0] add_77922;
  wire [31:0] array_update_77923[10][10];
  wire [31:0] array_index_77925[10];
  wire [31:0] array_index_77926[10];
  wire [31:0] smul_77930;
  wire [31:0] add_77932;
  wire [31:0] array_update_77934[10];
  wire [31:0] add_77935;
  wire [31:0] array_update_77936[10][10];
  wire [31:0] array_index_77938[10];
  wire [31:0] array_index_77939[10];
  wire [31:0] smul_77943;
  wire [31:0] add_77945;
  wire [31:0] array_update_77947[10];
  wire [31:0] add_77948;
  wire [31:0] array_update_77949[10][10];
  wire [31:0] array_index_77951[10];
  wire [31:0] array_index_77952[10];
  wire [31:0] smul_77956;
  wire [31:0] add_77958;
  wire [31:0] array_update_77959[10];
  wire [31:0] array_update_77960[10][10];
  wire [31:0] array_index_77962[10];
  wire [31:0] add_77964;
  wire [31:0] array_update_77965[10];
  wire [31:0] literal_77966;
  wire [31:0] array_update_77967[10][10];
  wire [31:0] array_index_77969[10];
  wire [31:0] array_index_77970[10];
  wire [31:0] smul_77974;
  wire [31:0] add_77976;
  wire [31:0] array_update_77978[10];
  wire [31:0] add_77979;
  wire [31:0] array_update_77980[10][10];
  wire [31:0] array_index_77982[10];
  wire [31:0] array_index_77983[10];
  wire [31:0] smul_77987;
  wire [31:0] add_77989;
  wire [31:0] array_update_77991[10];
  wire [31:0] add_77992;
  wire [31:0] array_update_77993[10][10];
  wire [31:0] array_index_77995[10];
  wire [31:0] array_index_77996[10];
  wire [31:0] smul_78000;
  wire [31:0] add_78002;
  wire [31:0] array_update_78004[10];
  wire [31:0] add_78005;
  wire [31:0] array_update_78006[10][10];
  wire [31:0] array_index_78008[10];
  wire [31:0] array_index_78009[10];
  wire [31:0] smul_78013;
  wire [31:0] add_78015;
  wire [31:0] array_update_78017[10];
  wire [31:0] add_78018;
  wire [31:0] array_update_78019[10][10];
  wire [31:0] array_index_78021[10];
  wire [31:0] array_index_78022[10];
  wire [31:0] smul_78026;
  wire [31:0] add_78028;
  wire [31:0] array_update_78030[10];
  wire [31:0] add_78031;
  wire [31:0] array_update_78032[10][10];
  wire [31:0] array_index_78034[10];
  wire [31:0] array_index_78035[10];
  wire [31:0] smul_78039;
  wire [31:0] add_78041;
  wire [31:0] array_update_78043[10];
  wire [31:0] add_78044;
  wire [31:0] array_update_78045[10][10];
  wire [31:0] array_index_78047[10];
  wire [31:0] array_index_78048[10];
  wire [31:0] smul_78052;
  wire [31:0] add_78054;
  wire [31:0] array_update_78056[10];
  wire [31:0] add_78057;
  wire [31:0] array_update_78058[10][10];
  wire [31:0] array_index_78060[10];
  wire [31:0] array_index_78061[10];
  wire [31:0] smul_78065;
  wire [31:0] add_78067;
  wire [31:0] array_update_78069[10];
  wire [31:0] add_78070;
  wire [31:0] array_update_78071[10][10];
  wire [31:0] array_index_78073[10];
  wire [31:0] array_index_78074[10];
  wire [31:0] smul_78078;
  wire [31:0] add_78080;
  wire [31:0] array_update_78082[10];
  wire [31:0] add_78083;
  wire [31:0] array_update_78084[10][10];
  wire [31:0] array_index_78086[10];
  wire [31:0] array_index_78087[10];
  wire [31:0] smul_78091;
  wire [31:0] add_78093;
  wire [31:0] array_update_78094[10];
  wire [31:0] array_update_78095[10][10];
  wire [31:0] array_index_78097[10];
  wire [31:0] add_78099;
  wire [31:0] array_update_78100[10];
  wire [31:0] literal_78101;
  wire [31:0] array_update_78102[10][10];
  wire [31:0] array_index_78104[10];
  wire [31:0] array_index_78105[10];
  wire [31:0] smul_78109;
  wire [31:0] add_78111;
  wire [31:0] array_update_78113[10];
  wire [31:0] add_78114;
  wire [31:0] array_update_78115[10][10];
  wire [31:0] array_index_78117[10];
  wire [31:0] array_index_78118[10];
  wire [31:0] smul_78122;
  wire [31:0] add_78124;
  wire [31:0] array_update_78126[10];
  wire [31:0] add_78127;
  wire [31:0] array_update_78128[10][10];
  wire [31:0] array_index_78130[10];
  wire [31:0] array_index_78131[10];
  wire [31:0] smul_78135;
  wire [31:0] add_78137;
  wire [31:0] array_update_78139[10];
  wire [31:0] add_78140;
  wire [31:0] array_update_78141[10][10];
  wire [31:0] array_index_78143[10];
  wire [31:0] array_index_78144[10];
  wire [31:0] smul_78148;
  wire [31:0] add_78150;
  wire [31:0] array_update_78152[10];
  wire [31:0] add_78153;
  wire [31:0] array_update_78154[10][10];
  wire [31:0] array_index_78156[10];
  wire [31:0] array_index_78157[10];
  wire [31:0] smul_78161;
  wire [31:0] add_78163;
  wire [31:0] array_update_78165[10];
  wire [31:0] add_78166;
  wire [31:0] array_update_78167[10][10];
  wire [31:0] array_index_78169[10];
  wire [31:0] array_index_78170[10];
  wire [31:0] smul_78174;
  wire [31:0] add_78176;
  wire [31:0] array_update_78178[10];
  wire [31:0] add_78179;
  wire [31:0] array_update_78180[10][10];
  wire [31:0] array_index_78182[10];
  wire [31:0] array_index_78183[10];
  wire [31:0] smul_78187;
  wire [31:0] add_78189;
  wire [31:0] array_update_78191[10];
  wire [31:0] add_78192;
  wire [31:0] array_update_78193[10][10];
  wire [31:0] array_index_78195[10];
  wire [31:0] array_index_78196[10];
  wire [31:0] smul_78200;
  wire [31:0] add_78202;
  wire [31:0] array_update_78204[10];
  wire [31:0] add_78205;
  wire [31:0] array_update_78206[10][10];
  wire [31:0] array_index_78208[10];
  wire [31:0] array_index_78209[10];
  wire [31:0] smul_78213;
  wire [31:0] add_78215;
  wire [31:0] array_update_78217[10];
  wire [31:0] add_78218;
  wire [31:0] array_update_78219[10][10];
  wire [31:0] array_index_78221[10];
  wire [31:0] array_index_78222[10];
  wire [31:0] smul_78226;
  wire [31:0] add_78228;
  wire [31:0] array_update_78229[10];
  wire [31:0] array_update_78230[10][10];
  wire [31:0] array_index_78232[10];
  wire [31:0] add_78234;
  wire [31:0] array_update_78235[10];
  wire [31:0] literal_78236;
  wire [31:0] array_update_78237[10][10];
  wire [31:0] array_index_78239[10];
  wire [31:0] array_index_78240[10];
  wire [31:0] smul_78244;
  wire [31:0] add_78246;
  wire [31:0] array_update_78248[10];
  wire [31:0] add_78249;
  wire [31:0] array_update_78250[10][10];
  wire [31:0] array_index_78252[10];
  wire [31:0] array_index_78253[10];
  wire [31:0] smul_78257;
  wire [31:0] add_78259;
  wire [31:0] array_update_78261[10];
  wire [31:0] add_78262;
  wire [31:0] array_update_78263[10][10];
  wire [31:0] array_index_78265[10];
  wire [31:0] array_index_78266[10];
  wire [31:0] smul_78270;
  wire [31:0] add_78272;
  wire [31:0] array_update_78274[10];
  wire [31:0] add_78275;
  wire [31:0] array_update_78276[10][10];
  wire [31:0] array_index_78278[10];
  wire [31:0] array_index_78279[10];
  wire [31:0] smul_78283;
  wire [31:0] add_78285;
  wire [31:0] array_update_78287[10];
  wire [31:0] add_78288;
  wire [31:0] array_update_78289[10][10];
  wire [31:0] array_index_78291[10];
  wire [31:0] array_index_78292[10];
  wire [31:0] smul_78296;
  wire [31:0] add_78298;
  wire [31:0] array_update_78300[10];
  wire [31:0] add_78301;
  wire [31:0] array_update_78302[10][10];
  wire [31:0] array_index_78304[10];
  wire [31:0] array_index_78305[10];
  wire [31:0] smul_78309;
  wire [31:0] add_78311;
  wire [31:0] array_update_78313[10];
  wire [31:0] add_78314;
  wire [31:0] array_update_78315[10][10];
  wire [31:0] array_index_78317[10];
  wire [31:0] array_index_78318[10];
  wire [31:0] smul_78322;
  wire [31:0] add_78324;
  wire [31:0] array_update_78326[10];
  wire [31:0] add_78327;
  wire [31:0] array_update_78328[10][10];
  wire [31:0] array_index_78330[10];
  wire [31:0] array_index_78331[10];
  wire [31:0] smul_78335;
  wire [31:0] add_78337;
  wire [31:0] array_update_78339[10];
  wire [31:0] add_78340;
  wire [31:0] array_update_78341[10][10];
  wire [31:0] array_index_78343[10];
  wire [31:0] array_index_78344[10];
  wire [31:0] smul_78348;
  wire [31:0] add_78350;
  wire [31:0] array_update_78352[10];
  wire [31:0] add_78353;
  wire [31:0] array_update_78354[10][10];
  wire [31:0] array_index_78356[10];
  wire [31:0] array_index_78357[10];
  wire [31:0] smul_78361;
  wire [31:0] add_78363;
  wire [31:0] array_update_78364[10];
  wire [31:0] array_update_78365[10][10];
  wire [31:0] array_index_78367[10];
  wire [31:0] add_78369;
  wire [31:0] array_update_78370[10];
  wire [31:0] literal_78371;
  wire [31:0] array_update_78372[10][10];
  wire [31:0] array_index_78374[10];
  wire [31:0] array_index_78375[10];
  wire [31:0] smul_78379;
  wire [31:0] add_78381;
  wire [31:0] array_update_78383[10];
  wire [31:0] add_78384;
  wire [31:0] array_update_78385[10][10];
  wire [31:0] array_index_78387[10];
  wire [31:0] array_index_78388[10];
  wire [31:0] smul_78392;
  wire [31:0] add_78394;
  wire [31:0] array_update_78396[10];
  wire [31:0] add_78397;
  wire [31:0] array_update_78398[10][10];
  wire [31:0] array_index_78400[10];
  wire [31:0] array_index_78401[10];
  wire [31:0] smul_78405;
  wire [31:0] add_78407;
  wire [31:0] array_update_78409[10];
  wire [31:0] add_78410;
  wire [31:0] array_update_78411[10][10];
  wire [31:0] array_index_78413[10];
  wire [31:0] array_index_78414[10];
  wire [31:0] smul_78418;
  wire [31:0] add_78420;
  wire [31:0] array_update_78422[10];
  wire [31:0] add_78423;
  wire [31:0] array_update_78424[10][10];
  wire [31:0] array_index_78426[10];
  wire [31:0] array_index_78427[10];
  wire [31:0] smul_78431;
  wire [31:0] add_78433;
  wire [31:0] array_update_78435[10];
  wire [31:0] add_78436;
  wire [31:0] array_update_78437[10][10];
  wire [31:0] array_index_78439[10];
  wire [31:0] array_index_78440[10];
  wire [31:0] smul_78444;
  wire [31:0] add_78446;
  wire [31:0] array_update_78448[10];
  wire [31:0] add_78449;
  wire [31:0] array_update_78450[10][10];
  wire [31:0] array_index_78452[10];
  wire [31:0] array_index_78453[10];
  wire [31:0] smul_78457;
  wire [31:0] add_78459;
  wire [31:0] array_update_78461[10];
  wire [31:0] add_78462;
  wire [31:0] array_update_78463[10][10];
  wire [31:0] array_index_78465[10];
  wire [31:0] array_index_78466[10];
  wire [31:0] smul_78470;
  wire [31:0] add_78472;
  wire [31:0] array_update_78474[10];
  wire [31:0] add_78475;
  wire [31:0] array_update_78476[10][10];
  wire [31:0] array_index_78478[10];
  wire [31:0] array_index_78479[10];
  wire [31:0] smul_78483;
  wire [31:0] add_78485;
  wire [31:0] array_update_78487[10];
  wire [31:0] add_78488;
  wire [31:0] array_update_78489[10][10];
  wire [31:0] array_index_78491[10];
  wire [31:0] array_index_78492[10];
  wire [31:0] smul_78496;
  wire [31:0] add_78498;
  wire [31:0] array_update_78499[10];
  wire [31:0] array_update_78500[10][10];
  wire [31:0] array_index_78502[10];
  wire [31:0] add_78504;
  wire [31:0] array_update_78505[10];
  wire [31:0] literal_78506;
  wire [31:0] array_update_78507[10][10];
  wire [31:0] array_index_78509[10];
  wire [31:0] array_index_78510[10];
  wire [31:0] smul_78514;
  wire [31:0] add_78516;
  wire [31:0] array_update_78518[10];
  wire [31:0] add_78519;
  wire [31:0] array_update_78520[10][10];
  wire [31:0] array_index_78522[10];
  wire [31:0] array_index_78523[10];
  wire [31:0] smul_78527;
  wire [31:0] add_78529;
  wire [31:0] array_update_78531[10];
  wire [31:0] add_78532;
  wire [31:0] array_update_78533[10][10];
  wire [31:0] array_index_78535[10];
  wire [31:0] array_index_78536[10];
  wire [31:0] smul_78540;
  wire [31:0] add_78542;
  wire [31:0] array_update_78544[10];
  wire [31:0] add_78545;
  wire [31:0] array_update_78546[10][10];
  wire [31:0] array_index_78548[10];
  wire [31:0] array_index_78549[10];
  wire [31:0] smul_78553;
  wire [31:0] add_78555;
  wire [31:0] array_update_78557[10];
  wire [31:0] add_78558;
  wire [31:0] array_update_78559[10][10];
  wire [31:0] array_index_78561[10];
  wire [31:0] array_index_78562[10];
  wire [31:0] smul_78566;
  wire [31:0] add_78568;
  wire [31:0] array_update_78570[10];
  wire [31:0] add_78571;
  wire [31:0] array_update_78572[10][10];
  wire [31:0] array_index_78574[10];
  wire [31:0] array_index_78575[10];
  wire [31:0] smul_78579;
  wire [31:0] add_78581;
  wire [31:0] array_update_78583[10];
  wire [31:0] add_78584;
  wire [31:0] array_update_78585[10][10];
  wire [31:0] array_index_78587[10];
  wire [31:0] array_index_78588[10];
  wire [31:0] smul_78592;
  wire [31:0] add_78594;
  wire [31:0] array_update_78596[10];
  wire [31:0] add_78597;
  wire [31:0] array_update_78598[10][10];
  wire [31:0] array_index_78600[10];
  wire [31:0] array_index_78601[10];
  wire [31:0] smul_78605;
  wire [31:0] add_78607;
  wire [31:0] array_update_78609[10];
  wire [31:0] add_78610;
  wire [31:0] array_update_78611[10][10];
  wire [31:0] array_index_78613[10];
  wire [31:0] array_index_78614[10];
  wire [31:0] smul_78618;
  wire [31:0] add_78620;
  wire [31:0] array_update_78622[10];
  wire [31:0] add_78623;
  wire [31:0] array_update_78624[10][10];
  wire [31:0] array_index_78626[10];
  wire [31:0] array_index_78627[10];
  wire [31:0] smul_78631;
  wire [31:0] add_78633;
  wire [31:0] array_update_78634[10];
  wire [31:0] array_update_78635[10][10];
  wire [31:0] array_index_78637[10];
  wire [31:0] add_78639;
  wire [31:0] array_update_78640[10];
  wire [31:0] literal_78641;
  wire [31:0] array_update_78642[10][10];
  wire [31:0] array_index_78644[10];
  wire [31:0] array_index_78645[10];
  wire [31:0] smul_78649;
  wire [31:0] add_78651;
  wire [31:0] array_update_78653[10];
  wire [31:0] add_78654;
  wire [31:0] array_update_78655[10][10];
  wire [31:0] array_index_78657[10];
  wire [31:0] array_index_78658[10];
  wire [31:0] smul_78662;
  wire [31:0] add_78664;
  wire [31:0] array_update_78666[10];
  wire [31:0] add_78667;
  wire [31:0] array_update_78668[10][10];
  wire [31:0] array_index_78670[10];
  wire [31:0] array_index_78671[10];
  wire [31:0] smul_78675;
  wire [31:0] add_78677;
  wire [31:0] array_update_78679[10];
  wire [31:0] add_78680;
  wire [31:0] array_update_78681[10][10];
  wire [31:0] array_index_78683[10];
  wire [31:0] array_index_78684[10];
  wire [31:0] smul_78688;
  wire [31:0] add_78690;
  wire [31:0] array_update_78692[10];
  wire [31:0] add_78693;
  wire [31:0] array_update_78694[10][10];
  wire [31:0] array_index_78696[10];
  wire [31:0] array_index_78697[10];
  wire [31:0] smul_78701;
  wire [31:0] add_78703;
  wire [31:0] array_update_78705[10];
  wire [31:0] add_78706;
  wire [31:0] array_update_78707[10][10];
  wire [31:0] array_index_78709[10];
  wire [31:0] array_index_78710[10];
  wire [31:0] smul_78714;
  wire [31:0] add_78716;
  wire [31:0] array_update_78718[10];
  wire [31:0] add_78719;
  wire [31:0] array_update_78720[10][10];
  wire [31:0] array_index_78722[10];
  wire [31:0] array_index_78723[10];
  wire [31:0] smul_78727;
  wire [31:0] add_78729;
  wire [31:0] array_update_78731[10];
  wire [31:0] add_78732;
  wire [31:0] array_update_78733[10][10];
  wire [31:0] array_index_78735[10];
  wire [31:0] array_index_78736[10];
  wire [31:0] smul_78740;
  wire [31:0] add_78742;
  wire [31:0] array_update_78744[10];
  wire [31:0] add_78745;
  wire [31:0] array_update_78746[10][10];
  wire [31:0] array_index_78748[10];
  wire [31:0] array_index_78749[10];
  wire [31:0] smul_78753;
  wire [31:0] add_78755;
  wire [31:0] array_update_78757[10];
  wire [31:0] add_78758;
  wire [31:0] array_update_78759[10][10];
  wire [31:0] array_index_78761[10];
  wire [31:0] array_index_78762[10];
  wire [31:0] smul_78766;
  wire [31:0] add_78768;
  wire [31:0] array_update_78769[10];
  wire [31:0] array_update_78771[10][10];
  wire [31:0] add_78772;
  wire [31:0] array_index_78773[10];
  wire [31:0] literal_78775;
  wire [31:0] array_update_78776[10];
  wire [31:0] literal_78777;
  wire [31:0] array_update_78778[10][10];
  wire [31:0] array_index_78779[10];
  wire [31:0] array_index_78780[10];
  wire [31:0] array_index_78781[10];
  wire [31:0] smul_78785;
  wire [31:0] add_78787;
  wire [31:0] array_update_78789[10];
  wire [31:0] add_78790;
  wire [31:0] array_update_78791[10][10];
  wire [31:0] array_index_78793[10];
  wire [31:0] array_index_78794[10];
  wire [31:0] smul_78798;
  wire [31:0] add_78800;
  wire [31:0] array_update_78802[10];
  wire [31:0] add_78803;
  wire [31:0] array_update_78804[10][10];
  wire [31:0] array_index_78806[10];
  wire [31:0] array_index_78807[10];
  wire [31:0] smul_78811;
  wire [31:0] add_78813;
  wire [31:0] array_update_78815[10];
  wire [31:0] add_78816;
  wire [31:0] array_update_78817[10][10];
  wire [31:0] array_index_78819[10];
  wire [31:0] array_index_78820[10];
  wire [31:0] smul_78824;
  wire [31:0] add_78826;
  wire [31:0] array_update_78828[10];
  wire [31:0] add_78829;
  wire [31:0] array_update_78830[10][10];
  wire [31:0] array_index_78832[10];
  wire [31:0] array_index_78833[10];
  wire [31:0] smul_78837;
  wire [31:0] add_78839;
  wire [31:0] array_update_78841[10];
  wire [31:0] add_78842;
  wire [31:0] array_update_78843[10][10];
  wire [31:0] array_index_78845[10];
  wire [31:0] array_index_78846[10];
  wire [31:0] smul_78850;
  wire [31:0] add_78852;
  wire [31:0] array_update_78854[10];
  wire [31:0] add_78855;
  wire [31:0] array_update_78856[10][10];
  wire [31:0] array_index_78858[10];
  wire [31:0] array_index_78859[10];
  wire [31:0] smul_78863;
  wire [31:0] add_78865;
  wire [31:0] array_update_78867[10];
  wire [31:0] add_78868;
  wire [31:0] array_update_78869[10][10];
  wire [31:0] array_index_78871[10];
  wire [31:0] array_index_78872[10];
  wire [31:0] smul_78876;
  wire [31:0] add_78878;
  wire [31:0] array_update_78880[10];
  wire [31:0] add_78881;
  wire [31:0] array_update_78882[10][10];
  wire [31:0] array_index_78884[10];
  wire [31:0] array_index_78885[10];
  wire [31:0] smul_78889;
  wire [31:0] add_78891;
  wire [31:0] array_update_78893[10];
  wire [31:0] add_78894;
  wire [31:0] array_update_78895[10][10];
  wire [31:0] array_index_78897[10];
  wire [31:0] array_index_78898[10];
  wire [31:0] smul_78902;
  wire [31:0] add_78904;
  wire [31:0] array_update_78905[10];
  wire [31:0] array_update_78906[10][10];
  wire [31:0] array_index_78908[10];
  wire [31:0] add_78910;
  wire [31:0] array_update_78911[10];
  wire [31:0] literal_78912;
  wire [31:0] array_update_78913[10][10];
  wire [31:0] array_index_78915[10];
  wire [31:0] array_index_78916[10];
  wire [31:0] smul_78920;
  wire [31:0] add_78922;
  wire [31:0] array_update_78924[10];
  wire [31:0] add_78925;
  wire [31:0] array_update_78926[10][10];
  wire [31:0] array_index_78928[10];
  wire [31:0] array_index_78929[10];
  wire [31:0] smul_78933;
  wire [31:0] add_78935;
  wire [31:0] array_update_78937[10];
  wire [31:0] add_78938;
  wire [31:0] array_update_78939[10][10];
  wire [31:0] array_index_78941[10];
  wire [31:0] array_index_78942[10];
  wire [31:0] smul_78946;
  wire [31:0] add_78948;
  wire [31:0] array_update_78950[10];
  wire [31:0] add_78951;
  wire [31:0] array_update_78952[10][10];
  wire [31:0] array_index_78954[10];
  wire [31:0] array_index_78955[10];
  wire [31:0] smul_78959;
  wire [31:0] add_78961;
  wire [31:0] array_update_78963[10];
  wire [31:0] add_78964;
  wire [31:0] array_update_78965[10][10];
  wire [31:0] array_index_78967[10];
  wire [31:0] array_index_78968[10];
  wire [31:0] smul_78972;
  wire [31:0] add_78974;
  wire [31:0] array_update_78976[10];
  wire [31:0] add_78977;
  wire [31:0] array_update_78978[10][10];
  wire [31:0] array_index_78980[10];
  wire [31:0] array_index_78981[10];
  wire [31:0] smul_78985;
  wire [31:0] add_78987;
  wire [31:0] array_update_78989[10];
  wire [31:0] add_78990;
  wire [31:0] array_update_78991[10][10];
  wire [31:0] array_index_78993[10];
  wire [31:0] array_index_78994[10];
  wire [31:0] smul_78998;
  wire [31:0] add_79000;
  wire [31:0] array_update_79002[10];
  wire [31:0] add_79003;
  wire [31:0] array_update_79004[10][10];
  wire [31:0] array_index_79006[10];
  wire [31:0] array_index_79007[10];
  wire [31:0] smul_79011;
  wire [31:0] add_79013;
  wire [31:0] array_update_79015[10];
  wire [31:0] add_79016;
  wire [31:0] array_update_79017[10][10];
  wire [31:0] array_index_79019[10];
  wire [31:0] array_index_79020[10];
  wire [31:0] smul_79024;
  wire [31:0] add_79026;
  wire [31:0] array_update_79028[10];
  wire [31:0] add_79029;
  wire [31:0] array_update_79030[10][10];
  wire [31:0] array_index_79032[10];
  wire [31:0] array_index_79033[10];
  wire [31:0] smul_79037;
  wire [31:0] add_79039;
  wire [31:0] array_update_79040[10];
  wire [31:0] array_update_79041[10][10];
  wire [31:0] array_index_79043[10];
  wire [31:0] add_79045;
  wire [31:0] array_update_79046[10];
  wire [31:0] literal_79047;
  wire [31:0] array_update_79048[10][10];
  wire [31:0] array_index_79050[10];
  wire [31:0] array_index_79051[10];
  wire [31:0] smul_79055;
  wire [31:0] add_79057;
  wire [31:0] array_update_79059[10];
  wire [31:0] add_79060;
  wire [31:0] array_update_79061[10][10];
  wire [31:0] array_index_79063[10];
  wire [31:0] array_index_79064[10];
  wire [31:0] smul_79068;
  wire [31:0] add_79070;
  wire [31:0] array_update_79072[10];
  wire [31:0] add_79073;
  wire [31:0] array_update_79074[10][10];
  wire [31:0] array_index_79076[10];
  wire [31:0] array_index_79077[10];
  wire [31:0] smul_79081;
  wire [31:0] add_79083;
  wire [31:0] array_update_79085[10];
  wire [31:0] add_79086;
  wire [31:0] array_update_79087[10][10];
  wire [31:0] array_index_79089[10];
  wire [31:0] array_index_79090[10];
  wire [31:0] smul_79094;
  wire [31:0] add_79096;
  wire [31:0] array_update_79098[10];
  wire [31:0] add_79099;
  wire [31:0] array_update_79100[10][10];
  wire [31:0] array_index_79102[10];
  wire [31:0] array_index_79103[10];
  wire [31:0] smul_79107;
  wire [31:0] add_79109;
  wire [31:0] array_update_79111[10];
  wire [31:0] add_79112;
  wire [31:0] array_update_79113[10][10];
  wire [31:0] array_index_79115[10];
  wire [31:0] array_index_79116[10];
  wire [31:0] smul_79120;
  wire [31:0] add_79122;
  wire [31:0] array_update_79124[10];
  wire [31:0] add_79125;
  wire [31:0] array_update_79126[10][10];
  wire [31:0] array_index_79128[10];
  wire [31:0] array_index_79129[10];
  wire [31:0] smul_79133;
  wire [31:0] add_79135;
  wire [31:0] array_update_79137[10];
  wire [31:0] add_79138;
  wire [31:0] array_update_79139[10][10];
  wire [31:0] array_index_79141[10];
  wire [31:0] array_index_79142[10];
  wire [31:0] smul_79146;
  wire [31:0] add_79148;
  wire [31:0] array_update_79150[10];
  wire [31:0] add_79151;
  wire [31:0] array_update_79152[10][10];
  wire [31:0] array_index_79154[10];
  wire [31:0] array_index_79155[10];
  wire [31:0] smul_79159;
  wire [31:0] add_79161;
  wire [31:0] array_update_79163[10];
  wire [31:0] add_79164;
  wire [31:0] array_update_79165[10][10];
  wire [31:0] array_index_79167[10];
  wire [31:0] array_index_79168[10];
  wire [31:0] smul_79172;
  wire [31:0] add_79174;
  wire [31:0] array_update_79175[10];
  wire [31:0] array_update_79176[10][10];
  wire [31:0] array_index_79178[10];
  wire [31:0] add_79180;
  wire [31:0] array_update_79181[10];
  wire [31:0] literal_79182;
  wire [31:0] array_update_79183[10][10];
  wire [31:0] array_index_79185[10];
  wire [31:0] array_index_79186[10];
  wire [31:0] smul_79190;
  wire [31:0] add_79192;
  wire [31:0] array_update_79194[10];
  wire [31:0] add_79195;
  wire [31:0] array_update_79196[10][10];
  wire [31:0] array_index_79198[10];
  wire [31:0] array_index_79199[10];
  wire [31:0] smul_79203;
  wire [31:0] add_79205;
  wire [31:0] array_update_79207[10];
  wire [31:0] add_79208;
  wire [31:0] array_update_79209[10][10];
  wire [31:0] array_index_79211[10];
  wire [31:0] array_index_79212[10];
  wire [31:0] smul_79216;
  wire [31:0] add_79218;
  wire [31:0] array_update_79220[10];
  wire [31:0] add_79221;
  wire [31:0] array_update_79222[10][10];
  wire [31:0] array_index_79224[10];
  wire [31:0] array_index_79225[10];
  wire [31:0] smul_79229;
  wire [31:0] add_79231;
  wire [31:0] array_update_79233[10];
  wire [31:0] add_79234;
  wire [31:0] array_update_79235[10][10];
  wire [31:0] array_index_79237[10];
  wire [31:0] array_index_79238[10];
  wire [31:0] smul_79242;
  wire [31:0] add_79244;
  wire [31:0] array_update_79246[10];
  wire [31:0] add_79247;
  wire [31:0] array_update_79248[10][10];
  wire [31:0] array_index_79250[10];
  wire [31:0] array_index_79251[10];
  wire [31:0] smul_79255;
  wire [31:0] add_79257;
  wire [31:0] array_update_79259[10];
  wire [31:0] add_79260;
  wire [31:0] array_update_79261[10][10];
  wire [31:0] array_index_79263[10];
  wire [31:0] array_index_79264[10];
  wire [31:0] smul_79268;
  wire [31:0] add_79270;
  wire [31:0] array_update_79272[10];
  wire [31:0] add_79273;
  wire [31:0] array_update_79274[10][10];
  wire [31:0] array_index_79276[10];
  wire [31:0] array_index_79277[10];
  wire [31:0] smul_79281;
  wire [31:0] add_79283;
  wire [31:0] array_update_79285[10];
  wire [31:0] add_79286;
  wire [31:0] array_update_79287[10][10];
  wire [31:0] array_index_79289[10];
  wire [31:0] array_index_79290[10];
  wire [31:0] smul_79294;
  wire [31:0] add_79296;
  wire [31:0] array_update_79298[10];
  wire [31:0] add_79299;
  wire [31:0] array_update_79300[10][10];
  wire [31:0] array_index_79302[10];
  wire [31:0] array_index_79303[10];
  wire [31:0] smul_79307;
  wire [31:0] add_79309;
  wire [31:0] array_update_79310[10];
  wire [31:0] array_update_79311[10][10];
  wire [31:0] array_index_79313[10];
  wire [31:0] add_79315;
  wire [31:0] array_update_79316[10];
  wire [31:0] literal_79317;
  wire [31:0] array_update_79318[10][10];
  wire [31:0] array_index_79320[10];
  wire [31:0] array_index_79321[10];
  wire [31:0] smul_79325;
  wire [31:0] add_79327;
  wire [31:0] array_update_79329[10];
  wire [31:0] add_79330;
  wire [31:0] array_update_79331[10][10];
  wire [31:0] array_index_79333[10];
  wire [31:0] array_index_79334[10];
  wire [31:0] smul_79338;
  wire [31:0] add_79340;
  wire [31:0] array_update_79342[10];
  wire [31:0] add_79343;
  wire [31:0] array_update_79344[10][10];
  wire [31:0] array_index_79346[10];
  wire [31:0] array_index_79347[10];
  wire [31:0] smul_79351;
  wire [31:0] add_79353;
  wire [31:0] array_update_79355[10];
  wire [31:0] add_79356;
  wire [31:0] array_update_79357[10][10];
  wire [31:0] array_index_79359[10];
  wire [31:0] array_index_79360[10];
  wire [31:0] smul_79364;
  wire [31:0] add_79366;
  wire [31:0] array_update_79368[10];
  wire [31:0] add_79369;
  wire [31:0] array_update_79370[10][10];
  wire [31:0] array_index_79372[10];
  wire [31:0] array_index_79373[10];
  wire [31:0] smul_79377;
  wire [31:0] add_79379;
  wire [31:0] array_update_79381[10];
  wire [31:0] add_79382;
  wire [31:0] array_update_79383[10][10];
  wire [31:0] array_index_79385[10];
  wire [31:0] array_index_79386[10];
  wire [31:0] smul_79390;
  wire [31:0] add_79392;
  wire [31:0] array_update_79394[10];
  wire [31:0] add_79395;
  wire [31:0] array_update_79396[10][10];
  wire [31:0] array_index_79398[10];
  wire [31:0] array_index_79399[10];
  wire [31:0] smul_79403;
  wire [31:0] add_79405;
  wire [31:0] array_update_79407[10];
  wire [31:0] add_79408;
  wire [31:0] array_update_79409[10][10];
  wire [31:0] array_index_79411[10];
  wire [31:0] array_index_79412[10];
  wire [31:0] smul_79416;
  wire [31:0] add_79418;
  wire [31:0] array_update_79420[10];
  wire [31:0] add_79421;
  wire [31:0] array_update_79422[10][10];
  wire [31:0] array_index_79424[10];
  wire [31:0] array_index_79425[10];
  wire [31:0] smul_79429;
  wire [31:0] add_79431;
  wire [31:0] array_update_79433[10];
  wire [31:0] add_79434;
  wire [31:0] array_update_79435[10][10];
  wire [31:0] array_index_79437[10];
  wire [31:0] array_index_79438[10];
  wire [31:0] smul_79442;
  wire [31:0] add_79444;
  wire [31:0] array_update_79445[10];
  wire [31:0] array_update_79446[10][10];
  wire [31:0] array_index_79448[10];
  wire [31:0] add_79450;
  wire [31:0] array_update_79451[10];
  wire [31:0] literal_79452;
  wire [31:0] array_update_79453[10][10];
  wire [31:0] array_index_79455[10];
  wire [31:0] array_index_79456[10];
  wire [31:0] smul_79460;
  wire [31:0] add_79462;
  wire [31:0] array_update_79464[10];
  wire [31:0] add_79465;
  wire [31:0] array_update_79466[10][10];
  wire [31:0] array_index_79468[10];
  wire [31:0] array_index_79469[10];
  wire [31:0] smul_79473;
  wire [31:0] add_79475;
  wire [31:0] array_update_79477[10];
  wire [31:0] add_79478;
  wire [31:0] array_update_79479[10][10];
  wire [31:0] array_index_79481[10];
  wire [31:0] array_index_79482[10];
  wire [31:0] smul_79486;
  wire [31:0] add_79488;
  wire [31:0] array_update_79490[10];
  wire [31:0] add_79491;
  wire [31:0] array_update_79492[10][10];
  wire [31:0] array_index_79494[10];
  wire [31:0] array_index_79495[10];
  wire [31:0] smul_79499;
  wire [31:0] add_79501;
  wire [31:0] array_update_79503[10];
  wire [31:0] add_79504;
  wire [31:0] array_update_79505[10][10];
  wire [31:0] array_index_79507[10];
  wire [31:0] array_index_79508[10];
  wire [31:0] smul_79512;
  wire [31:0] add_79514;
  wire [31:0] array_update_79516[10];
  wire [31:0] add_79517;
  wire [31:0] array_update_79518[10][10];
  wire [31:0] array_index_79520[10];
  wire [31:0] array_index_79521[10];
  wire [31:0] smul_79525;
  wire [31:0] add_79527;
  wire [31:0] array_update_79529[10];
  wire [31:0] add_79530;
  wire [31:0] array_update_79531[10][10];
  wire [31:0] array_index_79533[10];
  wire [31:0] array_index_79534[10];
  wire [31:0] smul_79538;
  wire [31:0] add_79540;
  wire [31:0] array_update_79542[10];
  wire [31:0] add_79543;
  wire [31:0] array_update_79544[10][10];
  wire [31:0] array_index_79546[10];
  wire [31:0] array_index_79547[10];
  wire [31:0] smul_79551;
  wire [31:0] add_79553;
  wire [31:0] array_update_79555[10];
  wire [31:0] add_79556;
  wire [31:0] array_update_79557[10][10];
  wire [31:0] array_index_79559[10];
  wire [31:0] array_index_79560[10];
  wire [31:0] smul_79564;
  wire [31:0] add_79566;
  wire [31:0] array_update_79568[10];
  wire [31:0] add_79569;
  wire [31:0] array_update_79570[10][10];
  wire [31:0] array_index_79572[10];
  wire [31:0] array_index_79573[10];
  wire [31:0] smul_79577;
  wire [31:0] add_79579;
  wire [31:0] array_update_79580[10];
  wire [31:0] array_update_79581[10][10];
  wire [31:0] array_index_79583[10];
  wire [31:0] add_79585;
  wire [31:0] array_update_79586[10];
  wire [31:0] literal_79587;
  wire [31:0] array_update_79588[10][10];
  wire [31:0] array_index_79590[10];
  wire [31:0] array_index_79591[10];
  wire [31:0] smul_79595;
  wire [31:0] add_79597;
  wire [31:0] array_update_79599[10];
  wire [31:0] add_79600;
  wire [31:0] array_update_79601[10][10];
  wire [31:0] array_index_79603[10];
  wire [31:0] array_index_79604[10];
  wire [31:0] smul_79608;
  wire [31:0] add_79610;
  wire [31:0] array_update_79612[10];
  wire [31:0] add_79613;
  wire [31:0] array_update_79614[10][10];
  wire [31:0] array_index_79616[10];
  wire [31:0] array_index_79617[10];
  wire [31:0] smul_79621;
  wire [31:0] add_79623;
  wire [31:0] array_update_79625[10];
  wire [31:0] add_79626;
  wire [31:0] array_update_79627[10][10];
  wire [31:0] array_index_79629[10];
  wire [31:0] array_index_79630[10];
  wire [31:0] smul_79634;
  wire [31:0] add_79636;
  wire [31:0] array_update_79638[10];
  wire [31:0] add_79639;
  wire [31:0] array_update_79640[10][10];
  wire [31:0] array_index_79642[10];
  wire [31:0] array_index_79643[10];
  wire [31:0] smul_79647;
  wire [31:0] add_79649;
  wire [31:0] array_update_79651[10];
  wire [31:0] add_79652;
  wire [31:0] array_update_79653[10][10];
  wire [31:0] array_index_79655[10];
  wire [31:0] array_index_79656[10];
  wire [31:0] smul_79660;
  wire [31:0] add_79662;
  wire [31:0] array_update_79664[10];
  wire [31:0] add_79665;
  wire [31:0] array_update_79666[10][10];
  wire [31:0] array_index_79668[10];
  wire [31:0] array_index_79669[10];
  wire [31:0] smul_79673;
  wire [31:0] add_79675;
  wire [31:0] array_update_79677[10];
  wire [31:0] add_79678;
  wire [31:0] array_update_79679[10][10];
  wire [31:0] array_index_79681[10];
  wire [31:0] array_index_79682[10];
  wire [31:0] smul_79686;
  wire [31:0] add_79688;
  wire [31:0] array_update_79690[10];
  wire [31:0] add_79691;
  wire [31:0] array_update_79692[10][10];
  wire [31:0] array_index_79694[10];
  wire [31:0] array_index_79695[10];
  wire [31:0] smul_79699;
  wire [31:0] add_79701;
  wire [31:0] array_update_79703[10];
  wire [31:0] add_79704;
  wire [31:0] array_update_79705[10][10];
  wire [31:0] array_index_79707[10];
  wire [31:0] array_index_79708[10];
  wire [31:0] smul_79712;
  wire [31:0] add_79714;
  wire [31:0] array_update_79715[10];
  wire [31:0] array_update_79716[10][10];
  wire [31:0] array_index_79718[10];
  wire [31:0] add_79720;
  wire [31:0] array_update_79721[10];
  wire [31:0] literal_79722;
  wire [31:0] array_update_79723[10][10];
  wire [31:0] array_index_79725[10];
  wire [31:0] array_index_79726[10];
  wire [31:0] smul_79730;
  wire [31:0] add_79732;
  wire [31:0] array_update_79734[10];
  wire [31:0] add_79735;
  wire [31:0] array_update_79736[10][10];
  wire [31:0] array_index_79738[10];
  wire [31:0] array_index_79739[10];
  wire [31:0] smul_79743;
  wire [31:0] add_79745;
  wire [31:0] array_update_79747[10];
  wire [31:0] add_79748;
  wire [31:0] array_update_79749[10][10];
  wire [31:0] array_index_79751[10];
  wire [31:0] array_index_79752[10];
  wire [31:0] smul_79756;
  wire [31:0] add_79758;
  wire [31:0] array_update_79760[10];
  wire [31:0] add_79761;
  wire [31:0] array_update_79762[10][10];
  wire [31:0] array_index_79764[10];
  wire [31:0] array_index_79765[10];
  wire [31:0] smul_79769;
  wire [31:0] add_79771;
  wire [31:0] array_update_79773[10];
  wire [31:0] add_79774;
  wire [31:0] array_update_79775[10][10];
  wire [31:0] array_index_79777[10];
  wire [31:0] array_index_79778[10];
  wire [31:0] smul_79782;
  wire [31:0] add_79784;
  wire [31:0] array_update_79786[10];
  wire [31:0] add_79787;
  wire [31:0] array_update_79788[10][10];
  wire [31:0] array_index_79790[10];
  wire [31:0] array_index_79791[10];
  wire [31:0] smul_79795;
  wire [31:0] add_79797;
  wire [31:0] array_update_79799[10];
  wire [31:0] add_79800;
  wire [31:0] array_update_79801[10][10];
  wire [31:0] array_index_79803[10];
  wire [31:0] array_index_79804[10];
  wire [31:0] smul_79808;
  wire [31:0] add_79810;
  wire [31:0] array_update_79812[10];
  wire [31:0] add_79813;
  wire [31:0] array_update_79814[10][10];
  wire [31:0] array_index_79816[10];
  wire [31:0] array_index_79817[10];
  wire [31:0] smul_79821;
  wire [31:0] add_79823;
  wire [31:0] array_update_79825[10];
  wire [31:0] add_79826;
  wire [31:0] array_update_79827[10][10];
  wire [31:0] array_index_79829[10];
  wire [31:0] array_index_79830[10];
  wire [31:0] smul_79834;
  wire [31:0] add_79836;
  wire [31:0] array_update_79838[10];
  wire [31:0] add_79839;
  wire [31:0] array_update_79840[10][10];
  wire [31:0] array_index_79842[10];
  wire [31:0] array_index_79843[10];
  wire [31:0] smul_79847;
  wire [31:0] add_79849;
  wire [31:0] array_update_79850[10];
  wire [31:0] array_update_79851[10][10];
  wire [31:0] array_index_79853[10];
  wire [31:0] add_79855;
  wire [31:0] array_update_79856[10];
  wire [31:0] literal_79857;
  wire [31:0] array_update_79858[10][10];
  wire [31:0] array_index_79860[10];
  wire [31:0] array_index_79861[10];
  wire [31:0] smul_79865;
  wire [31:0] add_79867;
  wire [31:0] array_update_79869[10];
  wire [31:0] add_79870;
  wire [31:0] array_update_79871[10][10];
  wire [31:0] array_index_79873[10];
  wire [31:0] array_index_79874[10];
  wire [31:0] smul_79878;
  wire [31:0] add_79880;
  wire [31:0] array_update_79882[10];
  wire [31:0] add_79883;
  wire [31:0] array_update_79884[10][10];
  wire [31:0] array_index_79886[10];
  wire [31:0] array_index_79887[10];
  wire [31:0] smul_79891;
  wire [31:0] add_79893;
  wire [31:0] array_update_79895[10];
  wire [31:0] add_79896;
  wire [31:0] array_update_79897[10][10];
  wire [31:0] array_index_79899[10];
  wire [31:0] array_index_79900[10];
  wire [31:0] smul_79904;
  wire [31:0] add_79906;
  wire [31:0] array_update_79908[10];
  wire [31:0] add_79909;
  wire [31:0] array_update_79910[10][10];
  wire [31:0] array_index_79912[10];
  wire [31:0] array_index_79913[10];
  wire [31:0] smul_79917;
  wire [31:0] add_79919;
  wire [31:0] array_update_79921[10];
  wire [31:0] add_79922;
  wire [31:0] array_update_79923[10][10];
  wire [31:0] array_index_79925[10];
  wire [31:0] array_index_79926[10];
  wire [31:0] smul_79930;
  wire [31:0] add_79932;
  wire [31:0] array_update_79934[10];
  wire [31:0] add_79935;
  wire [31:0] array_update_79936[10][10];
  wire [31:0] array_index_79938[10];
  wire [31:0] array_index_79939[10];
  wire [31:0] smul_79943;
  wire [31:0] add_79945;
  wire [31:0] array_update_79947[10];
  wire [31:0] add_79948;
  wire [31:0] array_update_79949[10][10];
  wire [31:0] array_index_79951[10];
  wire [31:0] array_index_79952[10];
  wire [31:0] smul_79956;
  wire [31:0] add_79958;
  wire [31:0] array_update_79960[10];
  wire [31:0] add_79961;
  wire [31:0] array_update_79962[10][10];
  wire [31:0] array_index_79964[10];
  wire [31:0] array_index_79965[10];
  wire [31:0] smul_79969;
  wire [31:0] add_79971;
  wire [31:0] array_update_79973[10];
  wire [31:0] add_79974;
  wire [31:0] array_update_79975[10][10];
  wire [31:0] array_index_79977[10];
  wire [31:0] array_index_79978[10];
  wire [31:0] smul_79982;
  wire [31:0] add_79984;
  wire [31:0] array_update_79985[10];
  wire [31:0] array_update_79986[10][10];
  wire [31:0] array_index_79988[10];
  wire [31:0] add_79990;
  wire [31:0] array_update_79991[10];
  wire [31:0] literal_79992;
  wire [31:0] array_update_79993[10][10];
  wire [31:0] array_index_79995[10];
  wire [31:0] array_index_79996[10];
  wire [31:0] smul_80000;
  wire [31:0] add_80002;
  wire [31:0] array_update_80004[10];
  wire [31:0] add_80005;
  wire [31:0] array_update_80006[10][10];
  wire [31:0] array_index_80008[10];
  wire [31:0] array_index_80009[10];
  wire [31:0] smul_80013;
  wire [31:0] add_80015;
  wire [31:0] array_update_80017[10];
  wire [31:0] add_80018;
  wire [31:0] array_update_80019[10][10];
  wire [31:0] array_index_80021[10];
  wire [31:0] array_index_80022[10];
  wire [31:0] smul_80026;
  wire [31:0] add_80028;
  wire [31:0] array_update_80030[10];
  wire [31:0] add_80031;
  wire [31:0] array_update_80032[10][10];
  wire [31:0] array_index_80034[10];
  wire [31:0] array_index_80035[10];
  wire [31:0] smul_80039;
  wire [31:0] add_80041;
  wire [31:0] array_update_80043[10];
  wire [31:0] add_80044;
  wire [31:0] array_update_80045[10][10];
  wire [31:0] array_index_80047[10];
  wire [31:0] array_index_80048[10];
  wire [31:0] smul_80052;
  wire [31:0] add_80054;
  wire [31:0] array_update_80056[10];
  wire [31:0] add_80057;
  wire [31:0] array_update_80058[10][10];
  wire [31:0] array_index_80060[10];
  wire [31:0] array_index_80061[10];
  wire [31:0] smul_80065;
  wire [31:0] add_80067;
  wire [31:0] array_update_80069[10];
  wire [31:0] add_80070;
  wire [31:0] array_update_80071[10][10];
  wire [31:0] array_index_80073[10];
  wire [31:0] array_index_80074[10];
  wire [31:0] smul_80078;
  wire [31:0] add_80080;
  wire [31:0] array_update_80082[10];
  wire [31:0] add_80083;
  wire [31:0] array_update_80084[10][10];
  wire [31:0] array_index_80086[10];
  wire [31:0] array_index_80087[10];
  wire [31:0] smul_80091;
  wire [31:0] add_80093;
  wire [31:0] array_update_80095[10];
  wire [31:0] add_80096;
  wire [31:0] array_update_80097[10][10];
  wire [31:0] array_index_80099[10];
  wire [31:0] array_index_80100[10];
  wire [31:0] smul_80104;
  wire [31:0] add_80106;
  wire [31:0] array_update_80108[10];
  wire [31:0] add_80109;
  wire [31:0] array_update_80110[10][10];
  wire [31:0] array_index_80112[10];
  wire [31:0] array_index_80113[10];
  wire [31:0] smul_80117;
  wire [31:0] add_80119;
  wire [31:0] array_update_80120[10];
  wire [31:0] array_update_80122[10][10];
  wire [31:0] add_80123;
  wire [31:0] array_index_80124[10];
  wire [31:0] literal_80126;
  wire [31:0] array_update_80127[10];
  wire [31:0] literal_80128;
  wire [31:0] array_update_80129[10][10];
  wire [31:0] array_index_80130[10];
  wire [31:0] array_index_80131[10];
  wire [31:0] array_index_80132[10];
  wire [31:0] smul_80136;
  wire [31:0] add_80138;
  wire [31:0] array_update_80140[10];
  wire [31:0] add_80141;
  wire [31:0] array_update_80142[10][10];
  wire [31:0] array_index_80144[10];
  wire [31:0] array_index_80145[10];
  wire [31:0] smul_80149;
  wire [31:0] add_80151;
  wire [31:0] array_update_80153[10];
  wire [31:0] add_80154;
  wire [31:0] array_update_80155[10][10];
  wire [31:0] array_index_80157[10];
  wire [31:0] array_index_80158[10];
  wire [31:0] smul_80162;
  wire [31:0] add_80164;
  wire [31:0] array_update_80166[10];
  wire [31:0] add_80167;
  wire [31:0] array_update_80168[10][10];
  wire [31:0] array_index_80170[10];
  wire [31:0] array_index_80171[10];
  wire [31:0] smul_80175;
  wire [31:0] add_80177;
  wire [31:0] array_update_80179[10];
  wire [31:0] add_80180;
  wire [31:0] array_update_80181[10][10];
  wire [31:0] array_index_80183[10];
  wire [31:0] array_index_80184[10];
  wire [31:0] smul_80188;
  wire [31:0] add_80190;
  wire [31:0] array_update_80192[10];
  wire [31:0] add_80193;
  wire [31:0] array_update_80194[10][10];
  wire [31:0] array_index_80196[10];
  wire [31:0] array_index_80197[10];
  wire [31:0] smul_80201;
  wire [31:0] add_80203;
  wire [31:0] array_update_80205[10];
  wire [31:0] add_80206;
  wire [31:0] array_update_80207[10][10];
  wire [31:0] array_index_80209[10];
  wire [31:0] array_index_80210[10];
  wire [31:0] smul_80214;
  wire [31:0] add_80216;
  wire [31:0] array_update_80218[10];
  wire [31:0] add_80219;
  wire [31:0] array_update_80220[10][10];
  wire [31:0] array_index_80222[10];
  wire [31:0] array_index_80223[10];
  wire [31:0] smul_80227;
  wire [31:0] add_80229;
  wire [31:0] array_update_80231[10];
  wire [31:0] add_80232;
  wire [31:0] array_update_80233[10][10];
  wire [31:0] array_index_80235[10];
  wire [31:0] array_index_80236[10];
  wire [31:0] smul_80240;
  wire [31:0] add_80242;
  wire [31:0] array_update_80244[10];
  wire [31:0] add_80245;
  wire [31:0] array_update_80246[10][10];
  wire [31:0] array_index_80248[10];
  wire [31:0] array_index_80249[10];
  wire [31:0] smul_80253;
  wire [31:0] add_80255;
  wire [31:0] array_update_80256[10];
  wire [31:0] array_update_80257[10][10];
  wire [31:0] array_index_80259[10];
  wire [31:0] add_80261;
  wire [31:0] array_update_80262[10];
  wire [31:0] literal_80263;
  wire [31:0] array_update_80264[10][10];
  wire [31:0] array_index_80266[10];
  wire [31:0] array_index_80267[10];
  wire [31:0] smul_80271;
  wire [31:0] add_80273;
  wire [31:0] array_update_80275[10];
  wire [31:0] add_80276;
  wire [31:0] array_update_80277[10][10];
  wire [31:0] array_index_80279[10];
  wire [31:0] array_index_80280[10];
  wire [31:0] smul_80284;
  wire [31:0] add_80286;
  wire [31:0] array_update_80288[10];
  wire [31:0] add_80289;
  wire [31:0] array_update_80290[10][10];
  wire [31:0] array_index_80292[10];
  wire [31:0] array_index_80293[10];
  wire [31:0] smul_80297;
  wire [31:0] add_80299;
  wire [31:0] array_update_80301[10];
  wire [31:0] add_80302;
  wire [31:0] array_update_80303[10][10];
  wire [31:0] array_index_80305[10];
  wire [31:0] array_index_80306[10];
  wire [31:0] smul_80310;
  wire [31:0] add_80312;
  wire [31:0] array_update_80314[10];
  wire [31:0] add_80315;
  wire [31:0] array_update_80316[10][10];
  wire [31:0] array_index_80318[10];
  wire [31:0] array_index_80319[10];
  wire [31:0] smul_80323;
  wire [31:0] add_80325;
  wire [31:0] array_update_80327[10];
  wire [31:0] add_80328;
  wire [31:0] array_update_80329[10][10];
  wire [31:0] array_index_80331[10];
  wire [31:0] array_index_80332[10];
  wire [31:0] smul_80336;
  wire [31:0] add_80338;
  wire [31:0] array_update_80340[10];
  wire [31:0] add_80341;
  wire [31:0] array_update_80342[10][10];
  wire [31:0] array_index_80344[10];
  wire [31:0] array_index_80345[10];
  wire [31:0] smul_80349;
  wire [31:0] add_80351;
  wire [31:0] array_update_80353[10];
  wire [31:0] add_80354;
  wire [31:0] array_update_80355[10][10];
  wire [31:0] array_index_80357[10];
  wire [31:0] array_index_80358[10];
  wire [31:0] smul_80362;
  wire [31:0] add_80364;
  wire [31:0] array_update_80366[10];
  wire [31:0] add_80367;
  wire [31:0] array_update_80368[10][10];
  wire [31:0] array_index_80370[10];
  wire [31:0] array_index_80371[10];
  wire [31:0] smul_80375;
  wire [31:0] add_80377;
  wire [31:0] array_update_80379[10];
  wire [31:0] add_80380;
  wire [31:0] array_update_80381[10][10];
  wire [31:0] array_index_80383[10];
  wire [31:0] array_index_80384[10];
  wire [31:0] smul_80388;
  wire [31:0] add_80390;
  wire [31:0] array_update_80391[10];
  wire [31:0] array_update_80392[10][10];
  wire [31:0] array_index_80394[10];
  wire [31:0] add_80396;
  wire [31:0] array_update_80397[10];
  wire [31:0] literal_80398;
  wire [31:0] array_update_80399[10][10];
  wire [31:0] array_index_80401[10];
  wire [31:0] array_index_80402[10];
  wire [31:0] smul_80406;
  wire [31:0] add_80408;
  wire [31:0] array_update_80410[10];
  wire [31:0] add_80411;
  wire [31:0] array_update_80412[10][10];
  wire [31:0] array_index_80414[10];
  wire [31:0] array_index_80415[10];
  wire [31:0] smul_80419;
  wire [31:0] add_80421;
  wire [31:0] array_update_80423[10];
  wire [31:0] add_80424;
  wire [31:0] array_update_80425[10][10];
  wire [31:0] array_index_80427[10];
  wire [31:0] array_index_80428[10];
  wire [31:0] smul_80432;
  wire [31:0] add_80434;
  wire [31:0] array_update_80436[10];
  wire [31:0] add_80437;
  wire [31:0] array_update_80438[10][10];
  wire [31:0] array_index_80440[10];
  wire [31:0] array_index_80441[10];
  wire [31:0] smul_80445;
  wire [31:0] add_80447;
  wire [31:0] array_update_80449[10];
  wire [31:0] add_80450;
  wire [31:0] array_update_80451[10][10];
  wire [31:0] array_index_80453[10];
  wire [31:0] array_index_80454[10];
  wire [31:0] smul_80458;
  wire [31:0] add_80460;
  wire [31:0] array_update_80462[10];
  wire [31:0] add_80463;
  wire [31:0] array_update_80464[10][10];
  wire [31:0] array_index_80466[10];
  wire [31:0] array_index_80467[10];
  wire [31:0] smul_80471;
  wire [31:0] add_80473;
  wire [31:0] array_update_80475[10];
  wire [31:0] add_80476;
  wire [31:0] array_update_80477[10][10];
  wire [31:0] array_index_80479[10];
  wire [31:0] array_index_80480[10];
  wire [31:0] smul_80484;
  wire [31:0] add_80486;
  wire [31:0] array_update_80488[10];
  wire [31:0] add_80489;
  wire [31:0] array_update_80490[10][10];
  wire [31:0] array_index_80492[10];
  wire [31:0] array_index_80493[10];
  wire [31:0] smul_80497;
  wire [31:0] add_80499;
  wire [31:0] array_update_80501[10];
  wire [31:0] add_80502;
  wire [31:0] array_update_80503[10][10];
  wire [31:0] array_index_80505[10];
  wire [31:0] array_index_80506[10];
  wire [31:0] smul_80510;
  wire [31:0] add_80512;
  wire [31:0] array_update_80514[10];
  wire [31:0] add_80515;
  wire [31:0] array_update_80516[10][10];
  wire [31:0] array_index_80518[10];
  wire [31:0] array_index_80519[10];
  wire [31:0] smul_80523;
  wire [31:0] add_80525;
  wire [31:0] array_update_80526[10];
  wire [31:0] array_update_80527[10][10];
  wire [31:0] array_index_80529[10];
  wire [31:0] add_80531;
  wire [31:0] array_update_80532[10];
  wire [31:0] literal_80533;
  wire [31:0] array_update_80534[10][10];
  wire [31:0] array_index_80536[10];
  wire [31:0] array_index_80537[10];
  wire [31:0] smul_80541;
  wire [31:0] add_80543;
  wire [31:0] array_update_80545[10];
  wire [31:0] add_80546;
  wire [31:0] array_update_80547[10][10];
  wire [31:0] array_index_80549[10];
  wire [31:0] array_index_80550[10];
  wire [31:0] smul_80554;
  wire [31:0] add_80556;
  wire [31:0] array_update_80558[10];
  wire [31:0] add_80559;
  wire [31:0] array_update_80560[10][10];
  wire [31:0] array_index_80562[10];
  wire [31:0] array_index_80563[10];
  wire [31:0] smul_80567;
  wire [31:0] add_80569;
  wire [31:0] array_update_80571[10];
  wire [31:0] add_80572;
  wire [31:0] array_update_80573[10][10];
  wire [31:0] array_index_80575[10];
  wire [31:0] array_index_80576[10];
  wire [31:0] smul_80580;
  wire [31:0] add_80582;
  wire [31:0] array_update_80584[10];
  wire [31:0] add_80585;
  wire [31:0] array_update_80586[10][10];
  wire [31:0] array_index_80588[10];
  wire [31:0] array_index_80589[10];
  wire [31:0] smul_80593;
  wire [31:0] add_80595;
  wire [31:0] array_update_80597[10];
  wire [31:0] add_80598;
  wire [31:0] array_update_80599[10][10];
  wire [31:0] array_index_80601[10];
  wire [31:0] array_index_80602[10];
  wire [31:0] smul_80606;
  wire [31:0] add_80608;
  wire [31:0] array_update_80610[10];
  wire [31:0] add_80611;
  wire [31:0] array_update_80612[10][10];
  wire [31:0] array_index_80614[10];
  wire [31:0] array_index_80615[10];
  wire [31:0] smul_80619;
  wire [31:0] add_80621;
  wire [31:0] array_update_80623[10];
  wire [31:0] add_80624;
  wire [31:0] array_update_80625[10][10];
  wire [31:0] array_index_80627[10];
  wire [31:0] array_index_80628[10];
  wire [31:0] smul_80632;
  wire [31:0] add_80634;
  wire [31:0] array_update_80636[10];
  wire [31:0] add_80637;
  wire [31:0] array_update_80638[10][10];
  wire [31:0] array_index_80640[10];
  wire [31:0] array_index_80641[10];
  wire [31:0] smul_80645;
  wire [31:0] add_80647;
  wire [31:0] array_update_80649[10];
  wire [31:0] add_80650;
  wire [31:0] array_update_80651[10][10];
  wire [31:0] array_index_80653[10];
  wire [31:0] array_index_80654[10];
  wire [31:0] smul_80658;
  wire [31:0] add_80660;
  wire [31:0] array_update_80661[10];
  wire [31:0] array_update_80662[10][10];
  wire [31:0] array_index_80664[10];
  wire [31:0] add_80666;
  wire [31:0] array_update_80667[10];
  wire [31:0] literal_80668;
  wire [31:0] array_update_80669[10][10];
  wire [31:0] array_index_80671[10];
  wire [31:0] array_index_80672[10];
  wire [31:0] smul_80676;
  wire [31:0] add_80678;
  wire [31:0] array_update_80680[10];
  wire [31:0] add_80681;
  wire [31:0] array_update_80682[10][10];
  wire [31:0] array_index_80684[10];
  wire [31:0] array_index_80685[10];
  wire [31:0] smul_80689;
  wire [31:0] add_80691;
  wire [31:0] array_update_80693[10];
  wire [31:0] add_80694;
  wire [31:0] array_update_80695[10][10];
  wire [31:0] array_index_80697[10];
  wire [31:0] array_index_80698[10];
  wire [31:0] smul_80702;
  wire [31:0] add_80704;
  wire [31:0] array_update_80706[10];
  wire [31:0] add_80707;
  wire [31:0] array_update_80708[10][10];
  wire [31:0] array_index_80710[10];
  wire [31:0] array_index_80711[10];
  wire [31:0] smul_80715;
  wire [31:0] add_80717;
  wire [31:0] array_update_80719[10];
  wire [31:0] add_80720;
  wire [31:0] array_update_80721[10][10];
  wire [31:0] array_index_80723[10];
  wire [31:0] array_index_80724[10];
  wire [31:0] smul_80728;
  wire [31:0] add_80730;
  wire [31:0] array_update_80732[10];
  wire [31:0] add_80733;
  wire [31:0] array_update_80734[10][10];
  wire [31:0] array_index_80736[10];
  wire [31:0] array_index_80737[10];
  wire [31:0] smul_80741;
  wire [31:0] add_80743;
  wire [31:0] array_update_80745[10];
  wire [31:0] add_80746;
  wire [31:0] array_update_80747[10][10];
  wire [31:0] array_index_80749[10];
  wire [31:0] array_index_80750[10];
  wire [31:0] smul_80754;
  wire [31:0] add_80756;
  wire [31:0] array_update_80758[10];
  wire [31:0] add_80759;
  wire [31:0] array_update_80760[10][10];
  wire [31:0] array_index_80762[10];
  wire [31:0] array_index_80763[10];
  wire [31:0] smul_80767;
  wire [31:0] add_80769;
  wire [31:0] array_update_80771[10];
  wire [31:0] add_80772;
  wire [31:0] array_update_80773[10][10];
  wire [31:0] array_index_80775[10];
  wire [31:0] array_index_80776[10];
  wire [31:0] smul_80780;
  wire [31:0] add_80782;
  wire [31:0] array_update_80784[10];
  wire [31:0] add_80785;
  wire [31:0] array_update_80786[10][10];
  wire [31:0] array_index_80788[10];
  wire [31:0] array_index_80789[10];
  wire [31:0] smul_80793;
  wire [31:0] add_80795;
  wire [31:0] array_update_80796[10];
  wire [31:0] array_update_80797[10][10];
  wire [31:0] array_index_80799[10];
  wire [31:0] add_80801;
  wire [31:0] array_update_80802[10];
  wire [31:0] literal_80803;
  wire [31:0] array_update_80804[10][10];
  wire [31:0] array_index_80806[10];
  wire [31:0] array_index_80807[10];
  wire [31:0] smul_80811;
  wire [31:0] add_80813;
  wire [31:0] array_update_80815[10];
  wire [31:0] add_80816;
  wire [31:0] array_update_80817[10][10];
  wire [31:0] array_index_80819[10];
  wire [31:0] array_index_80820[10];
  wire [31:0] smul_80824;
  wire [31:0] add_80826;
  wire [31:0] array_update_80828[10];
  wire [31:0] add_80829;
  wire [31:0] array_update_80830[10][10];
  wire [31:0] array_index_80832[10];
  wire [31:0] array_index_80833[10];
  wire [31:0] smul_80837;
  wire [31:0] add_80839;
  wire [31:0] array_update_80841[10];
  wire [31:0] add_80842;
  wire [31:0] array_update_80843[10][10];
  wire [31:0] array_index_80845[10];
  wire [31:0] array_index_80846[10];
  wire [31:0] smul_80850;
  wire [31:0] add_80852;
  wire [31:0] array_update_80854[10];
  wire [31:0] add_80855;
  wire [31:0] array_update_80856[10][10];
  wire [31:0] array_index_80858[10];
  wire [31:0] array_index_80859[10];
  wire [31:0] smul_80863;
  wire [31:0] add_80865;
  wire [31:0] array_update_80867[10];
  wire [31:0] add_80868;
  wire [31:0] array_update_80869[10][10];
  wire [31:0] array_index_80871[10];
  wire [31:0] array_index_80872[10];
  wire [31:0] smul_80876;
  wire [31:0] add_80878;
  wire [31:0] array_update_80880[10];
  wire [31:0] add_80881;
  wire [31:0] array_update_80882[10][10];
  wire [31:0] array_index_80884[10];
  wire [31:0] array_index_80885[10];
  wire [31:0] smul_80889;
  wire [31:0] add_80891;
  wire [31:0] array_update_80893[10];
  wire [31:0] add_80894;
  wire [31:0] array_update_80895[10][10];
  wire [31:0] array_index_80897[10];
  wire [31:0] array_index_80898[10];
  wire [31:0] smul_80902;
  wire [31:0] add_80904;
  wire [31:0] array_update_80906[10];
  wire [31:0] add_80907;
  wire [31:0] array_update_80908[10][10];
  wire [31:0] array_index_80910[10];
  wire [31:0] array_index_80911[10];
  wire [31:0] smul_80915;
  wire [31:0] add_80917;
  wire [31:0] array_update_80919[10];
  wire [31:0] add_80920;
  wire [31:0] array_update_80921[10][10];
  wire [31:0] array_index_80923[10];
  wire [31:0] array_index_80924[10];
  wire [31:0] smul_80928;
  wire [31:0] add_80930;
  wire [31:0] array_update_80931[10];
  wire [31:0] array_update_80932[10][10];
  wire [31:0] array_index_80934[10];
  wire [31:0] add_80936;
  wire [31:0] array_update_80937[10];
  wire [31:0] literal_80938;
  wire [31:0] array_update_80939[10][10];
  wire [31:0] array_index_80941[10];
  wire [31:0] array_index_80942[10];
  wire [31:0] smul_80946;
  wire [31:0] add_80948;
  wire [31:0] array_update_80950[10];
  wire [31:0] add_80951;
  wire [31:0] array_update_80952[10][10];
  wire [31:0] array_index_80954[10];
  wire [31:0] array_index_80955[10];
  wire [31:0] smul_80959;
  wire [31:0] add_80961;
  wire [31:0] array_update_80963[10];
  wire [31:0] add_80964;
  wire [31:0] array_update_80965[10][10];
  wire [31:0] array_index_80967[10];
  wire [31:0] array_index_80968[10];
  wire [31:0] smul_80972;
  wire [31:0] add_80974;
  wire [31:0] array_update_80976[10];
  wire [31:0] add_80977;
  wire [31:0] array_update_80978[10][10];
  wire [31:0] array_index_80980[10];
  wire [31:0] array_index_80981[10];
  wire [31:0] smul_80985;
  wire [31:0] add_80987;
  wire [31:0] array_update_80989[10];
  wire [31:0] add_80990;
  wire [31:0] array_update_80991[10][10];
  wire [31:0] array_index_80993[10];
  wire [31:0] array_index_80994[10];
  wire [31:0] smul_80998;
  wire [31:0] add_81000;
  wire [31:0] array_update_81002[10];
  wire [31:0] add_81003;
  wire [31:0] array_update_81004[10][10];
  wire [31:0] array_index_81006[10];
  wire [31:0] array_index_81007[10];
  wire [31:0] smul_81011;
  wire [31:0] add_81013;
  wire [31:0] array_update_81015[10];
  wire [31:0] add_81016;
  wire [31:0] array_update_81017[10][10];
  wire [31:0] array_index_81019[10];
  wire [31:0] array_index_81020[10];
  wire [31:0] smul_81024;
  wire [31:0] add_81026;
  wire [31:0] array_update_81028[10];
  wire [31:0] add_81029;
  wire [31:0] array_update_81030[10][10];
  wire [31:0] array_index_81032[10];
  wire [31:0] array_index_81033[10];
  wire [31:0] smul_81037;
  wire [31:0] add_81039;
  wire [31:0] array_update_81041[10];
  wire [31:0] add_81042;
  wire [31:0] array_update_81043[10][10];
  wire [31:0] array_index_81045[10];
  wire [31:0] array_index_81046[10];
  wire [31:0] smul_81050;
  wire [31:0] add_81052;
  wire [31:0] array_update_81054[10];
  wire [31:0] add_81055;
  wire [31:0] array_update_81056[10][10];
  wire [31:0] array_index_81058[10];
  wire [31:0] array_index_81059[10];
  wire [31:0] smul_81063;
  wire [31:0] add_81065;
  wire [31:0] array_update_81066[10];
  wire [31:0] array_update_81067[10][10];
  wire [31:0] array_index_81069[10];
  wire [31:0] add_81071;
  wire [31:0] array_update_81072[10];
  wire [31:0] literal_81073;
  wire [31:0] array_update_81074[10][10];
  wire [31:0] array_index_81076[10];
  wire [31:0] array_index_81077[10];
  wire [31:0] smul_81081;
  wire [31:0] add_81083;
  wire [31:0] array_update_81085[10];
  wire [31:0] add_81086;
  wire [31:0] array_update_81087[10][10];
  wire [31:0] array_index_81089[10];
  wire [31:0] array_index_81090[10];
  wire [31:0] smul_81094;
  wire [31:0] add_81096;
  wire [31:0] array_update_81098[10];
  wire [31:0] add_81099;
  wire [31:0] array_update_81100[10][10];
  wire [31:0] array_index_81102[10];
  wire [31:0] array_index_81103[10];
  wire [31:0] smul_81107;
  wire [31:0] add_81109;
  wire [31:0] array_update_81111[10];
  wire [31:0] add_81112;
  wire [31:0] array_update_81113[10][10];
  wire [31:0] array_index_81115[10];
  wire [31:0] array_index_81116[10];
  wire [31:0] smul_81120;
  wire [31:0] add_81122;
  wire [31:0] array_update_81124[10];
  wire [31:0] add_81125;
  wire [31:0] array_update_81126[10][10];
  wire [31:0] array_index_81128[10];
  wire [31:0] array_index_81129[10];
  wire [31:0] smul_81133;
  wire [31:0] add_81135;
  wire [31:0] array_update_81137[10];
  wire [31:0] add_81138;
  wire [31:0] array_update_81139[10][10];
  wire [31:0] array_index_81141[10];
  wire [31:0] array_index_81142[10];
  wire [31:0] smul_81146;
  wire [31:0] add_81148;
  wire [31:0] array_update_81150[10];
  wire [31:0] add_81151;
  wire [31:0] array_update_81152[10][10];
  wire [31:0] array_index_81154[10];
  wire [31:0] array_index_81155[10];
  wire [31:0] smul_81159;
  wire [31:0] add_81161;
  wire [31:0] array_update_81163[10];
  wire [31:0] add_81164;
  wire [31:0] array_update_81165[10][10];
  wire [31:0] array_index_81167[10];
  wire [31:0] array_index_81168[10];
  wire [31:0] smul_81172;
  wire [31:0] add_81174;
  wire [31:0] array_update_81176[10];
  wire [31:0] add_81177;
  wire [31:0] array_update_81178[10][10];
  wire [31:0] array_index_81180[10];
  wire [31:0] array_index_81181[10];
  wire [31:0] smul_81185;
  wire [31:0] add_81187;
  wire [31:0] array_update_81189[10];
  wire [31:0] add_81190;
  wire [31:0] array_update_81191[10][10];
  wire [31:0] array_index_81193[10];
  wire [31:0] array_index_81194[10];
  wire [31:0] smul_81198;
  wire [31:0] add_81200;
  wire [31:0] array_update_81201[10];
  wire [31:0] array_update_81202[10][10];
  wire [31:0] array_index_81204[10];
  wire [31:0] add_81206;
  wire [31:0] array_update_81207[10];
  wire [31:0] literal_81208;
  wire [31:0] array_update_81209[10][10];
  wire [31:0] array_index_81211[10];
  wire [31:0] array_index_81212[10];
  wire [31:0] smul_81216;
  wire [31:0] add_81218;
  wire [31:0] array_update_81220[10];
  wire [31:0] add_81221;
  wire [31:0] array_update_81222[10][10];
  wire [31:0] array_index_81224[10];
  wire [31:0] array_index_81225[10];
  wire [31:0] smul_81229;
  wire [31:0] add_81231;
  wire [31:0] array_update_81233[10];
  wire [31:0] add_81234;
  wire [31:0] array_update_81235[10][10];
  wire [31:0] array_index_81237[10];
  wire [31:0] array_index_81238[10];
  wire [31:0] smul_81242;
  wire [31:0] add_81244;
  wire [31:0] array_update_81246[10];
  wire [31:0] add_81247;
  wire [31:0] array_update_81248[10][10];
  wire [31:0] array_index_81250[10];
  wire [31:0] array_index_81251[10];
  wire [31:0] smul_81255;
  wire [31:0] add_81257;
  wire [31:0] array_update_81259[10];
  wire [31:0] add_81260;
  wire [31:0] array_update_81261[10][10];
  wire [31:0] array_index_81263[10];
  wire [31:0] array_index_81264[10];
  wire [31:0] smul_81268;
  wire [31:0] add_81270;
  wire [31:0] array_update_81272[10];
  wire [31:0] add_81273;
  wire [31:0] array_update_81274[10][10];
  wire [31:0] array_index_81276[10];
  wire [31:0] array_index_81277[10];
  wire [31:0] smul_81281;
  wire [31:0] add_81283;
  wire [31:0] array_update_81285[10];
  wire [31:0] add_81286;
  wire [31:0] array_update_81287[10][10];
  wire [31:0] array_index_81289[10];
  wire [31:0] array_index_81290[10];
  wire [31:0] smul_81294;
  wire [31:0] add_81296;
  wire [31:0] array_update_81298[10];
  wire [31:0] add_81299;
  wire [31:0] array_update_81300[10][10];
  wire [31:0] array_index_81302[10];
  wire [31:0] array_index_81303[10];
  wire [31:0] smul_81307;
  wire [31:0] add_81309;
  wire [31:0] array_update_81311[10];
  wire [31:0] add_81312;
  wire [31:0] array_update_81313[10][10];
  wire [31:0] array_index_81315[10];
  wire [31:0] array_index_81316[10];
  wire [31:0] smul_81320;
  wire [31:0] add_81322;
  wire [31:0] array_update_81324[10];
  wire [31:0] add_81325;
  wire [31:0] array_update_81326[10][10];
  wire [31:0] array_index_81328[10];
  wire [31:0] array_index_81329[10];
  wire [31:0] smul_81333;
  wire [31:0] add_81335;
  wire [31:0] array_update_81336[10];
  wire [31:0] array_update_81337[10][10];
  wire [31:0] array_index_81339[10];
  wire [31:0] add_81341;
  wire [31:0] array_update_81342[10];
  wire [31:0] literal_81343;
  wire [31:0] array_update_81344[10][10];
  wire [31:0] array_index_81346[10];
  wire [31:0] array_index_81347[10];
  wire [31:0] smul_81351;
  wire [31:0] add_81353;
  wire [31:0] array_update_81355[10];
  wire [31:0] add_81356;
  wire [31:0] array_update_81357[10][10];
  wire [31:0] array_index_81359[10];
  wire [31:0] array_index_81360[10];
  wire [31:0] smul_81364;
  wire [31:0] add_81366;
  wire [31:0] array_update_81368[10];
  wire [31:0] add_81369;
  wire [31:0] array_update_81370[10][10];
  wire [31:0] array_index_81372[10];
  wire [31:0] array_index_81373[10];
  wire [31:0] smul_81377;
  wire [31:0] add_81379;
  wire [31:0] array_update_81381[10];
  wire [31:0] add_81382;
  wire [31:0] array_update_81383[10][10];
  wire [31:0] array_index_81385[10];
  wire [31:0] array_index_81386[10];
  wire [31:0] smul_81390;
  wire [31:0] add_81392;
  wire [31:0] array_update_81394[10];
  wire [31:0] add_81395;
  wire [31:0] array_update_81396[10][10];
  wire [31:0] array_index_81398[10];
  wire [31:0] array_index_81399[10];
  wire [31:0] smul_81403;
  wire [31:0] add_81405;
  wire [31:0] array_update_81407[10];
  wire [31:0] add_81408;
  wire [31:0] array_update_81409[10][10];
  wire [31:0] array_index_81411[10];
  wire [31:0] array_index_81412[10];
  wire [31:0] smul_81416;
  wire [31:0] add_81418;
  wire [31:0] array_update_81420[10];
  wire [31:0] add_81421;
  wire [31:0] array_update_81422[10][10];
  wire [31:0] array_index_81424[10];
  wire [31:0] array_index_81425[10];
  wire [31:0] smul_81429;
  wire [31:0] add_81431;
  wire [31:0] array_update_81433[10];
  wire [31:0] add_81434;
  wire [31:0] array_update_81435[10][10];
  wire [31:0] array_index_81437[10];
  wire [31:0] array_index_81438[10];
  wire [31:0] smul_81442;
  wire [31:0] add_81444;
  wire [31:0] array_update_81446[10];
  wire [31:0] add_81447;
  wire [31:0] array_update_81448[10][10];
  wire [31:0] array_index_81450[10];
  wire [31:0] array_index_81451[10];
  wire [31:0] smul_81455;
  wire [31:0] add_81457;
  wire [31:0] array_update_81459[10];
  wire [31:0] add_81460;
  wire [31:0] array_update_81461[10][10];
  wire [31:0] array_index_81463[10];
  wire [31:0] array_index_81464[10];
  wire [31:0] smul_81468;
  wire [31:0] add_81470;
  wire [31:0] array_update_81471[10];
  wire [31:0] array_update_81473[10][10];
  wire [31:0] add_81474;
  wire [31:0] array_index_81475[10];
  wire [31:0] literal_81477;
  wire [31:0] array_update_81478[10];
  wire [31:0] literal_81479;
  wire [31:0] array_update_81480[10][10];
  wire [31:0] array_index_81481[10];
  wire [31:0] array_index_81482[10];
  wire [31:0] array_index_81483[10];
  wire [31:0] smul_81487;
  wire [31:0] add_81489;
  wire [31:0] array_update_81491[10];
  wire [31:0] add_81492;
  wire [31:0] array_update_81493[10][10];
  wire [31:0] array_index_81495[10];
  wire [31:0] array_index_81496[10];
  wire [31:0] smul_81500;
  wire [31:0] add_81502;
  wire [31:0] array_update_81504[10];
  wire [31:0] add_81505;
  wire [31:0] array_update_81506[10][10];
  wire [31:0] array_index_81508[10];
  wire [31:0] array_index_81509[10];
  wire [31:0] smul_81513;
  wire [31:0] add_81515;
  wire [31:0] array_update_81517[10];
  wire [31:0] add_81518;
  wire [31:0] array_update_81519[10][10];
  wire [31:0] array_index_81521[10];
  wire [31:0] array_index_81522[10];
  wire [31:0] smul_81526;
  wire [31:0] add_81528;
  wire [31:0] array_update_81530[10];
  wire [31:0] add_81531;
  wire [31:0] array_update_81532[10][10];
  wire [31:0] array_index_81534[10];
  wire [31:0] array_index_81535[10];
  wire [31:0] smul_81539;
  wire [31:0] add_81541;
  wire [31:0] array_update_81543[10];
  wire [31:0] add_81544;
  wire [31:0] array_update_81545[10][10];
  wire [31:0] array_index_81547[10];
  wire [31:0] array_index_81548[10];
  wire [31:0] smul_81552;
  wire [31:0] add_81554;
  wire [31:0] array_update_81556[10];
  wire [31:0] add_81557;
  wire [31:0] array_update_81558[10][10];
  wire [31:0] array_index_81560[10];
  wire [31:0] array_index_81561[10];
  wire [31:0] smul_81565;
  wire [31:0] add_81567;
  wire [31:0] array_update_81569[10];
  wire [31:0] add_81570;
  wire [31:0] array_update_81571[10][10];
  wire [31:0] array_index_81573[10];
  wire [31:0] array_index_81574[10];
  wire [31:0] smul_81578;
  wire [31:0] add_81580;
  wire [31:0] array_update_81582[10];
  wire [31:0] add_81583;
  wire [31:0] array_update_81584[10][10];
  wire [31:0] array_index_81586[10];
  wire [31:0] array_index_81587[10];
  wire [31:0] smul_81591;
  wire [31:0] add_81593;
  wire [31:0] array_update_81595[10];
  wire [31:0] add_81596;
  wire [31:0] array_update_81597[10][10];
  wire [31:0] array_index_81599[10];
  wire [31:0] array_index_81600[10];
  wire [31:0] smul_81604;
  wire [31:0] add_81606;
  wire [31:0] array_update_81607[10];
  wire [31:0] array_update_81608[10][10];
  wire [31:0] array_index_81610[10];
  wire [31:0] add_81612;
  wire [31:0] array_update_81613[10];
  wire [31:0] literal_81614;
  wire [31:0] array_update_81615[10][10];
  wire [31:0] array_index_81617[10];
  wire [31:0] array_index_81618[10];
  wire [31:0] smul_81622;
  wire [31:0] add_81624;
  wire [31:0] array_update_81626[10];
  wire [31:0] add_81627;
  wire [31:0] array_update_81628[10][10];
  wire [31:0] array_index_81630[10];
  wire [31:0] array_index_81631[10];
  wire [31:0] smul_81635;
  wire [31:0] add_81637;
  wire [31:0] array_update_81639[10];
  wire [31:0] add_81640;
  wire [31:0] array_update_81641[10][10];
  wire [31:0] array_index_81643[10];
  wire [31:0] array_index_81644[10];
  wire [31:0] smul_81648;
  wire [31:0] add_81650;
  wire [31:0] array_update_81652[10];
  wire [31:0] add_81653;
  wire [31:0] array_update_81654[10][10];
  wire [31:0] array_index_81656[10];
  wire [31:0] array_index_81657[10];
  wire [31:0] smul_81661;
  wire [31:0] add_81663;
  wire [31:0] array_update_81665[10];
  wire [31:0] add_81666;
  wire [31:0] array_update_81667[10][10];
  wire [31:0] array_index_81669[10];
  wire [31:0] array_index_81670[10];
  wire [31:0] smul_81674;
  wire [31:0] add_81676;
  wire [31:0] array_update_81678[10];
  wire [31:0] add_81679;
  wire [31:0] array_update_81680[10][10];
  wire [31:0] array_index_81682[10];
  wire [31:0] array_index_81683[10];
  wire [31:0] smul_81687;
  wire [31:0] add_81689;
  wire [31:0] array_update_81691[10];
  wire [31:0] add_81692;
  wire [31:0] array_update_81693[10][10];
  wire [31:0] array_index_81695[10];
  wire [31:0] array_index_81696[10];
  wire [31:0] smul_81700;
  wire [31:0] add_81702;
  wire [31:0] array_update_81704[10];
  wire [31:0] add_81705;
  wire [31:0] array_update_81706[10][10];
  wire [31:0] array_index_81708[10];
  wire [31:0] array_index_81709[10];
  wire [31:0] smul_81713;
  wire [31:0] add_81715;
  wire [31:0] array_update_81717[10];
  wire [31:0] add_81718;
  wire [31:0] array_update_81719[10][10];
  wire [31:0] array_index_81721[10];
  wire [31:0] array_index_81722[10];
  wire [31:0] smul_81726;
  wire [31:0] add_81728;
  wire [31:0] array_update_81730[10];
  wire [31:0] add_81731;
  wire [31:0] array_update_81732[10][10];
  wire [31:0] array_index_81734[10];
  wire [31:0] array_index_81735[10];
  wire [31:0] smul_81739;
  wire [31:0] add_81741;
  wire [31:0] array_update_81742[10];
  wire [31:0] array_update_81743[10][10];
  wire [31:0] array_index_81745[10];
  wire [31:0] add_81747;
  wire [31:0] array_update_81748[10];
  wire [31:0] literal_81749;
  wire [31:0] array_update_81750[10][10];
  wire [31:0] array_index_81752[10];
  wire [31:0] array_index_81753[10];
  wire [31:0] smul_81757;
  wire [31:0] add_81759;
  wire [31:0] array_update_81761[10];
  wire [31:0] add_81762;
  wire [31:0] array_update_81763[10][10];
  wire [31:0] array_index_81765[10];
  wire [31:0] array_index_81766[10];
  wire [31:0] smul_81770;
  wire [31:0] add_81772;
  wire [31:0] array_update_81774[10];
  wire [31:0] add_81775;
  wire [31:0] array_update_81776[10][10];
  wire [31:0] array_index_81778[10];
  wire [31:0] array_index_81779[10];
  wire [31:0] smul_81783;
  wire [31:0] add_81785;
  wire [31:0] array_update_81787[10];
  wire [31:0] add_81788;
  wire [31:0] array_update_81789[10][10];
  wire [31:0] array_index_81791[10];
  wire [31:0] array_index_81792[10];
  wire [31:0] smul_81796;
  wire [31:0] add_81798;
  wire [31:0] array_update_81800[10];
  wire [31:0] add_81801;
  wire [31:0] array_update_81802[10][10];
  wire [31:0] array_index_81804[10];
  wire [31:0] array_index_81805[10];
  wire [31:0] smul_81809;
  wire [31:0] add_81811;
  wire [31:0] array_update_81813[10];
  wire [31:0] add_81814;
  wire [31:0] array_update_81815[10][10];
  wire [31:0] array_index_81817[10];
  wire [31:0] array_index_81818[10];
  wire [31:0] smul_81822;
  wire [31:0] add_81824;
  wire [31:0] array_update_81826[10];
  wire [31:0] add_81827;
  wire [31:0] array_update_81828[10][10];
  wire [31:0] array_index_81830[10];
  wire [31:0] array_index_81831[10];
  wire [31:0] smul_81835;
  wire [31:0] add_81837;
  wire [31:0] array_update_81839[10];
  wire [31:0] add_81840;
  wire [31:0] array_update_81841[10][10];
  wire [31:0] array_index_81843[10];
  wire [31:0] array_index_81844[10];
  wire [31:0] smul_81848;
  wire [31:0] add_81850;
  wire [31:0] array_update_81852[10];
  wire [31:0] add_81853;
  wire [31:0] array_update_81854[10][10];
  wire [31:0] array_index_81856[10];
  wire [31:0] array_index_81857[10];
  wire [31:0] smul_81861;
  wire [31:0] add_81863;
  wire [31:0] array_update_81865[10];
  wire [31:0] add_81866;
  wire [31:0] array_update_81867[10][10];
  wire [31:0] array_index_81869[10];
  wire [31:0] array_index_81870[10];
  wire [31:0] smul_81874;
  wire [31:0] add_81876;
  wire [31:0] array_update_81877[10];
  wire [31:0] array_update_81878[10][10];
  wire [31:0] array_index_81880[10];
  wire [31:0] add_81882;
  wire [31:0] array_update_81883[10];
  wire [31:0] literal_81884;
  wire [31:0] array_update_81885[10][10];
  wire [31:0] array_index_81887[10];
  wire [31:0] array_index_81888[10];
  wire [31:0] smul_81892;
  wire [31:0] add_81894;
  wire [31:0] array_update_81896[10];
  wire [31:0] add_81897;
  wire [31:0] array_update_81898[10][10];
  wire [31:0] array_index_81900[10];
  wire [31:0] array_index_81901[10];
  wire [31:0] smul_81905;
  wire [31:0] add_81907;
  wire [31:0] array_update_81909[10];
  wire [31:0] add_81910;
  wire [31:0] array_update_81911[10][10];
  wire [31:0] array_index_81913[10];
  wire [31:0] array_index_81914[10];
  wire [31:0] smul_81918;
  wire [31:0] add_81920;
  wire [31:0] array_update_81922[10];
  wire [31:0] add_81923;
  wire [31:0] array_update_81924[10][10];
  wire [31:0] array_index_81926[10];
  wire [31:0] array_index_81927[10];
  wire [31:0] smul_81931;
  wire [31:0] add_81933;
  wire [31:0] array_update_81935[10];
  wire [31:0] add_81936;
  wire [31:0] array_update_81937[10][10];
  wire [31:0] array_index_81939[10];
  wire [31:0] array_index_81940[10];
  wire [31:0] smul_81944;
  wire [31:0] add_81946;
  wire [31:0] array_update_81948[10];
  wire [31:0] add_81949;
  wire [31:0] array_update_81950[10][10];
  wire [31:0] array_index_81952[10];
  wire [31:0] array_index_81953[10];
  wire [31:0] smul_81957;
  wire [31:0] add_81959;
  wire [31:0] array_update_81961[10];
  wire [31:0] add_81962;
  wire [31:0] array_update_81963[10][10];
  wire [31:0] array_index_81965[10];
  wire [31:0] array_index_81966[10];
  wire [31:0] smul_81970;
  wire [31:0] add_81972;
  wire [31:0] array_update_81974[10];
  wire [31:0] add_81975;
  wire [31:0] array_update_81976[10][10];
  wire [31:0] array_index_81978[10];
  wire [31:0] array_index_81979[10];
  wire [31:0] smul_81983;
  wire [31:0] add_81985;
  wire [31:0] array_update_81987[10];
  wire [31:0] add_81988;
  wire [31:0] array_update_81989[10][10];
  wire [31:0] array_index_81991[10];
  wire [31:0] array_index_81992[10];
  wire [31:0] smul_81996;
  wire [31:0] add_81998;
  wire [31:0] array_update_82000[10];
  wire [31:0] add_82001;
  wire [31:0] array_update_82002[10][10];
  wire [31:0] array_index_82004[10];
  wire [31:0] array_index_82005[10];
  wire [31:0] smul_82009;
  wire [31:0] add_82011;
  wire [31:0] array_update_82012[10];
  wire [31:0] array_update_82013[10][10];
  wire [31:0] array_index_82015[10];
  wire [31:0] add_82017;
  wire [31:0] array_update_82018[10];
  wire [31:0] literal_82019;
  wire [31:0] array_update_82020[10][10];
  wire [31:0] array_index_82022[10];
  wire [31:0] array_index_82023[10];
  wire [31:0] smul_82027;
  wire [31:0] add_82029;
  wire [31:0] array_update_82031[10];
  wire [31:0] add_82032;
  wire [31:0] array_update_82033[10][10];
  wire [31:0] array_index_82035[10];
  wire [31:0] array_index_82036[10];
  wire [31:0] smul_82040;
  wire [31:0] add_82042;
  wire [31:0] array_update_82044[10];
  wire [31:0] add_82045;
  wire [31:0] array_update_82046[10][10];
  wire [31:0] array_index_82048[10];
  wire [31:0] array_index_82049[10];
  wire [31:0] smul_82053;
  wire [31:0] add_82055;
  wire [31:0] array_update_82057[10];
  wire [31:0] add_82058;
  wire [31:0] array_update_82059[10][10];
  wire [31:0] array_index_82061[10];
  wire [31:0] array_index_82062[10];
  wire [31:0] smul_82066;
  wire [31:0] add_82068;
  wire [31:0] array_update_82070[10];
  wire [31:0] add_82071;
  wire [31:0] array_update_82072[10][10];
  wire [31:0] array_index_82074[10];
  wire [31:0] array_index_82075[10];
  wire [31:0] smul_82079;
  wire [31:0] add_82081;
  wire [31:0] array_update_82083[10];
  wire [31:0] add_82084;
  wire [31:0] array_update_82085[10][10];
  wire [31:0] array_index_82087[10];
  wire [31:0] array_index_82088[10];
  wire [31:0] smul_82092;
  wire [31:0] add_82094;
  wire [31:0] array_update_82096[10];
  wire [31:0] add_82097;
  wire [31:0] array_update_82098[10][10];
  wire [31:0] array_index_82100[10];
  wire [31:0] array_index_82101[10];
  wire [31:0] smul_82105;
  wire [31:0] add_82107;
  wire [31:0] array_update_82109[10];
  wire [31:0] add_82110;
  wire [31:0] array_update_82111[10][10];
  wire [31:0] array_index_82113[10];
  wire [31:0] array_index_82114[10];
  wire [31:0] smul_82118;
  wire [31:0] add_82120;
  wire [31:0] array_update_82122[10];
  wire [31:0] add_82123;
  wire [31:0] array_update_82124[10][10];
  wire [31:0] array_index_82126[10];
  wire [31:0] array_index_82127[10];
  wire [31:0] smul_82131;
  wire [31:0] add_82133;
  wire [31:0] array_update_82135[10];
  wire [31:0] add_82136;
  wire [31:0] array_update_82137[10][10];
  wire [31:0] array_index_82139[10];
  wire [31:0] array_index_82140[10];
  wire [31:0] smul_82144;
  wire [31:0] add_82146;
  wire [31:0] array_update_82147[10];
  wire [31:0] array_update_82148[10][10];
  wire [31:0] array_index_82150[10];
  wire [31:0] add_82152;
  wire [31:0] array_update_82153[10];
  wire [31:0] literal_82154;
  wire [31:0] array_update_82155[10][10];
  wire [31:0] array_index_82157[10];
  wire [31:0] array_index_82158[10];
  wire [31:0] smul_82162;
  wire [31:0] add_82164;
  wire [31:0] array_update_82166[10];
  wire [31:0] add_82167;
  wire [31:0] array_update_82168[10][10];
  wire [31:0] array_index_82170[10];
  wire [31:0] array_index_82171[10];
  wire [31:0] smul_82175;
  wire [31:0] add_82177;
  wire [31:0] array_update_82179[10];
  wire [31:0] add_82180;
  wire [31:0] array_update_82181[10][10];
  wire [31:0] array_index_82183[10];
  wire [31:0] array_index_82184[10];
  wire [31:0] smul_82188;
  wire [31:0] add_82190;
  wire [31:0] array_update_82192[10];
  wire [31:0] add_82193;
  wire [31:0] array_update_82194[10][10];
  wire [31:0] array_index_82196[10];
  wire [31:0] array_index_82197[10];
  wire [31:0] smul_82201;
  wire [31:0] add_82203;
  wire [31:0] array_update_82205[10];
  wire [31:0] add_82206;
  wire [31:0] array_update_82207[10][10];
  wire [31:0] array_index_82209[10];
  wire [31:0] array_index_82210[10];
  wire [31:0] smul_82214;
  wire [31:0] add_82216;
  wire [31:0] array_update_82218[10];
  wire [31:0] add_82219;
  wire [31:0] array_update_82220[10][10];
  wire [31:0] array_index_82222[10];
  wire [31:0] array_index_82223[10];
  wire [31:0] smul_82227;
  wire [31:0] add_82229;
  wire [31:0] array_update_82231[10];
  wire [31:0] add_82232;
  wire [31:0] array_update_82233[10][10];
  wire [31:0] array_index_82235[10];
  wire [31:0] array_index_82236[10];
  wire [31:0] smul_82240;
  wire [31:0] add_82242;
  wire [31:0] array_update_82244[10];
  wire [31:0] add_82245;
  wire [31:0] array_update_82246[10][10];
  wire [31:0] array_index_82248[10];
  wire [31:0] array_index_82249[10];
  wire [31:0] smul_82253;
  wire [31:0] add_82255;
  wire [31:0] array_update_82257[10];
  wire [31:0] add_82258;
  wire [31:0] array_update_82259[10][10];
  wire [31:0] array_index_82261[10];
  wire [31:0] array_index_82262[10];
  wire [31:0] smul_82266;
  wire [31:0] add_82268;
  wire [31:0] array_update_82270[10];
  wire [31:0] add_82271;
  wire [31:0] array_update_82272[10][10];
  wire [31:0] array_index_82274[10];
  wire [31:0] array_index_82275[10];
  wire [31:0] smul_82279;
  wire [31:0] add_82281;
  wire [31:0] array_update_82282[10];
  wire [31:0] array_update_82283[10][10];
  wire [31:0] array_index_82285[10];
  wire [31:0] add_82287;
  wire [31:0] array_update_82288[10];
  wire [31:0] literal_82289;
  wire [31:0] array_update_82290[10][10];
  wire [31:0] array_index_82292[10];
  wire [31:0] array_index_82293[10];
  wire [31:0] smul_82297;
  wire [31:0] add_82299;
  wire [31:0] array_update_82301[10];
  wire [31:0] add_82302;
  wire [31:0] array_update_82303[10][10];
  wire [31:0] array_index_82305[10];
  wire [31:0] array_index_82306[10];
  wire [31:0] smul_82310;
  wire [31:0] add_82312;
  wire [31:0] array_update_82314[10];
  wire [31:0] add_82315;
  wire [31:0] array_update_82316[10][10];
  wire [31:0] array_index_82318[10];
  wire [31:0] array_index_82319[10];
  wire [31:0] smul_82323;
  wire [31:0] add_82325;
  wire [31:0] array_update_82327[10];
  wire [31:0] add_82328;
  wire [31:0] array_update_82329[10][10];
  wire [31:0] array_index_82331[10];
  wire [31:0] array_index_82332[10];
  wire [31:0] smul_82336;
  wire [31:0] add_82338;
  wire [31:0] array_update_82340[10];
  wire [31:0] add_82341;
  wire [31:0] array_update_82342[10][10];
  wire [31:0] array_index_82344[10];
  wire [31:0] array_index_82345[10];
  wire [31:0] smul_82349;
  wire [31:0] add_82351;
  wire [31:0] array_update_82353[10];
  wire [31:0] add_82354;
  wire [31:0] array_update_82355[10][10];
  wire [31:0] array_index_82357[10];
  wire [31:0] array_index_82358[10];
  wire [31:0] smul_82362;
  wire [31:0] add_82364;
  wire [31:0] array_update_82366[10];
  wire [31:0] add_82367;
  wire [31:0] array_update_82368[10][10];
  wire [31:0] array_index_82370[10];
  wire [31:0] array_index_82371[10];
  wire [31:0] smul_82375;
  wire [31:0] add_82377;
  wire [31:0] array_update_82379[10];
  wire [31:0] add_82380;
  wire [31:0] array_update_82381[10][10];
  wire [31:0] array_index_82383[10];
  wire [31:0] array_index_82384[10];
  wire [31:0] smul_82388;
  wire [31:0] add_82390;
  wire [31:0] array_update_82392[10];
  wire [31:0] add_82393;
  wire [31:0] array_update_82394[10][10];
  wire [31:0] array_index_82396[10];
  wire [31:0] array_index_82397[10];
  wire [31:0] smul_82401;
  wire [31:0] add_82403;
  wire [31:0] array_update_82405[10];
  wire [31:0] add_82406;
  wire [31:0] array_update_82407[10][10];
  wire [31:0] array_index_82409[10];
  wire [31:0] array_index_82410[10];
  wire [31:0] smul_82414;
  wire [31:0] add_82416;
  wire [31:0] array_update_82417[10];
  wire [31:0] array_update_82418[10][10];
  wire [31:0] array_index_82420[10];
  wire [31:0] add_82422;
  wire [31:0] array_update_82423[10];
  wire [31:0] literal_82424;
  wire [31:0] array_update_82425[10][10];
  wire [31:0] array_index_82427[10];
  wire [31:0] array_index_82428[10];
  wire [31:0] smul_82432;
  wire [31:0] add_82434;
  wire [31:0] array_update_82436[10];
  wire [31:0] add_82437;
  wire [31:0] array_update_82438[10][10];
  wire [31:0] array_index_82440[10];
  wire [31:0] array_index_82441[10];
  wire [31:0] smul_82445;
  wire [31:0] add_82447;
  wire [31:0] array_update_82449[10];
  wire [31:0] add_82450;
  wire [31:0] array_update_82451[10][10];
  wire [31:0] array_index_82453[10];
  wire [31:0] array_index_82454[10];
  wire [31:0] smul_82458;
  wire [31:0] add_82460;
  wire [31:0] array_update_82462[10];
  wire [31:0] add_82463;
  wire [31:0] array_update_82464[10][10];
  wire [31:0] array_index_82466[10];
  wire [31:0] array_index_82467[10];
  wire [31:0] smul_82471;
  wire [31:0] add_82473;
  wire [31:0] array_update_82475[10];
  wire [31:0] add_82476;
  wire [31:0] array_update_82477[10][10];
  wire [31:0] array_index_82479[10];
  wire [31:0] array_index_82480[10];
  wire [31:0] smul_82484;
  wire [31:0] add_82486;
  wire [31:0] array_update_82488[10];
  wire [31:0] add_82489;
  wire [31:0] array_update_82490[10][10];
  wire [31:0] array_index_82492[10];
  wire [31:0] array_index_82493[10];
  wire [31:0] smul_82497;
  wire [31:0] add_82499;
  wire [31:0] array_update_82501[10];
  wire [31:0] add_82502;
  wire [31:0] array_update_82503[10][10];
  wire [31:0] array_index_82505[10];
  wire [31:0] array_index_82506[10];
  wire [31:0] smul_82510;
  wire [31:0] add_82512;
  wire [31:0] array_update_82514[10];
  wire [31:0] add_82515;
  wire [31:0] array_update_82516[10][10];
  wire [31:0] array_index_82518[10];
  wire [31:0] array_index_82519[10];
  wire [31:0] smul_82523;
  wire [31:0] add_82525;
  wire [31:0] array_update_82527[10];
  wire [31:0] add_82528;
  wire [31:0] array_update_82529[10][10];
  wire [31:0] array_index_82531[10];
  wire [31:0] array_index_82532[10];
  wire [31:0] smul_82536;
  wire [31:0] add_82538;
  wire [31:0] array_update_82540[10];
  wire [31:0] add_82541;
  wire [31:0] array_update_82542[10][10];
  wire [31:0] array_index_82544[10];
  wire [31:0] array_index_82545[10];
  wire [31:0] smul_82549;
  wire [31:0] add_82551;
  wire [31:0] array_update_82552[10];
  wire [31:0] array_update_82553[10][10];
  wire [31:0] array_index_82555[10];
  wire [31:0] add_82557;
  wire [31:0] array_update_82558[10];
  wire [31:0] literal_82559;
  wire [31:0] array_update_82560[10][10];
  wire [31:0] array_index_82562[10];
  wire [31:0] array_index_82563[10];
  wire [31:0] smul_82567;
  wire [31:0] add_82569;
  wire [31:0] array_update_82571[10];
  wire [31:0] add_82572;
  wire [31:0] array_update_82573[10][10];
  wire [31:0] array_index_82575[10];
  wire [31:0] array_index_82576[10];
  wire [31:0] smul_82580;
  wire [31:0] add_82582;
  wire [31:0] array_update_82584[10];
  wire [31:0] add_82585;
  wire [31:0] array_update_82586[10][10];
  wire [31:0] array_index_82588[10];
  wire [31:0] array_index_82589[10];
  wire [31:0] smul_82593;
  wire [31:0] add_82595;
  wire [31:0] array_update_82597[10];
  wire [31:0] add_82598;
  wire [31:0] array_update_82599[10][10];
  wire [31:0] array_index_82601[10];
  wire [31:0] array_index_82602[10];
  wire [31:0] smul_82606;
  wire [31:0] add_82608;
  wire [31:0] array_update_82610[10];
  wire [31:0] add_82611;
  wire [31:0] array_update_82612[10][10];
  wire [31:0] array_index_82614[10];
  wire [31:0] array_index_82615[10];
  wire [31:0] smul_82619;
  wire [31:0] add_82621;
  wire [31:0] array_update_82623[10];
  wire [31:0] add_82624;
  wire [31:0] array_update_82625[10][10];
  wire [31:0] array_index_82627[10];
  wire [31:0] array_index_82628[10];
  wire [31:0] smul_82632;
  wire [31:0] add_82634;
  wire [31:0] array_update_82636[10];
  wire [31:0] add_82637;
  wire [31:0] array_update_82638[10][10];
  wire [31:0] array_index_82640[10];
  wire [31:0] array_index_82641[10];
  wire [31:0] smul_82645;
  wire [31:0] add_82647;
  wire [31:0] array_update_82649[10];
  wire [31:0] add_82650;
  wire [31:0] array_update_82651[10][10];
  wire [31:0] array_index_82653[10];
  wire [31:0] array_index_82654[10];
  wire [31:0] smul_82658;
  wire [31:0] add_82660;
  wire [31:0] array_update_82662[10];
  wire [31:0] add_82663;
  wire [31:0] array_update_82664[10][10];
  wire [31:0] array_index_82666[10];
  wire [31:0] array_index_82667[10];
  wire [31:0] smul_82671;
  wire [31:0] add_82673;
  wire [31:0] array_update_82675[10];
  wire [31:0] add_82676;
  wire [31:0] array_update_82677[10][10];
  wire [31:0] array_index_82679[10];
  wire [31:0] array_index_82680[10];
  wire [31:0] smul_82684;
  wire [31:0] add_82686;
  wire [31:0] array_update_82687[10];
  wire [31:0] array_update_82688[10][10];
  wire [31:0] array_index_82690[10];
  wire [31:0] add_82692;
  wire [31:0] array_update_82693[10];
  wire [31:0] literal_82694;
  wire [31:0] array_update_82695[10][10];
  wire [31:0] array_index_82697[10];
  wire [31:0] array_index_82698[10];
  wire [31:0] smul_82702;
  wire [31:0] add_82704;
  wire [31:0] array_update_82706[10];
  wire [31:0] add_82707;
  wire [31:0] array_update_82708[10][10];
  wire [31:0] array_index_82710[10];
  wire [31:0] array_index_82711[10];
  wire [31:0] smul_82715;
  wire [31:0] add_82717;
  wire [31:0] array_update_82719[10];
  wire [31:0] add_82720;
  wire [31:0] array_update_82721[10][10];
  wire [31:0] array_index_82723[10];
  wire [31:0] array_index_82724[10];
  wire [31:0] smul_82728;
  wire [31:0] add_82730;
  wire [31:0] array_update_82732[10];
  wire [31:0] add_82733;
  wire [31:0] array_update_82734[10][10];
  wire [31:0] array_index_82736[10];
  wire [31:0] array_index_82737[10];
  wire [31:0] smul_82741;
  wire [31:0] add_82743;
  wire [31:0] array_update_82745[10];
  wire [31:0] add_82746;
  wire [31:0] array_update_82747[10][10];
  wire [31:0] array_index_82749[10];
  wire [31:0] array_index_82750[10];
  wire [31:0] smul_82754;
  wire [31:0] add_82756;
  wire [31:0] array_update_82758[10];
  wire [31:0] add_82759;
  wire [31:0] array_update_82760[10][10];
  wire [31:0] array_index_82762[10];
  wire [31:0] array_index_82763[10];
  wire [31:0] smul_82767;
  wire [31:0] add_82769;
  wire [31:0] array_update_82771[10];
  wire [31:0] add_82772;
  wire [31:0] array_update_82773[10][10];
  wire [31:0] array_index_82775[10];
  wire [31:0] array_index_82776[10];
  wire [31:0] smul_82780;
  wire [31:0] add_82782;
  wire [31:0] array_update_82784[10];
  wire [31:0] add_82785;
  wire [31:0] array_update_82786[10][10];
  wire [31:0] array_index_82788[10];
  wire [31:0] array_index_82789[10];
  wire [31:0] smul_82793;
  wire [31:0] add_82795;
  wire [31:0] array_update_82797[10];
  wire [31:0] add_82798;
  wire [31:0] array_update_82799[10][10];
  wire [31:0] array_index_82801[10];
  wire [31:0] array_index_82802[10];
  wire [31:0] smul_82806;
  wire [31:0] add_82808;
  wire [31:0] array_update_82810[10];
  wire [31:0] add_82811;
  wire [31:0] array_update_82812[10][10];
  wire [31:0] array_index_82814[10];
  wire [31:0] array_index_82815[10];
  wire [31:0] smul_82819;
  wire [31:0] add_82821;
  wire [31:0] array_update_82822[10];
  wire [31:0] array_update_82824[10][10];
  wire [31:0] add_82825;
  wire [31:0] array_index_82826[10];
  wire [31:0] literal_82828;
  wire [31:0] array_update_82829[10];
  wire [31:0] literal_82830;
  wire [31:0] array_update_82831[10][10];
  wire [31:0] array_index_82832[10];
  wire [31:0] array_index_82833[10];
  wire [31:0] array_index_82834[10];
  wire [31:0] smul_82838;
  wire [31:0] add_82840;
  wire [31:0] array_update_82842[10];
  wire [31:0] add_82843;
  wire [31:0] array_update_82844[10][10];
  wire [31:0] array_index_82846[10];
  wire [31:0] array_index_82847[10];
  wire [31:0] smul_82851;
  wire [31:0] add_82853;
  wire [31:0] array_update_82855[10];
  wire [31:0] add_82856;
  wire [31:0] array_update_82857[10][10];
  wire [31:0] array_index_82859[10];
  wire [31:0] array_index_82860[10];
  wire [31:0] smul_82864;
  wire [31:0] add_82866;
  wire [31:0] array_update_82868[10];
  wire [31:0] add_82869;
  wire [31:0] array_update_82870[10][10];
  wire [31:0] array_index_82872[10];
  wire [31:0] array_index_82873[10];
  wire [31:0] smul_82877;
  wire [31:0] add_82879;
  wire [31:0] array_update_82881[10];
  wire [31:0] add_82882;
  wire [31:0] array_update_82883[10][10];
  wire [31:0] array_index_82885[10];
  wire [31:0] array_index_82886[10];
  wire [31:0] smul_82890;
  wire [31:0] add_82892;
  wire [31:0] array_update_82894[10];
  wire [31:0] add_82895;
  wire [31:0] array_update_82896[10][10];
  wire [31:0] array_index_82898[10];
  wire [31:0] array_index_82899[10];
  wire [31:0] smul_82903;
  wire [31:0] add_82905;
  wire [31:0] array_update_82907[10];
  wire [31:0] add_82908;
  wire [31:0] array_update_82909[10][10];
  wire [31:0] array_index_82911[10];
  wire [31:0] array_index_82912[10];
  wire [31:0] smul_82916;
  wire [31:0] add_82918;
  wire [31:0] array_update_82920[10];
  wire [31:0] add_82921;
  wire [31:0] array_update_82922[10][10];
  wire [31:0] array_index_82924[10];
  wire [31:0] array_index_82925[10];
  wire [31:0] smul_82929;
  wire [31:0] add_82931;
  wire [31:0] array_update_82933[10];
  wire [31:0] add_82934;
  wire [31:0] array_update_82935[10][10];
  wire [31:0] array_index_82937[10];
  wire [31:0] array_index_82938[10];
  wire [31:0] smul_82942;
  wire [31:0] add_82944;
  wire [31:0] array_update_82946[10];
  wire [31:0] add_82947;
  wire [31:0] array_update_82948[10][10];
  wire [31:0] array_index_82950[10];
  wire [31:0] array_index_82951[10];
  wire [31:0] smul_82955;
  wire [31:0] add_82957;
  wire [31:0] array_update_82958[10];
  wire [31:0] array_update_82959[10][10];
  wire [31:0] array_index_82961[10];
  wire [31:0] add_82963;
  wire [31:0] array_update_82964[10];
  wire [31:0] literal_82965;
  wire [31:0] array_update_82966[10][10];
  wire [31:0] array_index_82968[10];
  wire [31:0] array_index_82969[10];
  wire [31:0] smul_82973;
  wire [31:0] add_82975;
  wire [31:0] array_update_82977[10];
  wire [31:0] add_82978;
  wire [31:0] array_update_82979[10][10];
  wire [31:0] array_index_82981[10];
  wire [31:0] array_index_82982[10];
  wire [31:0] smul_82986;
  wire [31:0] add_82988;
  wire [31:0] array_update_82990[10];
  wire [31:0] add_82991;
  wire [31:0] array_update_82992[10][10];
  wire [31:0] array_index_82994[10];
  wire [31:0] array_index_82995[10];
  wire [31:0] smul_82999;
  wire [31:0] add_83001;
  wire [31:0] array_update_83003[10];
  wire [31:0] add_83004;
  wire [31:0] array_update_83005[10][10];
  wire [31:0] array_index_83007[10];
  wire [31:0] array_index_83008[10];
  wire [31:0] smul_83012;
  wire [31:0] add_83014;
  wire [31:0] array_update_83016[10];
  wire [31:0] add_83017;
  wire [31:0] array_update_83018[10][10];
  wire [31:0] array_index_83020[10];
  wire [31:0] array_index_83021[10];
  wire [31:0] smul_83025;
  wire [31:0] add_83027;
  wire [31:0] array_update_83029[10];
  wire [31:0] add_83030;
  wire [31:0] array_update_83031[10][10];
  wire [31:0] array_index_83033[10];
  wire [31:0] array_index_83034[10];
  wire [31:0] smul_83038;
  wire [31:0] add_83040;
  wire [31:0] array_update_83042[10];
  wire [31:0] add_83043;
  wire [31:0] array_update_83044[10][10];
  wire [31:0] array_index_83046[10];
  wire [31:0] array_index_83047[10];
  wire [31:0] smul_83051;
  wire [31:0] add_83053;
  wire [31:0] array_update_83055[10];
  wire [31:0] add_83056;
  wire [31:0] array_update_83057[10][10];
  wire [31:0] array_index_83059[10];
  wire [31:0] array_index_83060[10];
  wire [31:0] smul_83064;
  wire [31:0] add_83066;
  wire [31:0] array_update_83068[10];
  wire [31:0] add_83069;
  wire [31:0] array_update_83070[10][10];
  wire [31:0] array_index_83072[10];
  wire [31:0] array_index_83073[10];
  wire [31:0] smul_83077;
  wire [31:0] add_83079;
  wire [31:0] array_update_83081[10];
  wire [31:0] add_83082;
  wire [31:0] array_update_83083[10][10];
  wire [31:0] array_index_83085[10];
  wire [31:0] array_index_83086[10];
  wire [31:0] smul_83090;
  wire [31:0] add_83092;
  wire [31:0] array_update_83093[10];
  wire [31:0] array_update_83094[10][10];
  wire [31:0] array_index_83096[10];
  wire [31:0] add_83098;
  wire [31:0] array_update_83099[10];
  wire [31:0] literal_83100;
  wire [31:0] array_update_83101[10][10];
  wire [31:0] array_index_83103[10];
  wire [31:0] array_index_83104[10];
  wire [31:0] smul_83108;
  wire [31:0] add_83110;
  wire [31:0] array_update_83112[10];
  wire [31:0] add_83113;
  wire [31:0] array_update_83114[10][10];
  wire [31:0] array_index_83116[10];
  wire [31:0] array_index_83117[10];
  wire [31:0] smul_83121;
  wire [31:0] add_83123;
  wire [31:0] array_update_83125[10];
  wire [31:0] add_83126;
  wire [31:0] array_update_83127[10][10];
  wire [31:0] array_index_83129[10];
  wire [31:0] array_index_83130[10];
  wire [31:0] smul_83134;
  wire [31:0] add_83136;
  wire [31:0] array_update_83138[10];
  wire [31:0] add_83139;
  wire [31:0] array_update_83140[10][10];
  wire [31:0] array_index_83142[10];
  wire [31:0] array_index_83143[10];
  wire [31:0] smul_83147;
  wire [31:0] add_83149;
  wire [31:0] array_update_83151[10];
  wire [31:0] add_83152;
  wire [31:0] array_update_83153[10][10];
  wire [31:0] array_index_83155[10];
  wire [31:0] array_index_83156[10];
  wire [31:0] smul_83160;
  wire [31:0] add_83162;
  wire [31:0] array_update_83164[10];
  wire [31:0] add_83165;
  wire [31:0] array_update_83166[10][10];
  wire [31:0] array_index_83168[10];
  wire [31:0] array_index_83169[10];
  wire [31:0] smul_83173;
  wire [31:0] add_83175;
  wire [31:0] array_update_83177[10];
  wire [31:0] add_83178;
  wire [31:0] array_update_83179[10][10];
  wire [31:0] array_index_83181[10];
  wire [31:0] array_index_83182[10];
  wire [31:0] smul_83186;
  wire [31:0] add_83188;
  wire [31:0] array_update_83190[10];
  wire [31:0] add_83191;
  wire [31:0] array_update_83192[10][10];
  wire [31:0] array_index_83194[10];
  wire [31:0] array_index_83195[10];
  wire [31:0] smul_83199;
  wire [31:0] add_83201;
  wire [31:0] array_update_83203[10];
  wire [31:0] add_83204;
  wire [31:0] array_update_83205[10][10];
  wire [31:0] array_index_83207[10];
  wire [31:0] array_index_83208[10];
  wire [31:0] smul_83212;
  wire [31:0] add_83214;
  wire [31:0] array_update_83216[10];
  wire [31:0] add_83217;
  wire [31:0] array_update_83218[10][10];
  wire [31:0] array_index_83220[10];
  wire [31:0] array_index_83221[10];
  wire [31:0] smul_83225;
  wire [31:0] add_83227;
  wire [31:0] array_update_83228[10];
  wire [31:0] array_update_83229[10][10];
  wire [31:0] array_index_83231[10];
  wire [31:0] add_83233;
  wire [31:0] array_update_83234[10];
  wire [31:0] literal_83235;
  wire [31:0] array_update_83236[10][10];
  wire [31:0] array_index_83238[10];
  wire [31:0] array_index_83239[10];
  wire [31:0] smul_83243;
  wire [31:0] add_83245;
  wire [31:0] array_update_83247[10];
  wire [31:0] add_83248;
  wire [31:0] array_update_83249[10][10];
  wire [31:0] array_index_83251[10];
  wire [31:0] array_index_83252[10];
  wire [31:0] smul_83256;
  wire [31:0] add_83258;
  wire [31:0] array_update_83260[10];
  wire [31:0] add_83261;
  wire [31:0] array_update_83262[10][10];
  wire [31:0] array_index_83264[10];
  wire [31:0] array_index_83265[10];
  wire [31:0] smul_83269;
  wire [31:0] add_83271;
  wire [31:0] array_update_83273[10];
  wire [31:0] add_83274;
  wire [31:0] array_update_83275[10][10];
  wire [31:0] array_index_83277[10];
  wire [31:0] array_index_83278[10];
  wire [31:0] smul_83282;
  wire [31:0] add_83284;
  wire [31:0] array_update_83286[10];
  wire [31:0] add_83287;
  wire [31:0] array_update_83288[10][10];
  wire [31:0] array_index_83290[10];
  wire [31:0] array_index_83291[10];
  wire [31:0] smul_83295;
  wire [31:0] add_83297;
  wire [31:0] array_update_83299[10];
  wire [31:0] add_83300;
  wire [31:0] array_update_83301[10][10];
  wire [31:0] array_index_83303[10];
  wire [31:0] array_index_83304[10];
  wire [31:0] smul_83308;
  wire [31:0] add_83310;
  wire [31:0] array_update_83312[10];
  wire [31:0] add_83313;
  wire [31:0] array_update_83314[10][10];
  wire [31:0] array_index_83316[10];
  wire [31:0] array_index_83317[10];
  wire [31:0] smul_83321;
  wire [31:0] add_83323;
  wire [31:0] array_update_83325[10];
  wire [31:0] add_83326;
  wire [31:0] array_update_83327[10][10];
  wire [31:0] array_index_83329[10];
  wire [31:0] array_index_83330[10];
  wire [31:0] smul_83334;
  wire [31:0] add_83336;
  wire [31:0] array_update_83338[10];
  wire [31:0] add_83339;
  wire [31:0] array_update_83340[10][10];
  wire [31:0] array_index_83342[10];
  wire [31:0] array_index_83343[10];
  wire [31:0] smul_83347;
  wire [31:0] add_83349;
  wire [31:0] array_update_83351[10];
  wire [31:0] add_83352;
  wire [31:0] array_update_83353[10][10];
  wire [31:0] array_index_83355[10];
  wire [31:0] array_index_83356[10];
  wire [31:0] smul_83360;
  wire [31:0] add_83362;
  wire [31:0] array_update_83363[10];
  wire [31:0] array_update_83364[10][10];
  wire [31:0] array_index_83366[10];
  wire [31:0] add_83368;
  wire [31:0] array_update_83369[10];
  wire [31:0] literal_83370;
  wire [31:0] array_update_83371[10][10];
  wire [31:0] array_index_83373[10];
  wire [31:0] array_index_83374[10];
  wire [31:0] smul_83378;
  wire [31:0] add_83380;
  wire [31:0] array_update_83382[10];
  wire [31:0] add_83383;
  wire [31:0] array_update_83384[10][10];
  wire [31:0] array_index_83386[10];
  wire [31:0] array_index_83387[10];
  wire [31:0] smul_83391;
  wire [31:0] add_83393;
  wire [31:0] array_update_83395[10];
  wire [31:0] add_83396;
  wire [31:0] array_update_83397[10][10];
  wire [31:0] array_index_83399[10];
  wire [31:0] array_index_83400[10];
  wire [31:0] smul_83404;
  wire [31:0] add_83406;
  wire [31:0] array_update_83408[10];
  wire [31:0] add_83409;
  wire [31:0] array_update_83410[10][10];
  wire [31:0] array_index_83412[10];
  wire [31:0] array_index_83413[10];
  wire [31:0] smul_83417;
  wire [31:0] add_83419;
  wire [31:0] array_update_83421[10];
  wire [31:0] add_83422;
  wire [31:0] array_update_83423[10][10];
  wire [31:0] array_index_83425[10];
  wire [31:0] array_index_83426[10];
  wire [31:0] smul_83430;
  wire [31:0] add_83432;
  wire [31:0] array_update_83434[10];
  wire [31:0] add_83435;
  wire [31:0] array_update_83436[10][10];
  wire [31:0] array_index_83438[10];
  wire [31:0] array_index_83439[10];
  wire [31:0] smul_83443;
  wire [31:0] add_83445;
  wire [31:0] array_update_83447[10];
  wire [31:0] add_83448;
  wire [31:0] array_update_83449[10][10];
  wire [31:0] array_index_83451[10];
  wire [31:0] array_index_83452[10];
  wire [31:0] smul_83456;
  wire [31:0] add_83458;
  wire [31:0] array_update_83460[10];
  wire [31:0] add_83461;
  wire [31:0] array_update_83462[10][10];
  wire [31:0] array_index_83464[10];
  wire [31:0] array_index_83465[10];
  wire [31:0] smul_83469;
  wire [31:0] add_83471;
  wire [31:0] array_update_83473[10];
  wire [31:0] add_83474;
  wire [31:0] array_update_83475[10][10];
  wire [31:0] array_index_83477[10];
  wire [31:0] array_index_83478[10];
  wire [31:0] smul_83482;
  wire [31:0] add_83484;
  wire [31:0] array_update_83486[10];
  wire [31:0] add_83487;
  wire [31:0] array_update_83488[10][10];
  wire [31:0] array_index_83490[10];
  wire [31:0] array_index_83491[10];
  wire [31:0] smul_83495;
  wire [31:0] add_83497;
  wire [31:0] array_update_83498[10];
  wire [31:0] array_update_83499[10][10];
  wire [31:0] array_index_83501[10];
  wire [31:0] add_83503;
  wire [31:0] array_update_83504[10];
  wire [31:0] literal_83505;
  wire [31:0] array_update_83506[10][10];
  wire [31:0] array_index_83508[10];
  wire [31:0] array_index_83509[10];
  wire [31:0] smul_83513;
  wire [31:0] add_83515;
  wire [31:0] array_update_83517[10];
  wire [31:0] add_83518;
  wire [31:0] array_update_83519[10][10];
  wire [31:0] array_index_83521[10];
  wire [31:0] array_index_83522[10];
  wire [31:0] smul_83526;
  wire [31:0] add_83528;
  wire [31:0] array_update_83530[10];
  wire [31:0] add_83531;
  wire [31:0] array_update_83532[10][10];
  wire [31:0] array_index_83534[10];
  wire [31:0] array_index_83535[10];
  wire [31:0] smul_83539;
  wire [31:0] add_83541;
  wire [31:0] array_update_83543[10];
  wire [31:0] add_83544;
  wire [31:0] array_update_83545[10][10];
  wire [31:0] array_index_83547[10];
  wire [31:0] array_index_83548[10];
  wire [31:0] smul_83552;
  wire [31:0] add_83554;
  wire [31:0] array_update_83556[10];
  wire [31:0] add_83557;
  wire [31:0] array_update_83558[10][10];
  wire [31:0] array_index_83560[10];
  wire [31:0] array_index_83561[10];
  wire [31:0] smul_83565;
  wire [31:0] add_83567;
  wire [31:0] array_update_83569[10];
  wire [31:0] add_83570;
  wire [31:0] array_update_83571[10][10];
  wire [31:0] array_index_83573[10];
  wire [31:0] array_index_83574[10];
  wire [31:0] smul_83578;
  wire [31:0] add_83580;
  wire [31:0] array_update_83582[10];
  wire [31:0] add_83583;
  wire [31:0] array_update_83584[10][10];
  wire [31:0] array_index_83586[10];
  wire [31:0] array_index_83587[10];
  wire [31:0] smul_83591;
  wire [31:0] add_83593;
  wire [31:0] array_update_83595[10];
  wire [31:0] add_83596;
  wire [31:0] array_update_83597[10][10];
  wire [31:0] array_index_83599[10];
  wire [31:0] array_index_83600[10];
  wire [31:0] smul_83604;
  wire [31:0] add_83606;
  wire [31:0] array_update_83608[10];
  wire [31:0] add_83609;
  wire [31:0] array_update_83610[10][10];
  wire [31:0] array_index_83612[10];
  wire [31:0] array_index_83613[10];
  wire [31:0] smul_83617;
  wire [31:0] add_83619;
  wire [31:0] array_update_83621[10];
  wire [31:0] add_83622;
  wire [31:0] array_update_83623[10][10];
  wire [31:0] array_index_83625[10];
  wire [31:0] array_index_83626[10];
  wire [31:0] smul_83630;
  wire [31:0] add_83632;
  wire [31:0] array_update_83633[10];
  wire [31:0] array_update_83634[10][10];
  wire [31:0] array_index_83636[10];
  wire [31:0] add_83638;
  wire [31:0] array_update_83639[10];
  wire [31:0] literal_83640;
  wire [31:0] array_update_83641[10][10];
  wire [31:0] array_index_83643[10];
  wire [31:0] array_index_83644[10];
  wire [31:0] smul_83648;
  wire [31:0] add_83650;
  wire [31:0] array_update_83652[10];
  wire [31:0] add_83653;
  wire [31:0] array_update_83654[10][10];
  wire [31:0] array_index_83656[10];
  wire [31:0] array_index_83657[10];
  wire [31:0] smul_83661;
  wire [31:0] add_83663;
  wire [31:0] array_update_83665[10];
  wire [31:0] add_83666;
  wire [31:0] array_update_83667[10][10];
  wire [31:0] array_index_83669[10];
  wire [31:0] array_index_83670[10];
  wire [31:0] smul_83674;
  wire [31:0] add_83676;
  wire [31:0] array_update_83678[10];
  wire [31:0] add_83679;
  wire [31:0] array_update_83680[10][10];
  wire [31:0] array_index_83682[10];
  wire [31:0] array_index_83683[10];
  wire [31:0] smul_83687;
  wire [31:0] add_83689;
  wire [31:0] array_update_83691[10];
  wire [31:0] add_83692;
  wire [31:0] array_update_83693[10][10];
  wire [31:0] array_index_83695[10];
  wire [31:0] array_index_83696[10];
  wire [31:0] smul_83700;
  wire [31:0] add_83702;
  wire [31:0] array_update_83704[10];
  wire [31:0] add_83705;
  wire [31:0] array_update_83706[10][10];
  wire [31:0] array_index_83708[10];
  wire [31:0] array_index_83709[10];
  wire [31:0] smul_83713;
  wire [31:0] add_83715;
  wire [31:0] array_update_83717[10];
  wire [31:0] add_83718;
  wire [31:0] array_update_83719[10][10];
  wire [31:0] array_index_83721[10];
  wire [31:0] array_index_83722[10];
  wire [31:0] smul_83726;
  wire [31:0] add_83728;
  wire [31:0] array_update_83730[10];
  wire [31:0] add_83731;
  wire [31:0] array_update_83732[10][10];
  wire [31:0] array_index_83734[10];
  wire [31:0] array_index_83735[10];
  wire [31:0] smul_83739;
  wire [31:0] add_83741;
  wire [31:0] array_update_83743[10];
  wire [31:0] add_83744;
  wire [31:0] array_update_83745[10][10];
  wire [31:0] array_index_83747[10];
  wire [31:0] array_index_83748[10];
  wire [31:0] smul_83752;
  wire [31:0] add_83754;
  wire [31:0] array_update_83756[10];
  wire [31:0] add_83757;
  wire [31:0] array_update_83758[10][10];
  wire [31:0] array_index_83760[10];
  wire [31:0] array_index_83761[10];
  wire [31:0] smul_83765;
  wire [31:0] add_83767;
  wire [31:0] array_update_83768[10];
  wire [31:0] array_update_83769[10][10];
  wire [31:0] array_index_83771[10];
  wire [31:0] add_83773;
  wire [31:0] array_update_83774[10];
  wire [31:0] literal_83775;
  wire [31:0] array_update_83776[10][10];
  wire [31:0] array_index_83778[10];
  wire [31:0] array_index_83779[10];
  wire [31:0] smul_83783;
  wire [31:0] add_83785;
  wire [31:0] array_update_83787[10];
  wire [31:0] add_83788;
  wire [31:0] array_update_83789[10][10];
  wire [31:0] array_index_83791[10];
  wire [31:0] array_index_83792[10];
  wire [31:0] smul_83796;
  wire [31:0] add_83798;
  wire [31:0] array_update_83800[10];
  wire [31:0] add_83801;
  wire [31:0] array_update_83802[10][10];
  wire [31:0] array_index_83804[10];
  wire [31:0] array_index_83805[10];
  wire [31:0] smul_83809;
  wire [31:0] add_83811;
  wire [31:0] array_update_83813[10];
  wire [31:0] add_83814;
  wire [31:0] array_update_83815[10][10];
  wire [31:0] array_index_83817[10];
  wire [31:0] array_index_83818[10];
  wire [31:0] smul_83822;
  wire [31:0] add_83824;
  wire [31:0] array_update_83826[10];
  wire [31:0] add_83827;
  wire [31:0] array_update_83828[10][10];
  wire [31:0] array_index_83830[10];
  wire [31:0] array_index_83831[10];
  wire [31:0] smul_83835;
  wire [31:0] add_83837;
  wire [31:0] array_update_83839[10];
  wire [31:0] add_83840;
  wire [31:0] array_update_83841[10][10];
  wire [31:0] array_index_83843[10];
  wire [31:0] array_index_83844[10];
  wire [31:0] smul_83848;
  wire [31:0] add_83850;
  wire [31:0] array_update_83852[10];
  wire [31:0] add_83853;
  wire [31:0] array_update_83854[10][10];
  wire [31:0] array_index_83856[10];
  wire [31:0] array_index_83857[10];
  wire [31:0] smul_83861;
  wire [31:0] add_83863;
  wire [31:0] array_update_83865[10];
  wire [31:0] add_83866;
  wire [31:0] array_update_83867[10][10];
  wire [31:0] array_index_83869[10];
  wire [31:0] array_index_83870[10];
  wire [31:0] smul_83874;
  wire [31:0] add_83876;
  wire [31:0] array_update_83878[10];
  wire [31:0] add_83879;
  wire [31:0] array_update_83880[10][10];
  wire [31:0] array_index_83882[10];
  wire [31:0] array_index_83883[10];
  wire [31:0] smul_83887;
  wire [31:0] add_83889;
  wire [31:0] array_update_83891[10];
  wire [31:0] add_83892;
  wire [31:0] array_update_83893[10][10];
  wire [31:0] array_index_83895[10];
  wire [31:0] array_index_83896[10];
  wire [31:0] smul_83900;
  wire [31:0] add_83902;
  wire [31:0] array_update_83903[10];
  wire [31:0] array_update_83904[10][10];
  wire [31:0] array_index_83906[10];
  wire [31:0] add_83908;
  wire [31:0] array_update_83909[10];
  wire [31:0] literal_83910;
  wire [31:0] array_update_83911[10][10];
  wire [31:0] array_index_83913[10];
  wire [31:0] array_index_83914[10];
  wire [31:0] smul_83918;
  wire [31:0] add_83920;
  wire [31:0] array_update_83922[10];
  wire [31:0] add_83923;
  wire [31:0] array_update_83924[10][10];
  wire [31:0] array_index_83926[10];
  wire [31:0] array_index_83927[10];
  wire [31:0] smul_83931;
  wire [31:0] add_83933;
  wire [31:0] array_update_83935[10];
  wire [31:0] add_83936;
  wire [31:0] array_update_83937[10][10];
  wire [31:0] array_index_83939[10];
  wire [31:0] array_index_83940[10];
  wire [31:0] smul_83944;
  wire [31:0] add_83946;
  wire [31:0] array_update_83948[10];
  wire [31:0] add_83949;
  wire [31:0] array_update_83950[10][10];
  wire [31:0] array_index_83952[10];
  wire [31:0] array_index_83953[10];
  wire [31:0] smul_83957;
  wire [31:0] add_83959;
  wire [31:0] array_update_83961[10];
  wire [31:0] add_83962;
  wire [31:0] array_update_83963[10][10];
  wire [31:0] array_index_83965[10];
  wire [31:0] array_index_83966[10];
  wire [31:0] smul_83970;
  wire [31:0] add_83972;
  wire [31:0] array_update_83974[10];
  wire [31:0] add_83975;
  wire [31:0] array_update_83976[10][10];
  wire [31:0] array_index_83978[10];
  wire [31:0] array_index_83979[10];
  wire [31:0] smul_83983;
  wire [31:0] add_83985;
  wire [31:0] array_update_83987[10];
  wire [31:0] add_83988;
  wire [31:0] array_update_83989[10][10];
  wire [31:0] array_index_83991[10];
  wire [31:0] array_index_83992[10];
  wire [31:0] smul_83996;
  wire [31:0] add_83998;
  wire [31:0] array_update_84000[10];
  wire [31:0] add_84001;
  wire [31:0] array_update_84002[10][10];
  wire [31:0] array_index_84004[10];
  wire [31:0] array_index_84005[10];
  wire [31:0] smul_84009;
  wire [31:0] add_84011;
  wire [31:0] array_update_84013[10];
  wire [31:0] add_84014;
  wire [31:0] array_update_84015[10][10];
  wire [31:0] array_index_84017[10];
  wire [31:0] array_index_84018[10];
  wire [31:0] smul_84022;
  wire [31:0] add_84024;
  wire [31:0] array_update_84026[10];
  wire [31:0] add_84027;
  wire [31:0] array_update_84028[10][10];
  wire [31:0] array_index_84030[10];
  wire [31:0] array_index_84031[10];
  wire [31:0] smul_84035;
  wire [31:0] add_84037;
  wire [31:0] array_update_84038[10];
  wire [31:0] array_update_84039[10][10];
  wire [31:0] array_index_84041[10];
  wire [31:0] add_84043;
  wire [31:0] array_update_84044[10];
  wire [31:0] literal_84045;
  wire [31:0] array_update_84046[10][10];
  wire [31:0] array_index_84048[10];
  wire [31:0] array_index_84049[10];
  wire [31:0] smul_84053;
  wire [31:0] add_84055;
  wire [31:0] array_update_84057[10];
  wire [31:0] add_84058;
  wire [31:0] array_update_84059[10][10];
  wire [31:0] array_index_84061[10];
  wire [31:0] array_index_84062[10];
  wire [31:0] smul_84066;
  wire [31:0] add_84068;
  wire [31:0] array_update_84070[10];
  wire [31:0] add_84071;
  wire [31:0] array_update_84072[10][10];
  wire [31:0] array_index_84074[10];
  wire [31:0] array_index_84075[10];
  wire [31:0] smul_84079;
  wire [31:0] add_84081;
  wire [31:0] array_update_84083[10];
  wire [31:0] add_84084;
  wire [31:0] array_update_84085[10][10];
  wire [31:0] array_index_84087[10];
  wire [31:0] array_index_84088[10];
  wire [31:0] smul_84092;
  wire [31:0] add_84094;
  wire [31:0] array_update_84096[10];
  wire [31:0] add_84097;
  wire [31:0] array_update_84098[10][10];
  wire [31:0] array_index_84100[10];
  wire [31:0] array_index_84101[10];
  wire [31:0] smul_84105;
  wire [31:0] add_84107;
  wire [31:0] array_update_84109[10];
  wire [31:0] add_84110;
  wire [31:0] array_update_84111[10][10];
  wire [31:0] array_index_84113[10];
  wire [31:0] array_index_84114[10];
  wire [31:0] smul_84118;
  wire [31:0] add_84120;
  wire [31:0] array_update_84122[10];
  wire [31:0] add_84123;
  wire [31:0] array_update_84124[10][10];
  wire [31:0] array_index_84126[10];
  wire [31:0] array_index_84127[10];
  wire [31:0] smul_84131;
  wire [31:0] add_84133;
  wire [31:0] array_update_84135[10];
  wire [31:0] add_84136;
  wire [31:0] array_update_84137[10][10];
  wire [31:0] array_index_84139[10];
  wire [31:0] array_index_84140[10];
  wire [31:0] smul_84144;
  wire [31:0] add_84146;
  wire [31:0] array_update_84148[10];
  wire [31:0] add_84149;
  wire [31:0] array_update_84150[10][10];
  wire [31:0] array_index_84152[10];
  wire [31:0] array_index_84153[10];
  wire [31:0] smul_84157;
  wire [31:0] add_84159;
  wire [31:0] array_update_84161[10];
  wire [31:0] add_84162;
  wire [31:0] array_update_84163[10][10];
  wire [31:0] array_index_84165[10];
  wire [31:0] array_index_84166[10];
  wire [31:0] smul_84170;
  wire [31:0] add_84172;
  wire [31:0] array_update_84173[10];
  wire [31:0] array_update_84175[10][10];
  wire [31:0] add_84176;
  wire [31:0] array_index_84177[10];
  wire [31:0] literal_84179;
  wire [31:0] array_update_84180[10];
  wire [31:0] literal_84181;
  wire [31:0] array_update_84182[10][10];
  wire [31:0] array_index_84183[10];
  wire [31:0] array_index_84184[10];
  wire [31:0] array_index_84185[10];
  wire [31:0] smul_84189;
  wire [31:0] add_84191;
  wire [31:0] array_update_84193[10];
  wire [31:0] add_84194;
  wire [31:0] array_update_84195[10][10];
  wire [31:0] array_index_84197[10];
  wire [31:0] array_index_84198[10];
  wire [31:0] smul_84202;
  wire [31:0] add_84204;
  wire [31:0] array_update_84206[10];
  wire [31:0] add_84207;
  wire [31:0] array_update_84208[10][10];
  wire [31:0] array_index_84210[10];
  wire [31:0] array_index_84211[10];
  wire [31:0] smul_84215;
  wire [31:0] add_84217;
  wire [31:0] array_update_84219[10];
  wire [31:0] add_84220;
  wire [31:0] array_update_84221[10][10];
  wire [31:0] array_index_84223[10];
  wire [31:0] array_index_84224[10];
  wire [31:0] smul_84228;
  wire [31:0] add_84230;
  wire [31:0] array_update_84232[10];
  wire [31:0] add_84233;
  wire [31:0] array_update_84234[10][10];
  wire [31:0] array_index_84236[10];
  wire [31:0] array_index_84237[10];
  wire [31:0] smul_84241;
  wire [31:0] add_84243;
  wire [31:0] array_update_84245[10];
  wire [31:0] add_84246;
  wire [31:0] array_update_84247[10][10];
  wire [31:0] array_index_84249[10];
  wire [31:0] array_index_84250[10];
  wire [31:0] smul_84254;
  wire [31:0] add_84256;
  wire [31:0] array_update_84258[10];
  wire [31:0] add_84259;
  wire [31:0] array_update_84260[10][10];
  wire [31:0] array_index_84262[10];
  wire [31:0] array_index_84263[10];
  wire [31:0] smul_84267;
  wire [31:0] add_84269;
  wire [31:0] array_update_84271[10];
  wire [31:0] add_84272;
  wire [31:0] array_update_84273[10][10];
  wire [31:0] array_index_84275[10];
  wire [31:0] array_index_84276[10];
  wire [31:0] smul_84280;
  wire [31:0] add_84282;
  wire [31:0] array_update_84284[10];
  wire [31:0] add_84285;
  wire [31:0] array_update_84286[10][10];
  wire [31:0] array_index_84288[10];
  wire [31:0] array_index_84289[10];
  wire [31:0] smul_84293;
  wire [31:0] add_84295;
  wire [31:0] array_update_84297[10];
  wire [31:0] add_84298;
  wire [31:0] array_update_84299[10][10];
  wire [31:0] array_index_84301[10];
  wire [31:0] array_index_84302[10];
  wire [31:0] smul_84306;
  wire [31:0] add_84308;
  wire [31:0] array_update_84309[10];
  wire [31:0] array_update_84310[10][10];
  wire [31:0] array_index_84312[10];
  wire [31:0] add_84314;
  wire [31:0] array_update_84315[10];
  wire [31:0] literal_84316;
  wire [31:0] array_update_84317[10][10];
  wire [31:0] array_index_84319[10];
  wire [31:0] array_index_84320[10];
  wire [31:0] smul_84324;
  wire [31:0] add_84326;
  wire [31:0] array_update_84328[10];
  wire [31:0] add_84329;
  wire [31:0] array_update_84330[10][10];
  wire [31:0] array_index_84332[10];
  wire [31:0] array_index_84333[10];
  wire [31:0] smul_84337;
  wire [31:0] add_84339;
  wire [31:0] array_update_84341[10];
  wire [31:0] add_84342;
  wire [31:0] array_update_84343[10][10];
  wire [31:0] array_index_84345[10];
  wire [31:0] array_index_84346[10];
  wire [31:0] smul_84350;
  wire [31:0] add_84352;
  wire [31:0] array_update_84354[10];
  wire [31:0] add_84355;
  wire [31:0] array_update_84356[10][10];
  wire [31:0] array_index_84358[10];
  wire [31:0] array_index_84359[10];
  wire [31:0] smul_84363;
  wire [31:0] add_84365;
  wire [31:0] array_update_84367[10];
  wire [31:0] add_84368;
  wire [31:0] array_update_84369[10][10];
  wire [31:0] array_index_84371[10];
  wire [31:0] array_index_84372[10];
  wire [31:0] smul_84376;
  wire [31:0] add_84378;
  wire [31:0] array_update_84380[10];
  wire [31:0] add_84381;
  wire [31:0] array_update_84382[10][10];
  wire [31:0] array_index_84384[10];
  wire [31:0] array_index_84385[10];
  wire [31:0] smul_84389;
  wire [31:0] add_84391;
  wire [31:0] array_update_84393[10];
  wire [31:0] add_84394;
  wire [31:0] array_update_84395[10][10];
  wire [31:0] array_index_84397[10];
  wire [31:0] array_index_84398[10];
  wire [31:0] smul_84402;
  wire [31:0] add_84404;
  wire [31:0] array_update_84406[10];
  wire [31:0] add_84407;
  wire [31:0] array_update_84408[10][10];
  wire [31:0] array_index_84410[10];
  wire [31:0] array_index_84411[10];
  wire [31:0] smul_84415;
  wire [31:0] add_84417;
  wire [31:0] array_update_84419[10];
  wire [31:0] add_84420;
  wire [31:0] array_update_84421[10][10];
  wire [31:0] array_index_84423[10];
  wire [31:0] array_index_84424[10];
  wire [31:0] smul_84428;
  wire [31:0] add_84430;
  wire [31:0] array_update_84432[10];
  wire [31:0] add_84433;
  wire [31:0] array_update_84434[10][10];
  wire [31:0] array_index_84436[10];
  wire [31:0] array_index_84437[10];
  wire [31:0] smul_84441;
  wire [31:0] add_84443;
  wire [31:0] array_update_84444[10];
  wire [31:0] array_update_84445[10][10];
  wire [31:0] array_index_84447[10];
  wire [31:0] add_84449;
  wire [31:0] array_update_84450[10];
  wire [31:0] literal_84451;
  wire [31:0] array_update_84452[10][10];
  wire [31:0] array_index_84454[10];
  wire [31:0] array_index_84455[10];
  wire [31:0] smul_84459;
  wire [31:0] add_84461;
  wire [31:0] array_update_84463[10];
  wire [31:0] add_84464;
  wire [31:0] array_update_84465[10][10];
  wire [31:0] array_index_84467[10];
  wire [31:0] array_index_84468[10];
  wire [31:0] smul_84472;
  wire [31:0] add_84474;
  wire [31:0] array_update_84476[10];
  wire [31:0] add_84477;
  wire [31:0] array_update_84478[10][10];
  wire [31:0] array_index_84480[10];
  wire [31:0] array_index_84481[10];
  wire [31:0] smul_84485;
  wire [31:0] add_84487;
  wire [31:0] array_update_84489[10];
  wire [31:0] add_84490;
  wire [31:0] array_update_84491[10][10];
  wire [31:0] array_index_84493[10];
  wire [31:0] array_index_84494[10];
  wire [31:0] smul_84498;
  wire [31:0] add_84500;
  wire [31:0] array_update_84502[10];
  wire [31:0] add_84503;
  wire [31:0] array_update_84504[10][10];
  wire [31:0] array_index_84506[10];
  wire [31:0] array_index_84507[10];
  wire [31:0] smul_84511;
  wire [31:0] add_84513;
  wire [31:0] array_update_84515[10];
  wire [31:0] add_84516;
  wire [31:0] array_update_84517[10][10];
  wire [31:0] array_index_84519[10];
  wire [31:0] array_index_84520[10];
  wire [31:0] smul_84524;
  wire [31:0] add_84526;
  wire [31:0] array_update_84528[10];
  wire [31:0] add_84529;
  wire [31:0] array_update_84530[10][10];
  wire [31:0] array_index_84532[10];
  wire [31:0] array_index_84533[10];
  wire [31:0] smul_84537;
  wire [31:0] add_84539;
  wire [31:0] array_update_84541[10];
  wire [31:0] add_84542;
  wire [31:0] array_update_84543[10][10];
  wire [31:0] array_index_84545[10];
  wire [31:0] array_index_84546[10];
  wire [31:0] smul_84550;
  wire [31:0] add_84552;
  wire [31:0] array_update_84554[10];
  wire [31:0] add_84555;
  wire [31:0] array_update_84556[10][10];
  wire [31:0] array_index_84558[10];
  wire [31:0] array_index_84559[10];
  wire [31:0] smul_84563;
  wire [31:0] add_84565;
  wire [31:0] array_update_84567[10];
  wire [31:0] add_84568;
  wire [31:0] array_update_84569[10][10];
  wire [31:0] array_index_84571[10];
  wire [31:0] array_index_84572[10];
  wire [31:0] smul_84576;
  wire [31:0] add_84578;
  wire [31:0] array_update_84579[10];
  wire [31:0] array_update_84580[10][10];
  wire [31:0] array_index_84582[10];
  wire [31:0] add_84584;
  wire [31:0] array_update_84585[10];
  wire [31:0] literal_84586;
  wire [31:0] array_update_84587[10][10];
  wire [31:0] array_index_84589[10];
  wire [31:0] array_index_84590[10];
  wire [31:0] smul_84594;
  wire [31:0] add_84596;
  wire [31:0] array_update_84598[10];
  wire [31:0] add_84599;
  wire [31:0] array_update_84600[10][10];
  wire [31:0] array_index_84602[10];
  wire [31:0] array_index_84603[10];
  wire [31:0] smul_84607;
  wire [31:0] add_84609;
  wire [31:0] array_update_84611[10];
  wire [31:0] add_84612;
  wire [31:0] array_update_84613[10][10];
  wire [31:0] array_index_84615[10];
  wire [31:0] array_index_84616[10];
  wire [31:0] smul_84620;
  wire [31:0] add_84622;
  wire [31:0] array_update_84624[10];
  wire [31:0] add_84625;
  wire [31:0] array_update_84626[10][10];
  wire [31:0] array_index_84628[10];
  wire [31:0] array_index_84629[10];
  wire [31:0] smul_84633;
  wire [31:0] add_84635;
  wire [31:0] array_update_84637[10];
  wire [31:0] add_84638;
  wire [31:0] array_update_84639[10][10];
  wire [31:0] array_index_84641[10];
  wire [31:0] array_index_84642[10];
  wire [31:0] smul_84646;
  wire [31:0] add_84648;
  wire [31:0] array_update_84650[10];
  wire [31:0] add_84651;
  wire [31:0] array_update_84652[10][10];
  wire [31:0] array_index_84654[10];
  wire [31:0] array_index_84655[10];
  wire [31:0] smul_84659;
  wire [31:0] add_84661;
  wire [31:0] array_update_84663[10];
  wire [31:0] add_84664;
  wire [31:0] array_update_84665[10][10];
  wire [31:0] array_index_84667[10];
  wire [31:0] array_index_84668[10];
  wire [31:0] smul_84672;
  wire [31:0] add_84674;
  wire [31:0] array_update_84676[10];
  wire [31:0] add_84677;
  wire [31:0] array_update_84678[10][10];
  wire [31:0] array_index_84680[10];
  wire [31:0] array_index_84681[10];
  wire [31:0] smul_84685;
  wire [31:0] add_84687;
  wire [31:0] array_update_84689[10];
  wire [31:0] add_84690;
  wire [31:0] array_update_84691[10][10];
  wire [31:0] array_index_84693[10];
  wire [31:0] array_index_84694[10];
  wire [31:0] smul_84698;
  wire [31:0] add_84700;
  wire [31:0] array_update_84702[10];
  wire [31:0] add_84703;
  wire [31:0] array_update_84704[10][10];
  wire [31:0] array_index_84706[10];
  wire [31:0] array_index_84707[10];
  wire [31:0] smul_84711;
  wire [31:0] add_84713;
  wire [31:0] array_update_84714[10];
  wire [31:0] array_update_84715[10][10];
  wire [31:0] array_index_84717[10];
  wire [31:0] add_84719;
  wire [31:0] array_update_84720[10];
  wire [31:0] literal_84721;
  wire [31:0] array_update_84722[10][10];
  wire [31:0] array_index_84724[10];
  wire [31:0] array_index_84725[10];
  wire [31:0] smul_84729;
  wire [31:0] add_84731;
  wire [31:0] array_update_84733[10];
  wire [31:0] add_84734;
  wire [31:0] array_update_84735[10][10];
  wire [31:0] array_index_84737[10];
  wire [31:0] array_index_84738[10];
  wire [31:0] smul_84742;
  wire [31:0] add_84744;
  wire [31:0] array_update_84746[10];
  wire [31:0] add_84747;
  wire [31:0] array_update_84748[10][10];
  wire [31:0] array_index_84750[10];
  wire [31:0] array_index_84751[10];
  wire [31:0] smul_84755;
  wire [31:0] add_84757;
  wire [31:0] array_update_84759[10];
  wire [31:0] add_84760;
  wire [31:0] array_update_84761[10][10];
  wire [31:0] array_index_84763[10];
  wire [31:0] array_index_84764[10];
  wire [31:0] smul_84768;
  wire [31:0] add_84770;
  wire [31:0] array_update_84772[10];
  wire [31:0] add_84773;
  wire [31:0] array_update_84774[10][10];
  wire [31:0] array_index_84776[10];
  wire [31:0] array_index_84777[10];
  wire [31:0] smul_84781;
  wire [31:0] add_84783;
  wire [31:0] array_update_84785[10];
  wire [31:0] add_84786;
  wire [31:0] array_update_84787[10][10];
  wire [31:0] array_index_84789[10];
  wire [31:0] array_index_84790[10];
  wire [31:0] smul_84794;
  wire [31:0] add_84796;
  wire [31:0] array_update_84798[10];
  wire [31:0] add_84799;
  wire [31:0] array_update_84800[10][10];
  wire [31:0] array_index_84802[10];
  wire [31:0] array_index_84803[10];
  wire [31:0] smul_84807;
  wire [31:0] add_84809;
  wire [31:0] array_update_84811[10];
  wire [31:0] add_84812;
  wire [31:0] array_update_84813[10][10];
  wire [31:0] array_index_84815[10];
  wire [31:0] array_index_84816[10];
  wire [31:0] smul_84820;
  wire [31:0] add_84822;
  wire [31:0] array_update_84824[10];
  wire [31:0] add_84825;
  wire [31:0] array_update_84826[10][10];
  wire [31:0] array_index_84828[10];
  wire [31:0] array_index_84829[10];
  wire [31:0] smul_84833;
  wire [31:0] add_84835;
  wire [31:0] array_update_84837[10];
  wire [31:0] add_84838;
  wire [31:0] array_update_84839[10][10];
  wire [31:0] array_index_84841[10];
  wire [31:0] array_index_84842[10];
  wire [31:0] smul_84846;
  wire [31:0] add_84848;
  wire [31:0] array_update_84849[10];
  wire [31:0] array_update_84850[10][10];
  wire [31:0] array_index_84852[10];
  wire [31:0] add_84854;
  wire [31:0] array_update_84855[10];
  wire [31:0] literal_84856;
  wire [31:0] array_update_84857[10][10];
  wire [31:0] array_index_84859[10];
  wire [31:0] array_index_84860[10];
  wire [31:0] smul_84864;
  wire [31:0] add_84866;
  wire [31:0] array_update_84868[10];
  wire [31:0] add_84869;
  wire [31:0] array_update_84870[10][10];
  wire [31:0] array_index_84872[10];
  wire [31:0] array_index_84873[10];
  wire [31:0] smul_84877;
  wire [31:0] add_84879;
  wire [31:0] array_update_84881[10];
  wire [31:0] add_84882;
  wire [31:0] array_update_84883[10][10];
  wire [31:0] array_index_84885[10];
  wire [31:0] array_index_84886[10];
  wire [31:0] smul_84890;
  wire [31:0] add_84892;
  wire [31:0] array_update_84894[10];
  wire [31:0] add_84895;
  wire [31:0] array_update_84896[10][10];
  wire [31:0] array_index_84898[10];
  wire [31:0] array_index_84899[10];
  wire [31:0] smul_84903;
  wire [31:0] add_84905;
  wire [31:0] array_update_84907[10];
  wire [31:0] add_84908;
  wire [31:0] array_update_84909[10][10];
  wire [31:0] array_index_84911[10];
  wire [31:0] array_index_84912[10];
  wire [31:0] smul_84916;
  wire [31:0] add_84918;
  wire [31:0] array_update_84920[10];
  wire [31:0] add_84921;
  wire [31:0] array_update_84922[10][10];
  wire [31:0] array_index_84924[10];
  wire [31:0] array_index_84925[10];
  wire [31:0] smul_84929;
  wire [31:0] add_84931;
  wire [31:0] array_update_84933[10];
  wire [31:0] add_84934;
  wire [31:0] array_update_84935[10][10];
  wire [31:0] array_index_84937[10];
  wire [31:0] array_index_84938[10];
  wire [31:0] smul_84942;
  wire [31:0] add_84944;
  wire [31:0] array_update_84946[10];
  wire [31:0] add_84947;
  wire [31:0] array_update_84948[10][10];
  wire [31:0] array_index_84950[10];
  wire [31:0] array_index_84951[10];
  wire [31:0] smul_84955;
  wire [31:0] add_84957;
  wire [31:0] array_update_84959[10];
  wire [31:0] add_84960;
  wire [31:0] array_update_84961[10][10];
  wire [31:0] array_index_84963[10];
  wire [31:0] array_index_84964[10];
  wire [31:0] smul_84968;
  wire [31:0] add_84970;
  wire [31:0] array_update_84972[10];
  wire [31:0] add_84973;
  wire [31:0] array_update_84974[10][10];
  wire [31:0] array_index_84976[10];
  wire [31:0] array_index_84977[10];
  wire [31:0] smul_84981;
  wire [31:0] add_84983;
  wire [31:0] array_update_84984[10];
  wire [31:0] array_update_84985[10][10];
  wire [31:0] array_index_84987[10];
  wire [31:0] add_84989;
  wire [31:0] array_update_84990[10];
  wire [31:0] literal_84991;
  wire [31:0] array_update_84992[10][10];
  wire [31:0] array_index_84994[10];
  wire [31:0] array_index_84995[10];
  wire [31:0] smul_84999;
  wire [31:0] add_85001;
  wire [31:0] array_update_85003[10];
  wire [31:0] add_85004;
  wire [31:0] array_update_85005[10][10];
  wire [31:0] array_index_85007[10];
  wire [31:0] array_index_85008[10];
  wire [31:0] smul_85012;
  wire [31:0] add_85014;
  wire [31:0] array_update_85016[10];
  wire [31:0] add_85017;
  wire [31:0] array_update_85018[10][10];
  wire [31:0] array_index_85020[10];
  wire [31:0] array_index_85021[10];
  wire [31:0] smul_85025;
  wire [31:0] add_85027;
  wire [31:0] array_update_85029[10];
  wire [31:0] add_85030;
  wire [31:0] array_update_85031[10][10];
  wire [31:0] array_index_85033[10];
  wire [31:0] array_index_85034[10];
  wire [31:0] smul_85038;
  wire [31:0] add_85040;
  wire [31:0] array_update_85042[10];
  wire [31:0] add_85043;
  wire [31:0] array_update_85044[10][10];
  wire [31:0] array_index_85046[10];
  wire [31:0] array_index_85047[10];
  wire [31:0] smul_85051;
  wire [31:0] add_85053;
  wire [31:0] array_update_85055[10];
  wire [31:0] add_85056;
  wire [31:0] array_update_85057[10][10];
  wire [31:0] array_index_85059[10];
  wire [31:0] array_index_85060[10];
  wire [31:0] smul_85064;
  wire [31:0] add_85066;
  wire [31:0] array_update_85068[10];
  wire [31:0] add_85069;
  wire [31:0] array_update_85070[10][10];
  wire [31:0] array_index_85072[10];
  wire [31:0] array_index_85073[10];
  wire [31:0] smul_85077;
  wire [31:0] add_85079;
  wire [31:0] array_update_85081[10];
  wire [31:0] add_85082;
  wire [31:0] array_update_85083[10][10];
  wire [31:0] array_index_85085[10];
  wire [31:0] array_index_85086[10];
  wire [31:0] smul_85090;
  wire [31:0] add_85092;
  wire [31:0] array_update_85094[10];
  wire [31:0] add_85095;
  wire [31:0] array_update_85096[10][10];
  wire [31:0] array_index_85098[10];
  wire [31:0] array_index_85099[10];
  wire [31:0] smul_85103;
  wire [31:0] add_85105;
  wire [31:0] array_update_85107[10];
  wire [31:0] add_85108;
  wire [31:0] array_update_85109[10][10];
  wire [31:0] array_index_85111[10];
  wire [31:0] array_index_85112[10];
  wire [31:0] smul_85116;
  wire [31:0] add_85118;
  wire [31:0] array_update_85119[10];
  wire [31:0] array_update_85120[10][10];
  wire [31:0] array_index_85122[10];
  wire [31:0] add_85124;
  wire [31:0] array_update_85125[10];
  wire [31:0] literal_85126;
  wire [31:0] array_update_85127[10][10];
  wire [31:0] array_index_85129[10];
  wire [31:0] array_index_85130[10];
  wire [31:0] smul_85134;
  wire [31:0] add_85136;
  wire [31:0] array_update_85138[10];
  wire [31:0] add_85139;
  wire [31:0] array_update_85140[10][10];
  wire [31:0] array_index_85142[10];
  wire [31:0] array_index_85143[10];
  wire [31:0] smul_85147;
  wire [31:0] add_85149;
  wire [31:0] array_update_85151[10];
  wire [31:0] add_85152;
  wire [31:0] array_update_85153[10][10];
  wire [31:0] array_index_85155[10];
  wire [31:0] array_index_85156[10];
  wire [31:0] smul_85160;
  wire [31:0] add_85162;
  wire [31:0] array_update_85164[10];
  wire [31:0] add_85165;
  wire [31:0] array_update_85166[10][10];
  wire [31:0] array_index_85168[10];
  wire [31:0] array_index_85169[10];
  wire [31:0] smul_85173;
  wire [31:0] add_85175;
  wire [31:0] array_update_85177[10];
  wire [31:0] add_85178;
  wire [31:0] array_update_85179[10][10];
  wire [31:0] array_index_85181[10];
  wire [31:0] array_index_85182[10];
  wire [31:0] smul_85186;
  wire [31:0] add_85188;
  wire [31:0] array_update_85190[10];
  wire [31:0] add_85191;
  wire [31:0] array_update_85192[10][10];
  wire [31:0] array_index_85194[10];
  wire [31:0] array_index_85195[10];
  wire [31:0] smul_85199;
  wire [31:0] add_85201;
  wire [31:0] array_update_85203[10];
  wire [31:0] add_85204;
  wire [31:0] array_update_85205[10][10];
  wire [31:0] array_index_85207[10];
  wire [31:0] array_index_85208[10];
  wire [31:0] smul_85212;
  wire [31:0] add_85214;
  wire [31:0] array_update_85216[10];
  wire [31:0] add_85217;
  wire [31:0] array_update_85218[10][10];
  wire [31:0] array_index_85220[10];
  wire [31:0] array_index_85221[10];
  wire [31:0] smul_85225;
  wire [31:0] add_85227;
  wire [31:0] array_update_85229[10];
  wire [31:0] add_85230;
  wire [31:0] array_update_85231[10][10];
  wire [31:0] array_index_85233[10];
  wire [31:0] array_index_85234[10];
  wire [31:0] smul_85238;
  wire [31:0] add_85240;
  wire [31:0] array_update_85242[10];
  wire [31:0] add_85243;
  wire [31:0] array_update_85244[10][10];
  wire [31:0] array_index_85246[10];
  wire [31:0] array_index_85247[10];
  wire [31:0] smul_85251;
  wire [31:0] add_85253;
  wire [31:0] array_update_85254[10];
  wire [31:0] array_update_85255[10][10];
  wire [31:0] array_index_85257[10];
  wire [31:0] add_85259;
  wire [31:0] array_update_85260[10];
  wire [31:0] literal_85261;
  wire [31:0] array_update_85262[10][10];
  wire [31:0] array_index_85264[10];
  wire [31:0] array_index_85265[10];
  wire [31:0] smul_85269;
  wire [31:0] add_85271;
  wire [31:0] array_update_85273[10];
  wire [31:0] add_85274;
  wire [31:0] array_update_85275[10][10];
  wire [31:0] array_index_85277[10];
  wire [31:0] array_index_85278[10];
  wire [31:0] smul_85282;
  wire [31:0] add_85284;
  wire [31:0] array_update_85286[10];
  wire [31:0] add_85287;
  wire [31:0] array_update_85288[10][10];
  wire [31:0] array_index_85290[10];
  wire [31:0] array_index_85291[10];
  wire [31:0] smul_85295;
  wire [31:0] add_85297;
  wire [31:0] array_update_85299[10];
  wire [31:0] add_85300;
  wire [31:0] array_update_85301[10][10];
  wire [31:0] array_index_85303[10];
  wire [31:0] array_index_85304[10];
  wire [31:0] smul_85308;
  wire [31:0] add_85310;
  wire [31:0] array_update_85312[10];
  wire [31:0] add_85313;
  wire [31:0] array_update_85314[10][10];
  wire [31:0] array_index_85316[10];
  wire [31:0] array_index_85317[10];
  wire [31:0] smul_85321;
  wire [31:0] add_85323;
  wire [31:0] array_update_85325[10];
  wire [31:0] add_85326;
  wire [31:0] array_update_85327[10][10];
  wire [31:0] array_index_85329[10];
  wire [31:0] array_index_85330[10];
  wire [31:0] smul_85334;
  wire [31:0] add_85336;
  wire [31:0] array_update_85338[10];
  wire [31:0] add_85339;
  wire [31:0] array_update_85340[10][10];
  wire [31:0] array_index_85342[10];
  wire [31:0] array_index_85343[10];
  wire [31:0] smul_85347;
  wire [31:0] add_85349;
  wire [31:0] array_update_85351[10];
  wire [31:0] add_85352;
  wire [31:0] array_update_85353[10][10];
  wire [31:0] array_index_85355[10];
  wire [31:0] array_index_85356[10];
  wire [31:0] smul_85360;
  wire [31:0] add_85362;
  wire [31:0] array_update_85364[10];
  wire [31:0] add_85365;
  wire [31:0] array_update_85366[10][10];
  wire [31:0] array_index_85368[10];
  wire [31:0] array_index_85369[10];
  wire [31:0] smul_85373;
  wire [31:0] add_85375;
  wire [31:0] array_update_85377[10];
  wire [31:0] add_85378;
  wire [31:0] array_update_85379[10][10];
  wire [31:0] array_index_85381[10];
  wire [31:0] array_index_85383[10];
  wire [31:0] smul_85388;
  wire [31:0] add_85391;
  wire [31:0] array_update_85393[10];
  wire [31:0] array_update_85397[10][10];
  wire [31:0] array_index_85401[10];
  wire [31:0] add_85403;
  wire [31:0] array_update_85407[10];
  wire [31:0] literal_85408;
  wire [31:0] array_update_85411[10][10];
  wire [31:0] array_index_85413[10];
  wire [31:0] array_index_85417[10];
  wire [31:0] smul_85423;
  wire [31:0] add_85428;
  wire [31:0] array_update_85432[10];
  wire [31:0] add_85433;
  wire [31:0] array_update_85437[10][10];
  wire [31:0] array_index_85439[10];
  wire [31:0] array_index_85442[10];
  wire [31:0] smul_85449;
  wire [31:0] add_85453;
  wire [31:0] array_update_85458[10];
  wire [31:0] add_85459;
  wire [31:0] array_update_85462[10][10];
  wire [31:0] array_index_85464[10];
  wire [31:0] array_index_85468[10];
  wire [31:0] smul_85474;
  wire [31:0] add_85479;
  wire [31:0] array_update_85502[10];
  wire [31:0] add_85503;
  wire [31:0] array_update_85524[10][10];
  wire [31:0] array_index_85526[10];
  wire [31:0] array_index_85557[10];
  wire [31:0] smul_85581;
  wire [31:0] add_85613;
  wire [31:0] array_update_85635[10];
  wire [31:0] add_85636;
  wire [31:0] array_update_85667[10][10];
  wire [31:0] array_index_85669[10];
  wire [31:0] array_index_85690[10];
  wire [31:0] smul_85724;
  wire [31:0] add_85746;
  wire [31:0] array_update_85778[10];
  wire [31:0] add_85779;
  wire [31:0] array_update_85800[10][10];
  wire [31:0] array_index_85802[10];
  wire [31:0] array_index_85833[10];
  wire [31:0] smul_85857;
  wire [31:0] add_85889;
  wire [31:0] array_update_85911[10];
  wire [31:0] add_85912;
  wire [31:0] array_update_85943[10][10];
  wire [31:0] array_index_85945[10];
  wire [31:0] array_index_85966[10];
  wire [31:0] smul_85991;
  wire [31:0] add_86203;
  wire [31:0] array_update_86405[10];
  wire [31:0] add_86406;
  wire [31:0] array_update_86707[10][10];
  wire [31:0] array_index_86709[10];
  wire [31:0] array_index_86910[10];
  wire [31:0] smul_87214;
  wire [31:0] add_87416;
  wire [31:0] array_update_87718[10];
  wire [31:0] add_87719;
  wire [31:0] array_update_87920[10][10];
  wire [31:0] array_index_87922[10];
  wire [31:0] array_index_88245[10];
  wire [31:0] literal_88243;
  wire [31:0] smul_88471;
  wire [31:0] literal_88223;
  wire [31:0] literal_88225;
  wire [31:0] literal_88227;
  wire [31:0] literal_88229;
  wire [31:0] literal_88231;
  wire [31:0] literal_88233;
  wire [31:0] literal_88235;
  wire [31:0] literal_88237;
  wire [31:0] literal_88239;
  wire [31:0] add_88468;
  wire [31:0] literal_88241;
  wire [31:0] add_88795;
  wire [31:0] add_88448;
  wire [31:0] add_88450;
  wire [31:0] add_88452;
  wire [31:0] add_88454;
  wire [31:0] add_88456;
  wire [31:0] add_88458;
  wire [31:0] add_88460;
  wire [31:0] add_88462;
  wire [31:0] add_88464;
  wire [31:0] add_88792;
  wire [31:0] add_88466;
  wire [31:0] array_update_89019[10];
  wire [31:0] add_89020;
  wire [31:0] add_88772;
  wire [31:0] add_88774;
  wire [31:0] add_88776;
  wire [31:0] add_88778;
  wire [31:0] add_88780;
  wire [31:0] add_88782;
  wire [31:0] add_88784;
  wire [31:0] add_88786;
  wire [31:0] add_88788;
  wire [31:0] add_89017;
  wire [31:0] add_88790;
  wire [31:0] array_update_89343[10][10];
  wire [31:0] array_index_89345[10];
  wire [31:0] add_88997;
  wire [31:0] add_88999;
  wire [31:0] add_89001;
  wire [31:0] add_89003;
  wire [31:0] add_89005;
  wire [31:0] add_89007;
  wire [31:0] add_89009;
  wire [31:0] add_89011;
  wire [31:0] add_89013;
  wire [31:0] add_89341;
  wire [31:0] add_89015;
  wire [31:0] array_index_89572[10];
  wire [31:0] add_89321;
  wire [31:0] add_89323;
  wire [31:0] add_89325;
  wire [31:0] add_89327;
  wire [31:0] add_89329;
  wire [31:0] add_89331;
  wire [31:0] add_89333;
  wire [31:0] add_89335;
  wire [31:0] add_89337;
  wire [31:0] add_89566;
  wire [31:0] add_89339;
  wire [31:0] smul_89899;
  wire [31:0] add_89546;
  wire [31:0] add_89548;
  wire [31:0] add_89550;
  wire [31:0] add_89552;
  wire [31:0] add_89554;
  wire [31:0] add_89556;
  wire [31:0] add_89558;
  wire [31:0] add_89560;
  wire [31:0] add_89562;
  wire [31:0] add_89895;
  wire [31:0] add_89564;
  wire [31:0] add_90127;
  wire [31:0] add_89875;
  wire [31:0] add_89877;
  wire [31:0] add_89879;
  wire [31:0] add_89881;
  wire [31:0] add_89883;
  wire [31:0] add_89885;
  wire [31:0] add_89887;
  wire [31:0] add_89889;
  wire [31:0] add_89891;
  wire [31:0] add_90120;
  wire [31:0] add_89893;
  wire [31:0] array_update_90451[10];
  wire [31:0] add_90100;
  wire [31:0] add_90102;
  wire [31:0] add_90104;
  wire [31:0] add_90106;
  wire [31:0] add_90108;
  wire [31:0] add_90110;
  wire [31:0] add_90112;
  wire [31:0] add_90114;
  wire [31:0] add_90116;
  wire [31:0] add_90448;
  wire [31:0] add_90118;
  wire [31:0] array_update_90811[10][10];
  wire [31:0] add_90428;
  wire [31:0] add_90430;
  wire [31:0] add_90432;
  wire [31:0] add_90434;
  wire [31:0] add_90436;
  wire [31:0] add_90438;
  wire [31:0] add_90440;
  wire [31:0] add_90442;
  wire [31:0] add_90444;
  wire [31:0] add_90805;
  wire [31:0] add_90446;
  wire [31:0] array_index_91514[10];
  wire [31:0] add_90785;
  wire [31:0] array_index_91524[10];
  wire [31:0] add_90787;
  wire [31:0] array_index_91534[10];
  wire [31:0] add_90789;
  wire [31:0] array_index_91544[10];
  wire [31:0] add_90791;
  wire [31:0] array_index_91554[10];
  wire [31:0] add_90793;
  wire [31:0] array_index_91564[10];
  wire [31:0] add_90795;
  wire [31:0] array_index_91574[10];
  wire [31:0] add_90797;
  wire [31:0] array_index_91584[10];
  wire [31:0] add_90799;
  wire [31:0] array_index_91594[10];
  wire [31:0] add_90801;
  wire [31:0] array_index_91604[10];
  wire [31:0] add_90803;
  assign literal_70997 = 32'h0000_0000;
  assign literal_70999 = 32'h0000_0000;
  assign array_index_71000 = literal_70996[literal_70997 > 32'h0000_0009 ? 4'h9 : literal_70997[3:0]];
  assign literal_71001 = 32'h0000_0000;
  assign array_index_71002 = literal_70998[literal_70999 > 32'h0000_0009 ? 4'h9 : literal_70999[3:0]];
  assign literal_71003 = 32'h0000_0000;
  assign array_update_71004[0] = literal_71001 == 32'h0000_0000 ? TestBlock__A_op0 : array_index_71000[0];
  assign array_update_71004[1] = literal_71001 == 32'h0000_0001 ? TestBlock__A_op0 : array_index_71000[1];
  assign array_update_71004[2] = literal_71001 == 32'h0000_0002 ? TestBlock__A_op0 : array_index_71000[2];
  assign array_update_71004[3] = literal_71001 == 32'h0000_0003 ? TestBlock__A_op0 : array_index_71000[3];
  assign array_update_71004[4] = literal_71001 == 32'h0000_0004 ? TestBlock__A_op0 : array_index_71000[4];
  assign array_update_71004[5] = literal_71001 == 32'h0000_0005 ? TestBlock__A_op0 : array_index_71000[5];
  assign array_update_71004[6] = literal_71001 == 32'h0000_0006 ? TestBlock__A_op0 : array_index_71000[6];
  assign array_update_71004[7] = literal_71001 == 32'h0000_0007 ? TestBlock__A_op0 : array_index_71000[7];
  assign array_update_71004[8] = literal_71001 == 32'h0000_0008 ? TestBlock__A_op0 : array_index_71000[8];
  assign array_update_71004[9] = literal_71001 == 32'h0000_0009 ? TestBlock__A_op0 : array_index_71000[9];
  assign array_update_71005[0] = literal_71003 == 32'h0000_0000 ? TestBlock__B_op0 : array_index_71002[0];
  assign array_update_71005[1] = literal_71003 == 32'h0000_0001 ? TestBlock__B_op0 : array_index_71002[1];
  assign array_update_71005[2] = literal_71003 == 32'h0000_0002 ? TestBlock__B_op0 : array_index_71002[2];
  assign array_update_71005[3] = literal_71003 == 32'h0000_0003 ? TestBlock__B_op0 : array_index_71002[3];
  assign array_update_71005[4] = literal_71003 == 32'h0000_0004 ? TestBlock__B_op0 : array_index_71002[4];
  assign array_update_71005[5] = literal_71003 == 32'h0000_0005 ? TestBlock__B_op0 : array_index_71002[5];
  assign array_update_71005[6] = literal_71003 == 32'h0000_0006 ? TestBlock__B_op0 : array_index_71002[6];
  assign array_update_71005[7] = literal_71003 == 32'h0000_0007 ? TestBlock__B_op0 : array_index_71002[7];
  assign array_update_71005[8] = literal_71003 == 32'h0000_0008 ? TestBlock__B_op0 : array_index_71002[8];
  assign array_update_71005[9] = literal_71003 == 32'h0000_0009 ? TestBlock__B_op0 : array_index_71002[9];
  assign array_update_71006[0] = literal_70997 == 32'h0000_0000 ? array_update_71004 : literal_70996[0];
  assign array_update_71006[1] = literal_70997 == 32'h0000_0001 ? array_update_71004 : literal_70996[1];
  assign array_update_71006[2] = literal_70997 == 32'h0000_0002 ? array_update_71004 : literal_70996[2];
  assign array_update_71006[3] = literal_70997 == 32'h0000_0003 ? array_update_71004 : literal_70996[3];
  assign array_update_71006[4] = literal_70997 == 32'h0000_0004 ? array_update_71004 : literal_70996[4];
  assign array_update_71006[5] = literal_70997 == 32'h0000_0005 ? array_update_71004 : literal_70996[5];
  assign array_update_71006[6] = literal_70997 == 32'h0000_0006 ? array_update_71004 : literal_70996[6];
  assign array_update_71006[7] = literal_70997 == 32'h0000_0007 ? array_update_71004 : literal_70996[7];
  assign array_update_71006[8] = literal_70997 == 32'h0000_0008 ? array_update_71004 : literal_70996[8];
  assign array_update_71006[9] = literal_70997 == 32'h0000_0009 ? array_update_71004 : literal_70996[9];
  assign array_update_71008[0] = literal_70999 == 32'h0000_0000 ? array_update_71005 : literal_70998[0];
  assign array_update_71008[1] = literal_70999 == 32'h0000_0001 ? array_update_71005 : literal_70998[1];
  assign array_update_71008[2] = literal_70999 == 32'h0000_0002 ? array_update_71005 : literal_70998[2];
  assign array_update_71008[3] = literal_70999 == 32'h0000_0003 ? array_update_71005 : literal_70998[3];
  assign array_update_71008[4] = literal_70999 == 32'h0000_0004 ? array_update_71005 : literal_70998[4];
  assign array_update_71008[5] = literal_70999 == 32'h0000_0005 ? array_update_71005 : literal_70998[5];
  assign array_update_71008[6] = literal_70999 == 32'h0000_0006 ? array_update_71005 : literal_70998[6];
  assign array_update_71008[7] = literal_70999 == 32'h0000_0007 ? array_update_71005 : literal_70998[7];
  assign array_update_71008[8] = literal_70999 == 32'h0000_0008 ? array_update_71005 : literal_70998[8];
  assign array_update_71008[9] = literal_70999 == 32'h0000_0009 ? array_update_71005 : literal_70998[9];
  assign array_index_71010 = array_update_71006[literal_70997 > 32'h0000_0009 ? 4'h9 : literal_70997[3:0]];
  assign add_71011 = literal_71001 + 32'h0000_0001;
  assign array_index_71012 = array_update_71008[literal_70999 > 32'h0000_0009 ? 4'h9 : literal_70999[3:0]];
  assign add_71013 = literal_71003 + 32'h0000_0001;
  assign array_update_71014[0] = add_71011 == 32'h0000_0000 ? TestBlock__A_op1 : array_index_71010[0];
  assign array_update_71014[1] = add_71011 == 32'h0000_0001 ? TestBlock__A_op1 : array_index_71010[1];
  assign array_update_71014[2] = add_71011 == 32'h0000_0002 ? TestBlock__A_op1 : array_index_71010[2];
  assign array_update_71014[3] = add_71011 == 32'h0000_0003 ? TestBlock__A_op1 : array_index_71010[3];
  assign array_update_71014[4] = add_71011 == 32'h0000_0004 ? TestBlock__A_op1 : array_index_71010[4];
  assign array_update_71014[5] = add_71011 == 32'h0000_0005 ? TestBlock__A_op1 : array_index_71010[5];
  assign array_update_71014[6] = add_71011 == 32'h0000_0006 ? TestBlock__A_op1 : array_index_71010[6];
  assign array_update_71014[7] = add_71011 == 32'h0000_0007 ? TestBlock__A_op1 : array_index_71010[7];
  assign array_update_71014[8] = add_71011 == 32'h0000_0008 ? TestBlock__A_op1 : array_index_71010[8];
  assign array_update_71014[9] = add_71011 == 32'h0000_0009 ? TestBlock__A_op1 : array_index_71010[9];
  assign array_update_71015[0] = add_71013 == 32'h0000_0000 ? TestBlock__B_op1 : array_index_71012[0];
  assign array_update_71015[1] = add_71013 == 32'h0000_0001 ? TestBlock__B_op1 : array_index_71012[1];
  assign array_update_71015[2] = add_71013 == 32'h0000_0002 ? TestBlock__B_op1 : array_index_71012[2];
  assign array_update_71015[3] = add_71013 == 32'h0000_0003 ? TestBlock__B_op1 : array_index_71012[3];
  assign array_update_71015[4] = add_71013 == 32'h0000_0004 ? TestBlock__B_op1 : array_index_71012[4];
  assign array_update_71015[5] = add_71013 == 32'h0000_0005 ? TestBlock__B_op1 : array_index_71012[5];
  assign array_update_71015[6] = add_71013 == 32'h0000_0006 ? TestBlock__B_op1 : array_index_71012[6];
  assign array_update_71015[7] = add_71013 == 32'h0000_0007 ? TestBlock__B_op1 : array_index_71012[7];
  assign array_update_71015[8] = add_71013 == 32'h0000_0008 ? TestBlock__B_op1 : array_index_71012[8];
  assign array_update_71015[9] = add_71013 == 32'h0000_0009 ? TestBlock__B_op1 : array_index_71012[9];
  assign array_update_71016[0] = literal_70997 == 32'h0000_0000 ? array_update_71014 : array_update_71006[0];
  assign array_update_71016[1] = literal_70997 == 32'h0000_0001 ? array_update_71014 : array_update_71006[1];
  assign array_update_71016[2] = literal_70997 == 32'h0000_0002 ? array_update_71014 : array_update_71006[2];
  assign array_update_71016[3] = literal_70997 == 32'h0000_0003 ? array_update_71014 : array_update_71006[3];
  assign array_update_71016[4] = literal_70997 == 32'h0000_0004 ? array_update_71014 : array_update_71006[4];
  assign array_update_71016[5] = literal_70997 == 32'h0000_0005 ? array_update_71014 : array_update_71006[5];
  assign array_update_71016[6] = literal_70997 == 32'h0000_0006 ? array_update_71014 : array_update_71006[6];
  assign array_update_71016[7] = literal_70997 == 32'h0000_0007 ? array_update_71014 : array_update_71006[7];
  assign array_update_71016[8] = literal_70997 == 32'h0000_0008 ? array_update_71014 : array_update_71006[8];
  assign array_update_71016[9] = literal_70997 == 32'h0000_0009 ? array_update_71014 : array_update_71006[9];
  assign array_update_71018[0] = literal_70999 == 32'h0000_0000 ? array_update_71015 : array_update_71008[0];
  assign array_update_71018[1] = literal_70999 == 32'h0000_0001 ? array_update_71015 : array_update_71008[1];
  assign array_update_71018[2] = literal_70999 == 32'h0000_0002 ? array_update_71015 : array_update_71008[2];
  assign array_update_71018[3] = literal_70999 == 32'h0000_0003 ? array_update_71015 : array_update_71008[3];
  assign array_update_71018[4] = literal_70999 == 32'h0000_0004 ? array_update_71015 : array_update_71008[4];
  assign array_update_71018[5] = literal_70999 == 32'h0000_0005 ? array_update_71015 : array_update_71008[5];
  assign array_update_71018[6] = literal_70999 == 32'h0000_0006 ? array_update_71015 : array_update_71008[6];
  assign array_update_71018[7] = literal_70999 == 32'h0000_0007 ? array_update_71015 : array_update_71008[7];
  assign array_update_71018[8] = literal_70999 == 32'h0000_0008 ? array_update_71015 : array_update_71008[8];
  assign array_update_71018[9] = literal_70999 == 32'h0000_0009 ? array_update_71015 : array_update_71008[9];
  assign array_index_71020 = array_update_71016[literal_70997 > 32'h0000_0009 ? 4'h9 : literal_70997[3:0]];
  assign add_71021 = add_71011 + 32'h0000_0001;
  assign array_index_71022 = array_update_71018[literal_70999 > 32'h0000_0009 ? 4'h9 : literal_70999[3:0]];
  assign add_71023 = add_71013 + 32'h0000_0001;
  assign array_update_71024[0] = add_71021 == 32'h0000_0000 ? TestBlock__A_op2 : array_index_71020[0];
  assign array_update_71024[1] = add_71021 == 32'h0000_0001 ? TestBlock__A_op2 : array_index_71020[1];
  assign array_update_71024[2] = add_71021 == 32'h0000_0002 ? TestBlock__A_op2 : array_index_71020[2];
  assign array_update_71024[3] = add_71021 == 32'h0000_0003 ? TestBlock__A_op2 : array_index_71020[3];
  assign array_update_71024[4] = add_71021 == 32'h0000_0004 ? TestBlock__A_op2 : array_index_71020[4];
  assign array_update_71024[5] = add_71021 == 32'h0000_0005 ? TestBlock__A_op2 : array_index_71020[5];
  assign array_update_71024[6] = add_71021 == 32'h0000_0006 ? TestBlock__A_op2 : array_index_71020[6];
  assign array_update_71024[7] = add_71021 == 32'h0000_0007 ? TestBlock__A_op2 : array_index_71020[7];
  assign array_update_71024[8] = add_71021 == 32'h0000_0008 ? TestBlock__A_op2 : array_index_71020[8];
  assign array_update_71024[9] = add_71021 == 32'h0000_0009 ? TestBlock__A_op2 : array_index_71020[9];
  assign array_update_71025[0] = add_71023 == 32'h0000_0000 ? TestBlock__B_op2 : array_index_71022[0];
  assign array_update_71025[1] = add_71023 == 32'h0000_0001 ? TestBlock__B_op2 : array_index_71022[1];
  assign array_update_71025[2] = add_71023 == 32'h0000_0002 ? TestBlock__B_op2 : array_index_71022[2];
  assign array_update_71025[3] = add_71023 == 32'h0000_0003 ? TestBlock__B_op2 : array_index_71022[3];
  assign array_update_71025[4] = add_71023 == 32'h0000_0004 ? TestBlock__B_op2 : array_index_71022[4];
  assign array_update_71025[5] = add_71023 == 32'h0000_0005 ? TestBlock__B_op2 : array_index_71022[5];
  assign array_update_71025[6] = add_71023 == 32'h0000_0006 ? TestBlock__B_op2 : array_index_71022[6];
  assign array_update_71025[7] = add_71023 == 32'h0000_0007 ? TestBlock__B_op2 : array_index_71022[7];
  assign array_update_71025[8] = add_71023 == 32'h0000_0008 ? TestBlock__B_op2 : array_index_71022[8];
  assign array_update_71025[9] = add_71023 == 32'h0000_0009 ? TestBlock__B_op2 : array_index_71022[9];
  assign array_update_71026[0] = literal_70997 == 32'h0000_0000 ? array_update_71024 : array_update_71016[0];
  assign array_update_71026[1] = literal_70997 == 32'h0000_0001 ? array_update_71024 : array_update_71016[1];
  assign array_update_71026[2] = literal_70997 == 32'h0000_0002 ? array_update_71024 : array_update_71016[2];
  assign array_update_71026[3] = literal_70997 == 32'h0000_0003 ? array_update_71024 : array_update_71016[3];
  assign array_update_71026[4] = literal_70997 == 32'h0000_0004 ? array_update_71024 : array_update_71016[4];
  assign array_update_71026[5] = literal_70997 == 32'h0000_0005 ? array_update_71024 : array_update_71016[5];
  assign array_update_71026[6] = literal_70997 == 32'h0000_0006 ? array_update_71024 : array_update_71016[6];
  assign array_update_71026[7] = literal_70997 == 32'h0000_0007 ? array_update_71024 : array_update_71016[7];
  assign array_update_71026[8] = literal_70997 == 32'h0000_0008 ? array_update_71024 : array_update_71016[8];
  assign array_update_71026[9] = literal_70997 == 32'h0000_0009 ? array_update_71024 : array_update_71016[9];
  assign array_update_71028[0] = literal_70999 == 32'h0000_0000 ? array_update_71025 : array_update_71018[0];
  assign array_update_71028[1] = literal_70999 == 32'h0000_0001 ? array_update_71025 : array_update_71018[1];
  assign array_update_71028[2] = literal_70999 == 32'h0000_0002 ? array_update_71025 : array_update_71018[2];
  assign array_update_71028[3] = literal_70999 == 32'h0000_0003 ? array_update_71025 : array_update_71018[3];
  assign array_update_71028[4] = literal_70999 == 32'h0000_0004 ? array_update_71025 : array_update_71018[4];
  assign array_update_71028[5] = literal_70999 == 32'h0000_0005 ? array_update_71025 : array_update_71018[5];
  assign array_update_71028[6] = literal_70999 == 32'h0000_0006 ? array_update_71025 : array_update_71018[6];
  assign array_update_71028[7] = literal_70999 == 32'h0000_0007 ? array_update_71025 : array_update_71018[7];
  assign array_update_71028[8] = literal_70999 == 32'h0000_0008 ? array_update_71025 : array_update_71018[8];
  assign array_update_71028[9] = literal_70999 == 32'h0000_0009 ? array_update_71025 : array_update_71018[9];
  assign array_index_71030 = array_update_71026[literal_70997 > 32'h0000_0009 ? 4'h9 : literal_70997[3:0]];
  assign add_71031 = add_71021 + 32'h0000_0001;
  assign array_index_71032 = array_update_71028[literal_70999 > 32'h0000_0009 ? 4'h9 : literal_70999[3:0]];
  assign add_71033 = add_71023 + 32'h0000_0001;
  assign array_update_71034[0] = add_71031 == 32'h0000_0000 ? TestBlock__A_op3 : array_index_71030[0];
  assign array_update_71034[1] = add_71031 == 32'h0000_0001 ? TestBlock__A_op3 : array_index_71030[1];
  assign array_update_71034[2] = add_71031 == 32'h0000_0002 ? TestBlock__A_op3 : array_index_71030[2];
  assign array_update_71034[3] = add_71031 == 32'h0000_0003 ? TestBlock__A_op3 : array_index_71030[3];
  assign array_update_71034[4] = add_71031 == 32'h0000_0004 ? TestBlock__A_op3 : array_index_71030[4];
  assign array_update_71034[5] = add_71031 == 32'h0000_0005 ? TestBlock__A_op3 : array_index_71030[5];
  assign array_update_71034[6] = add_71031 == 32'h0000_0006 ? TestBlock__A_op3 : array_index_71030[6];
  assign array_update_71034[7] = add_71031 == 32'h0000_0007 ? TestBlock__A_op3 : array_index_71030[7];
  assign array_update_71034[8] = add_71031 == 32'h0000_0008 ? TestBlock__A_op3 : array_index_71030[8];
  assign array_update_71034[9] = add_71031 == 32'h0000_0009 ? TestBlock__A_op3 : array_index_71030[9];
  assign array_update_71035[0] = add_71033 == 32'h0000_0000 ? TestBlock__B_op3 : array_index_71032[0];
  assign array_update_71035[1] = add_71033 == 32'h0000_0001 ? TestBlock__B_op3 : array_index_71032[1];
  assign array_update_71035[2] = add_71033 == 32'h0000_0002 ? TestBlock__B_op3 : array_index_71032[2];
  assign array_update_71035[3] = add_71033 == 32'h0000_0003 ? TestBlock__B_op3 : array_index_71032[3];
  assign array_update_71035[4] = add_71033 == 32'h0000_0004 ? TestBlock__B_op3 : array_index_71032[4];
  assign array_update_71035[5] = add_71033 == 32'h0000_0005 ? TestBlock__B_op3 : array_index_71032[5];
  assign array_update_71035[6] = add_71033 == 32'h0000_0006 ? TestBlock__B_op3 : array_index_71032[6];
  assign array_update_71035[7] = add_71033 == 32'h0000_0007 ? TestBlock__B_op3 : array_index_71032[7];
  assign array_update_71035[8] = add_71033 == 32'h0000_0008 ? TestBlock__B_op3 : array_index_71032[8];
  assign array_update_71035[9] = add_71033 == 32'h0000_0009 ? TestBlock__B_op3 : array_index_71032[9];
  assign array_update_71036[0] = literal_70997 == 32'h0000_0000 ? array_update_71034 : array_update_71026[0];
  assign array_update_71036[1] = literal_70997 == 32'h0000_0001 ? array_update_71034 : array_update_71026[1];
  assign array_update_71036[2] = literal_70997 == 32'h0000_0002 ? array_update_71034 : array_update_71026[2];
  assign array_update_71036[3] = literal_70997 == 32'h0000_0003 ? array_update_71034 : array_update_71026[3];
  assign array_update_71036[4] = literal_70997 == 32'h0000_0004 ? array_update_71034 : array_update_71026[4];
  assign array_update_71036[5] = literal_70997 == 32'h0000_0005 ? array_update_71034 : array_update_71026[5];
  assign array_update_71036[6] = literal_70997 == 32'h0000_0006 ? array_update_71034 : array_update_71026[6];
  assign array_update_71036[7] = literal_70997 == 32'h0000_0007 ? array_update_71034 : array_update_71026[7];
  assign array_update_71036[8] = literal_70997 == 32'h0000_0008 ? array_update_71034 : array_update_71026[8];
  assign array_update_71036[9] = literal_70997 == 32'h0000_0009 ? array_update_71034 : array_update_71026[9];
  assign array_update_71038[0] = literal_70999 == 32'h0000_0000 ? array_update_71035 : array_update_71028[0];
  assign array_update_71038[1] = literal_70999 == 32'h0000_0001 ? array_update_71035 : array_update_71028[1];
  assign array_update_71038[2] = literal_70999 == 32'h0000_0002 ? array_update_71035 : array_update_71028[2];
  assign array_update_71038[3] = literal_70999 == 32'h0000_0003 ? array_update_71035 : array_update_71028[3];
  assign array_update_71038[4] = literal_70999 == 32'h0000_0004 ? array_update_71035 : array_update_71028[4];
  assign array_update_71038[5] = literal_70999 == 32'h0000_0005 ? array_update_71035 : array_update_71028[5];
  assign array_update_71038[6] = literal_70999 == 32'h0000_0006 ? array_update_71035 : array_update_71028[6];
  assign array_update_71038[7] = literal_70999 == 32'h0000_0007 ? array_update_71035 : array_update_71028[7];
  assign array_update_71038[8] = literal_70999 == 32'h0000_0008 ? array_update_71035 : array_update_71028[8];
  assign array_update_71038[9] = literal_70999 == 32'h0000_0009 ? array_update_71035 : array_update_71028[9];
  assign array_index_71040 = array_update_71036[literal_70997 > 32'h0000_0009 ? 4'h9 : literal_70997[3:0]];
  assign add_71041 = add_71031 + 32'h0000_0001;
  assign array_index_71042 = array_update_71038[literal_70999 > 32'h0000_0009 ? 4'h9 : literal_70999[3:0]];
  assign add_71043 = add_71033 + 32'h0000_0001;
  assign array_update_71044[0] = add_71041 == 32'h0000_0000 ? TestBlock__A_op4 : array_index_71040[0];
  assign array_update_71044[1] = add_71041 == 32'h0000_0001 ? TestBlock__A_op4 : array_index_71040[1];
  assign array_update_71044[2] = add_71041 == 32'h0000_0002 ? TestBlock__A_op4 : array_index_71040[2];
  assign array_update_71044[3] = add_71041 == 32'h0000_0003 ? TestBlock__A_op4 : array_index_71040[3];
  assign array_update_71044[4] = add_71041 == 32'h0000_0004 ? TestBlock__A_op4 : array_index_71040[4];
  assign array_update_71044[5] = add_71041 == 32'h0000_0005 ? TestBlock__A_op4 : array_index_71040[5];
  assign array_update_71044[6] = add_71041 == 32'h0000_0006 ? TestBlock__A_op4 : array_index_71040[6];
  assign array_update_71044[7] = add_71041 == 32'h0000_0007 ? TestBlock__A_op4 : array_index_71040[7];
  assign array_update_71044[8] = add_71041 == 32'h0000_0008 ? TestBlock__A_op4 : array_index_71040[8];
  assign array_update_71044[9] = add_71041 == 32'h0000_0009 ? TestBlock__A_op4 : array_index_71040[9];
  assign array_update_71045[0] = add_71043 == 32'h0000_0000 ? TestBlock__B_op4 : array_index_71042[0];
  assign array_update_71045[1] = add_71043 == 32'h0000_0001 ? TestBlock__B_op4 : array_index_71042[1];
  assign array_update_71045[2] = add_71043 == 32'h0000_0002 ? TestBlock__B_op4 : array_index_71042[2];
  assign array_update_71045[3] = add_71043 == 32'h0000_0003 ? TestBlock__B_op4 : array_index_71042[3];
  assign array_update_71045[4] = add_71043 == 32'h0000_0004 ? TestBlock__B_op4 : array_index_71042[4];
  assign array_update_71045[5] = add_71043 == 32'h0000_0005 ? TestBlock__B_op4 : array_index_71042[5];
  assign array_update_71045[6] = add_71043 == 32'h0000_0006 ? TestBlock__B_op4 : array_index_71042[6];
  assign array_update_71045[7] = add_71043 == 32'h0000_0007 ? TestBlock__B_op4 : array_index_71042[7];
  assign array_update_71045[8] = add_71043 == 32'h0000_0008 ? TestBlock__B_op4 : array_index_71042[8];
  assign array_update_71045[9] = add_71043 == 32'h0000_0009 ? TestBlock__B_op4 : array_index_71042[9];
  assign array_update_71046[0] = literal_70997 == 32'h0000_0000 ? array_update_71044 : array_update_71036[0];
  assign array_update_71046[1] = literal_70997 == 32'h0000_0001 ? array_update_71044 : array_update_71036[1];
  assign array_update_71046[2] = literal_70997 == 32'h0000_0002 ? array_update_71044 : array_update_71036[2];
  assign array_update_71046[3] = literal_70997 == 32'h0000_0003 ? array_update_71044 : array_update_71036[3];
  assign array_update_71046[4] = literal_70997 == 32'h0000_0004 ? array_update_71044 : array_update_71036[4];
  assign array_update_71046[5] = literal_70997 == 32'h0000_0005 ? array_update_71044 : array_update_71036[5];
  assign array_update_71046[6] = literal_70997 == 32'h0000_0006 ? array_update_71044 : array_update_71036[6];
  assign array_update_71046[7] = literal_70997 == 32'h0000_0007 ? array_update_71044 : array_update_71036[7];
  assign array_update_71046[8] = literal_70997 == 32'h0000_0008 ? array_update_71044 : array_update_71036[8];
  assign array_update_71046[9] = literal_70997 == 32'h0000_0009 ? array_update_71044 : array_update_71036[9];
  assign array_update_71048[0] = literal_70999 == 32'h0000_0000 ? array_update_71045 : array_update_71038[0];
  assign array_update_71048[1] = literal_70999 == 32'h0000_0001 ? array_update_71045 : array_update_71038[1];
  assign array_update_71048[2] = literal_70999 == 32'h0000_0002 ? array_update_71045 : array_update_71038[2];
  assign array_update_71048[3] = literal_70999 == 32'h0000_0003 ? array_update_71045 : array_update_71038[3];
  assign array_update_71048[4] = literal_70999 == 32'h0000_0004 ? array_update_71045 : array_update_71038[4];
  assign array_update_71048[5] = literal_70999 == 32'h0000_0005 ? array_update_71045 : array_update_71038[5];
  assign array_update_71048[6] = literal_70999 == 32'h0000_0006 ? array_update_71045 : array_update_71038[6];
  assign array_update_71048[7] = literal_70999 == 32'h0000_0007 ? array_update_71045 : array_update_71038[7];
  assign array_update_71048[8] = literal_70999 == 32'h0000_0008 ? array_update_71045 : array_update_71038[8];
  assign array_update_71048[9] = literal_70999 == 32'h0000_0009 ? array_update_71045 : array_update_71038[9];
  assign array_index_71050 = array_update_71046[literal_70997 > 32'h0000_0009 ? 4'h9 : literal_70997[3:0]];
  assign add_71051 = add_71041 + 32'h0000_0001;
  assign array_index_71052 = array_update_71048[literal_70999 > 32'h0000_0009 ? 4'h9 : literal_70999[3:0]];
  assign add_71053 = add_71043 + 32'h0000_0001;
  assign array_update_71054[0] = add_71051 == 32'h0000_0000 ? TestBlock__A_op5 : array_index_71050[0];
  assign array_update_71054[1] = add_71051 == 32'h0000_0001 ? TestBlock__A_op5 : array_index_71050[1];
  assign array_update_71054[2] = add_71051 == 32'h0000_0002 ? TestBlock__A_op5 : array_index_71050[2];
  assign array_update_71054[3] = add_71051 == 32'h0000_0003 ? TestBlock__A_op5 : array_index_71050[3];
  assign array_update_71054[4] = add_71051 == 32'h0000_0004 ? TestBlock__A_op5 : array_index_71050[4];
  assign array_update_71054[5] = add_71051 == 32'h0000_0005 ? TestBlock__A_op5 : array_index_71050[5];
  assign array_update_71054[6] = add_71051 == 32'h0000_0006 ? TestBlock__A_op5 : array_index_71050[6];
  assign array_update_71054[7] = add_71051 == 32'h0000_0007 ? TestBlock__A_op5 : array_index_71050[7];
  assign array_update_71054[8] = add_71051 == 32'h0000_0008 ? TestBlock__A_op5 : array_index_71050[8];
  assign array_update_71054[9] = add_71051 == 32'h0000_0009 ? TestBlock__A_op5 : array_index_71050[9];
  assign array_update_71055[0] = add_71053 == 32'h0000_0000 ? TestBlock__B_op5 : array_index_71052[0];
  assign array_update_71055[1] = add_71053 == 32'h0000_0001 ? TestBlock__B_op5 : array_index_71052[1];
  assign array_update_71055[2] = add_71053 == 32'h0000_0002 ? TestBlock__B_op5 : array_index_71052[2];
  assign array_update_71055[3] = add_71053 == 32'h0000_0003 ? TestBlock__B_op5 : array_index_71052[3];
  assign array_update_71055[4] = add_71053 == 32'h0000_0004 ? TestBlock__B_op5 : array_index_71052[4];
  assign array_update_71055[5] = add_71053 == 32'h0000_0005 ? TestBlock__B_op5 : array_index_71052[5];
  assign array_update_71055[6] = add_71053 == 32'h0000_0006 ? TestBlock__B_op5 : array_index_71052[6];
  assign array_update_71055[7] = add_71053 == 32'h0000_0007 ? TestBlock__B_op5 : array_index_71052[7];
  assign array_update_71055[8] = add_71053 == 32'h0000_0008 ? TestBlock__B_op5 : array_index_71052[8];
  assign array_update_71055[9] = add_71053 == 32'h0000_0009 ? TestBlock__B_op5 : array_index_71052[9];
  assign array_update_71056[0] = literal_70997 == 32'h0000_0000 ? array_update_71054 : array_update_71046[0];
  assign array_update_71056[1] = literal_70997 == 32'h0000_0001 ? array_update_71054 : array_update_71046[1];
  assign array_update_71056[2] = literal_70997 == 32'h0000_0002 ? array_update_71054 : array_update_71046[2];
  assign array_update_71056[3] = literal_70997 == 32'h0000_0003 ? array_update_71054 : array_update_71046[3];
  assign array_update_71056[4] = literal_70997 == 32'h0000_0004 ? array_update_71054 : array_update_71046[4];
  assign array_update_71056[5] = literal_70997 == 32'h0000_0005 ? array_update_71054 : array_update_71046[5];
  assign array_update_71056[6] = literal_70997 == 32'h0000_0006 ? array_update_71054 : array_update_71046[6];
  assign array_update_71056[7] = literal_70997 == 32'h0000_0007 ? array_update_71054 : array_update_71046[7];
  assign array_update_71056[8] = literal_70997 == 32'h0000_0008 ? array_update_71054 : array_update_71046[8];
  assign array_update_71056[9] = literal_70997 == 32'h0000_0009 ? array_update_71054 : array_update_71046[9];
  assign array_update_71058[0] = literal_70999 == 32'h0000_0000 ? array_update_71055 : array_update_71048[0];
  assign array_update_71058[1] = literal_70999 == 32'h0000_0001 ? array_update_71055 : array_update_71048[1];
  assign array_update_71058[2] = literal_70999 == 32'h0000_0002 ? array_update_71055 : array_update_71048[2];
  assign array_update_71058[3] = literal_70999 == 32'h0000_0003 ? array_update_71055 : array_update_71048[3];
  assign array_update_71058[4] = literal_70999 == 32'h0000_0004 ? array_update_71055 : array_update_71048[4];
  assign array_update_71058[5] = literal_70999 == 32'h0000_0005 ? array_update_71055 : array_update_71048[5];
  assign array_update_71058[6] = literal_70999 == 32'h0000_0006 ? array_update_71055 : array_update_71048[6];
  assign array_update_71058[7] = literal_70999 == 32'h0000_0007 ? array_update_71055 : array_update_71048[7];
  assign array_update_71058[8] = literal_70999 == 32'h0000_0008 ? array_update_71055 : array_update_71048[8];
  assign array_update_71058[9] = literal_70999 == 32'h0000_0009 ? array_update_71055 : array_update_71048[9];
  assign array_index_71060 = array_update_71056[literal_70997 > 32'h0000_0009 ? 4'h9 : literal_70997[3:0]];
  assign add_71061 = add_71051 + 32'h0000_0001;
  assign array_index_71062 = array_update_71058[literal_70999 > 32'h0000_0009 ? 4'h9 : literal_70999[3:0]];
  assign add_71063 = add_71053 + 32'h0000_0001;
  assign array_update_71064[0] = add_71061 == 32'h0000_0000 ? TestBlock__A_op6 : array_index_71060[0];
  assign array_update_71064[1] = add_71061 == 32'h0000_0001 ? TestBlock__A_op6 : array_index_71060[1];
  assign array_update_71064[2] = add_71061 == 32'h0000_0002 ? TestBlock__A_op6 : array_index_71060[2];
  assign array_update_71064[3] = add_71061 == 32'h0000_0003 ? TestBlock__A_op6 : array_index_71060[3];
  assign array_update_71064[4] = add_71061 == 32'h0000_0004 ? TestBlock__A_op6 : array_index_71060[4];
  assign array_update_71064[5] = add_71061 == 32'h0000_0005 ? TestBlock__A_op6 : array_index_71060[5];
  assign array_update_71064[6] = add_71061 == 32'h0000_0006 ? TestBlock__A_op6 : array_index_71060[6];
  assign array_update_71064[7] = add_71061 == 32'h0000_0007 ? TestBlock__A_op6 : array_index_71060[7];
  assign array_update_71064[8] = add_71061 == 32'h0000_0008 ? TestBlock__A_op6 : array_index_71060[8];
  assign array_update_71064[9] = add_71061 == 32'h0000_0009 ? TestBlock__A_op6 : array_index_71060[9];
  assign array_update_71065[0] = add_71063 == 32'h0000_0000 ? TestBlock__B_op6 : array_index_71062[0];
  assign array_update_71065[1] = add_71063 == 32'h0000_0001 ? TestBlock__B_op6 : array_index_71062[1];
  assign array_update_71065[2] = add_71063 == 32'h0000_0002 ? TestBlock__B_op6 : array_index_71062[2];
  assign array_update_71065[3] = add_71063 == 32'h0000_0003 ? TestBlock__B_op6 : array_index_71062[3];
  assign array_update_71065[4] = add_71063 == 32'h0000_0004 ? TestBlock__B_op6 : array_index_71062[4];
  assign array_update_71065[5] = add_71063 == 32'h0000_0005 ? TestBlock__B_op6 : array_index_71062[5];
  assign array_update_71065[6] = add_71063 == 32'h0000_0006 ? TestBlock__B_op6 : array_index_71062[6];
  assign array_update_71065[7] = add_71063 == 32'h0000_0007 ? TestBlock__B_op6 : array_index_71062[7];
  assign array_update_71065[8] = add_71063 == 32'h0000_0008 ? TestBlock__B_op6 : array_index_71062[8];
  assign array_update_71065[9] = add_71063 == 32'h0000_0009 ? TestBlock__B_op6 : array_index_71062[9];
  assign array_update_71066[0] = literal_70997 == 32'h0000_0000 ? array_update_71064 : array_update_71056[0];
  assign array_update_71066[1] = literal_70997 == 32'h0000_0001 ? array_update_71064 : array_update_71056[1];
  assign array_update_71066[2] = literal_70997 == 32'h0000_0002 ? array_update_71064 : array_update_71056[2];
  assign array_update_71066[3] = literal_70997 == 32'h0000_0003 ? array_update_71064 : array_update_71056[3];
  assign array_update_71066[4] = literal_70997 == 32'h0000_0004 ? array_update_71064 : array_update_71056[4];
  assign array_update_71066[5] = literal_70997 == 32'h0000_0005 ? array_update_71064 : array_update_71056[5];
  assign array_update_71066[6] = literal_70997 == 32'h0000_0006 ? array_update_71064 : array_update_71056[6];
  assign array_update_71066[7] = literal_70997 == 32'h0000_0007 ? array_update_71064 : array_update_71056[7];
  assign array_update_71066[8] = literal_70997 == 32'h0000_0008 ? array_update_71064 : array_update_71056[8];
  assign array_update_71066[9] = literal_70997 == 32'h0000_0009 ? array_update_71064 : array_update_71056[9];
  assign array_update_71068[0] = literal_70999 == 32'h0000_0000 ? array_update_71065 : array_update_71058[0];
  assign array_update_71068[1] = literal_70999 == 32'h0000_0001 ? array_update_71065 : array_update_71058[1];
  assign array_update_71068[2] = literal_70999 == 32'h0000_0002 ? array_update_71065 : array_update_71058[2];
  assign array_update_71068[3] = literal_70999 == 32'h0000_0003 ? array_update_71065 : array_update_71058[3];
  assign array_update_71068[4] = literal_70999 == 32'h0000_0004 ? array_update_71065 : array_update_71058[4];
  assign array_update_71068[5] = literal_70999 == 32'h0000_0005 ? array_update_71065 : array_update_71058[5];
  assign array_update_71068[6] = literal_70999 == 32'h0000_0006 ? array_update_71065 : array_update_71058[6];
  assign array_update_71068[7] = literal_70999 == 32'h0000_0007 ? array_update_71065 : array_update_71058[7];
  assign array_update_71068[8] = literal_70999 == 32'h0000_0008 ? array_update_71065 : array_update_71058[8];
  assign array_update_71068[9] = literal_70999 == 32'h0000_0009 ? array_update_71065 : array_update_71058[9];
  assign array_index_71070 = array_update_71066[literal_70997 > 32'h0000_0009 ? 4'h9 : literal_70997[3:0]];
  assign add_71071 = add_71061 + 32'h0000_0001;
  assign array_index_71072 = array_update_71068[literal_70999 > 32'h0000_0009 ? 4'h9 : literal_70999[3:0]];
  assign add_71073 = add_71063 + 32'h0000_0001;
  assign array_update_71074[0] = add_71071 == 32'h0000_0000 ? TestBlock__A_op7 : array_index_71070[0];
  assign array_update_71074[1] = add_71071 == 32'h0000_0001 ? TestBlock__A_op7 : array_index_71070[1];
  assign array_update_71074[2] = add_71071 == 32'h0000_0002 ? TestBlock__A_op7 : array_index_71070[2];
  assign array_update_71074[3] = add_71071 == 32'h0000_0003 ? TestBlock__A_op7 : array_index_71070[3];
  assign array_update_71074[4] = add_71071 == 32'h0000_0004 ? TestBlock__A_op7 : array_index_71070[4];
  assign array_update_71074[5] = add_71071 == 32'h0000_0005 ? TestBlock__A_op7 : array_index_71070[5];
  assign array_update_71074[6] = add_71071 == 32'h0000_0006 ? TestBlock__A_op7 : array_index_71070[6];
  assign array_update_71074[7] = add_71071 == 32'h0000_0007 ? TestBlock__A_op7 : array_index_71070[7];
  assign array_update_71074[8] = add_71071 == 32'h0000_0008 ? TestBlock__A_op7 : array_index_71070[8];
  assign array_update_71074[9] = add_71071 == 32'h0000_0009 ? TestBlock__A_op7 : array_index_71070[9];
  assign array_update_71075[0] = add_71073 == 32'h0000_0000 ? TestBlock__B_op7 : array_index_71072[0];
  assign array_update_71075[1] = add_71073 == 32'h0000_0001 ? TestBlock__B_op7 : array_index_71072[1];
  assign array_update_71075[2] = add_71073 == 32'h0000_0002 ? TestBlock__B_op7 : array_index_71072[2];
  assign array_update_71075[3] = add_71073 == 32'h0000_0003 ? TestBlock__B_op7 : array_index_71072[3];
  assign array_update_71075[4] = add_71073 == 32'h0000_0004 ? TestBlock__B_op7 : array_index_71072[4];
  assign array_update_71075[5] = add_71073 == 32'h0000_0005 ? TestBlock__B_op7 : array_index_71072[5];
  assign array_update_71075[6] = add_71073 == 32'h0000_0006 ? TestBlock__B_op7 : array_index_71072[6];
  assign array_update_71075[7] = add_71073 == 32'h0000_0007 ? TestBlock__B_op7 : array_index_71072[7];
  assign array_update_71075[8] = add_71073 == 32'h0000_0008 ? TestBlock__B_op7 : array_index_71072[8];
  assign array_update_71075[9] = add_71073 == 32'h0000_0009 ? TestBlock__B_op7 : array_index_71072[9];
  assign array_update_71076[0] = literal_70997 == 32'h0000_0000 ? array_update_71074 : array_update_71066[0];
  assign array_update_71076[1] = literal_70997 == 32'h0000_0001 ? array_update_71074 : array_update_71066[1];
  assign array_update_71076[2] = literal_70997 == 32'h0000_0002 ? array_update_71074 : array_update_71066[2];
  assign array_update_71076[3] = literal_70997 == 32'h0000_0003 ? array_update_71074 : array_update_71066[3];
  assign array_update_71076[4] = literal_70997 == 32'h0000_0004 ? array_update_71074 : array_update_71066[4];
  assign array_update_71076[5] = literal_70997 == 32'h0000_0005 ? array_update_71074 : array_update_71066[5];
  assign array_update_71076[6] = literal_70997 == 32'h0000_0006 ? array_update_71074 : array_update_71066[6];
  assign array_update_71076[7] = literal_70997 == 32'h0000_0007 ? array_update_71074 : array_update_71066[7];
  assign array_update_71076[8] = literal_70997 == 32'h0000_0008 ? array_update_71074 : array_update_71066[8];
  assign array_update_71076[9] = literal_70997 == 32'h0000_0009 ? array_update_71074 : array_update_71066[9];
  assign array_update_71078[0] = literal_70999 == 32'h0000_0000 ? array_update_71075 : array_update_71068[0];
  assign array_update_71078[1] = literal_70999 == 32'h0000_0001 ? array_update_71075 : array_update_71068[1];
  assign array_update_71078[2] = literal_70999 == 32'h0000_0002 ? array_update_71075 : array_update_71068[2];
  assign array_update_71078[3] = literal_70999 == 32'h0000_0003 ? array_update_71075 : array_update_71068[3];
  assign array_update_71078[4] = literal_70999 == 32'h0000_0004 ? array_update_71075 : array_update_71068[4];
  assign array_update_71078[5] = literal_70999 == 32'h0000_0005 ? array_update_71075 : array_update_71068[5];
  assign array_update_71078[6] = literal_70999 == 32'h0000_0006 ? array_update_71075 : array_update_71068[6];
  assign array_update_71078[7] = literal_70999 == 32'h0000_0007 ? array_update_71075 : array_update_71068[7];
  assign array_update_71078[8] = literal_70999 == 32'h0000_0008 ? array_update_71075 : array_update_71068[8];
  assign array_update_71078[9] = literal_70999 == 32'h0000_0009 ? array_update_71075 : array_update_71068[9];
  assign array_index_71080 = array_update_71076[literal_70997 > 32'h0000_0009 ? 4'h9 : literal_70997[3:0]];
  assign add_71081 = add_71071 + 32'h0000_0001;
  assign array_index_71082 = array_update_71078[literal_70999 > 32'h0000_0009 ? 4'h9 : literal_70999[3:0]];
  assign add_71083 = add_71073 + 32'h0000_0001;
  assign array_update_71084[0] = add_71081 == 32'h0000_0000 ? TestBlock__A_op8 : array_index_71080[0];
  assign array_update_71084[1] = add_71081 == 32'h0000_0001 ? TestBlock__A_op8 : array_index_71080[1];
  assign array_update_71084[2] = add_71081 == 32'h0000_0002 ? TestBlock__A_op8 : array_index_71080[2];
  assign array_update_71084[3] = add_71081 == 32'h0000_0003 ? TestBlock__A_op8 : array_index_71080[3];
  assign array_update_71084[4] = add_71081 == 32'h0000_0004 ? TestBlock__A_op8 : array_index_71080[4];
  assign array_update_71084[5] = add_71081 == 32'h0000_0005 ? TestBlock__A_op8 : array_index_71080[5];
  assign array_update_71084[6] = add_71081 == 32'h0000_0006 ? TestBlock__A_op8 : array_index_71080[6];
  assign array_update_71084[7] = add_71081 == 32'h0000_0007 ? TestBlock__A_op8 : array_index_71080[7];
  assign array_update_71084[8] = add_71081 == 32'h0000_0008 ? TestBlock__A_op8 : array_index_71080[8];
  assign array_update_71084[9] = add_71081 == 32'h0000_0009 ? TestBlock__A_op8 : array_index_71080[9];
  assign array_update_71085[0] = add_71083 == 32'h0000_0000 ? TestBlock__B_op8 : array_index_71082[0];
  assign array_update_71085[1] = add_71083 == 32'h0000_0001 ? TestBlock__B_op8 : array_index_71082[1];
  assign array_update_71085[2] = add_71083 == 32'h0000_0002 ? TestBlock__B_op8 : array_index_71082[2];
  assign array_update_71085[3] = add_71083 == 32'h0000_0003 ? TestBlock__B_op8 : array_index_71082[3];
  assign array_update_71085[4] = add_71083 == 32'h0000_0004 ? TestBlock__B_op8 : array_index_71082[4];
  assign array_update_71085[5] = add_71083 == 32'h0000_0005 ? TestBlock__B_op8 : array_index_71082[5];
  assign array_update_71085[6] = add_71083 == 32'h0000_0006 ? TestBlock__B_op8 : array_index_71082[6];
  assign array_update_71085[7] = add_71083 == 32'h0000_0007 ? TestBlock__B_op8 : array_index_71082[7];
  assign array_update_71085[8] = add_71083 == 32'h0000_0008 ? TestBlock__B_op8 : array_index_71082[8];
  assign array_update_71085[9] = add_71083 == 32'h0000_0009 ? TestBlock__B_op8 : array_index_71082[9];
  assign array_update_71086[0] = literal_70997 == 32'h0000_0000 ? array_update_71084 : array_update_71076[0];
  assign array_update_71086[1] = literal_70997 == 32'h0000_0001 ? array_update_71084 : array_update_71076[1];
  assign array_update_71086[2] = literal_70997 == 32'h0000_0002 ? array_update_71084 : array_update_71076[2];
  assign array_update_71086[3] = literal_70997 == 32'h0000_0003 ? array_update_71084 : array_update_71076[3];
  assign array_update_71086[4] = literal_70997 == 32'h0000_0004 ? array_update_71084 : array_update_71076[4];
  assign array_update_71086[5] = literal_70997 == 32'h0000_0005 ? array_update_71084 : array_update_71076[5];
  assign array_update_71086[6] = literal_70997 == 32'h0000_0006 ? array_update_71084 : array_update_71076[6];
  assign array_update_71086[7] = literal_70997 == 32'h0000_0007 ? array_update_71084 : array_update_71076[7];
  assign array_update_71086[8] = literal_70997 == 32'h0000_0008 ? array_update_71084 : array_update_71076[8];
  assign array_update_71086[9] = literal_70997 == 32'h0000_0009 ? array_update_71084 : array_update_71076[9];
  assign array_update_71088[0] = literal_70999 == 32'h0000_0000 ? array_update_71085 : array_update_71078[0];
  assign array_update_71088[1] = literal_70999 == 32'h0000_0001 ? array_update_71085 : array_update_71078[1];
  assign array_update_71088[2] = literal_70999 == 32'h0000_0002 ? array_update_71085 : array_update_71078[2];
  assign array_update_71088[3] = literal_70999 == 32'h0000_0003 ? array_update_71085 : array_update_71078[3];
  assign array_update_71088[4] = literal_70999 == 32'h0000_0004 ? array_update_71085 : array_update_71078[4];
  assign array_update_71088[5] = literal_70999 == 32'h0000_0005 ? array_update_71085 : array_update_71078[5];
  assign array_update_71088[6] = literal_70999 == 32'h0000_0006 ? array_update_71085 : array_update_71078[6];
  assign array_update_71088[7] = literal_70999 == 32'h0000_0007 ? array_update_71085 : array_update_71078[7];
  assign array_update_71088[8] = literal_70999 == 32'h0000_0008 ? array_update_71085 : array_update_71078[8];
  assign array_update_71088[9] = literal_70999 == 32'h0000_0009 ? array_update_71085 : array_update_71078[9];
  assign array_index_71090 = array_update_71086[literal_70997 > 32'h0000_0009 ? 4'h9 : literal_70997[3:0]];
  assign add_71091 = add_71081 + 32'h0000_0001;
  assign array_index_71092 = array_update_71088[literal_70999 > 32'h0000_0009 ? 4'h9 : literal_70999[3:0]];
  assign add_71093 = add_71083 + 32'h0000_0001;
  assign array_update_71094[0] = add_71091 == 32'h0000_0000 ? TestBlock__A_op9 : array_index_71090[0];
  assign array_update_71094[1] = add_71091 == 32'h0000_0001 ? TestBlock__A_op9 : array_index_71090[1];
  assign array_update_71094[2] = add_71091 == 32'h0000_0002 ? TestBlock__A_op9 : array_index_71090[2];
  assign array_update_71094[3] = add_71091 == 32'h0000_0003 ? TestBlock__A_op9 : array_index_71090[3];
  assign array_update_71094[4] = add_71091 == 32'h0000_0004 ? TestBlock__A_op9 : array_index_71090[4];
  assign array_update_71094[5] = add_71091 == 32'h0000_0005 ? TestBlock__A_op9 : array_index_71090[5];
  assign array_update_71094[6] = add_71091 == 32'h0000_0006 ? TestBlock__A_op9 : array_index_71090[6];
  assign array_update_71094[7] = add_71091 == 32'h0000_0007 ? TestBlock__A_op9 : array_index_71090[7];
  assign array_update_71094[8] = add_71091 == 32'h0000_0008 ? TestBlock__A_op9 : array_index_71090[8];
  assign array_update_71094[9] = add_71091 == 32'h0000_0009 ? TestBlock__A_op9 : array_index_71090[9];
  assign array_update_71096[0] = add_71093 == 32'h0000_0000 ? TestBlock__B_op9 : array_index_71092[0];
  assign array_update_71096[1] = add_71093 == 32'h0000_0001 ? TestBlock__B_op9 : array_index_71092[1];
  assign array_update_71096[2] = add_71093 == 32'h0000_0002 ? TestBlock__B_op9 : array_index_71092[2];
  assign array_update_71096[3] = add_71093 == 32'h0000_0003 ? TestBlock__B_op9 : array_index_71092[3];
  assign array_update_71096[4] = add_71093 == 32'h0000_0004 ? TestBlock__B_op9 : array_index_71092[4];
  assign array_update_71096[5] = add_71093 == 32'h0000_0005 ? TestBlock__B_op9 : array_index_71092[5];
  assign array_update_71096[6] = add_71093 == 32'h0000_0006 ? TestBlock__B_op9 : array_index_71092[6];
  assign array_update_71096[7] = add_71093 == 32'h0000_0007 ? TestBlock__B_op9 : array_index_71092[7];
  assign array_update_71096[8] = add_71093 == 32'h0000_0008 ? TestBlock__B_op9 : array_index_71092[8];
  assign array_update_71096[9] = add_71093 == 32'h0000_0009 ? TestBlock__B_op9 : array_index_71092[9];
  assign array_update_71098[0] = literal_70997 == 32'h0000_0000 ? array_update_71094 : array_update_71086[0];
  assign array_update_71098[1] = literal_70997 == 32'h0000_0001 ? array_update_71094 : array_update_71086[1];
  assign array_update_71098[2] = literal_70997 == 32'h0000_0002 ? array_update_71094 : array_update_71086[2];
  assign array_update_71098[3] = literal_70997 == 32'h0000_0003 ? array_update_71094 : array_update_71086[3];
  assign array_update_71098[4] = literal_70997 == 32'h0000_0004 ? array_update_71094 : array_update_71086[4];
  assign array_update_71098[5] = literal_70997 == 32'h0000_0005 ? array_update_71094 : array_update_71086[5];
  assign array_update_71098[6] = literal_70997 == 32'h0000_0006 ? array_update_71094 : array_update_71086[6];
  assign array_update_71098[7] = literal_70997 == 32'h0000_0007 ? array_update_71094 : array_update_71086[7];
  assign array_update_71098[8] = literal_70997 == 32'h0000_0008 ? array_update_71094 : array_update_71086[8];
  assign array_update_71098[9] = literal_70997 == 32'h0000_0009 ? array_update_71094 : array_update_71086[9];
  assign add_71099 = literal_70997 + 32'h0000_0001;
  assign array_update_71100[0] = literal_70999 == 32'h0000_0000 ? array_update_71096 : array_update_71088[0];
  assign array_update_71100[1] = literal_70999 == 32'h0000_0001 ? array_update_71096 : array_update_71088[1];
  assign array_update_71100[2] = literal_70999 == 32'h0000_0002 ? array_update_71096 : array_update_71088[2];
  assign array_update_71100[3] = literal_70999 == 32'h0000_0003 ? array_update_71096 : array_update_71088[3];
  assign array_update_71100[4] = literal_70999 == 32'h0000_0004 ? array_update_71096 : array_update_71088[4];
  assign array_update_71100[5] = literal_70999 == 32'h0000_0005 ? array_update_71096 : array_update_71088[5];
  assign array_update_71100[6] = literal_70999 == 32'h0000_0006 ? array_update_71096 : array_update_71088[6];
  assign array_update_71100[7] = literal_70999 == 32'h0000_0007 ? array_update_71096 : array_update_71088[7];
  assign array_update_71100[8] = literal_70999 == 32'h0000_0008 ? array_update_71096 : array_update_71088[8];
  assign array_update_71100[9] = literal_70999 == 32'h0000_0009 ? array_update_71096 : array_update_71088[9];
  assign add_71101 = literal_70999 + 32'h0000_0001;
  assign array_index_71102 = array_update_71098[add_71099 > 32'h0000_0009 ? 4'h9 : add_71099[3:0]];
  assign literal_71103 = 32'h0000_0000;
  assign array_index_71104 = array_update_71100[add_71101 > 32'h0000_0009 ? 4'h9 : add_71101[3:0]];
  assign literal_71105 = 32'h0000_0000;
  assign array_update_71106[0] = literal_71103 == 32'h0000_0000 ? TestBlock__A_op10 : array_index_71102[0];
  assign array_update_71106[1] = literal_71103 == 32'h0000_0001 ? TestBlock__A_op10 : array_index_71102[1];
  assign array_update_71106[2] = literal_71103 == 32'h0000_0002 ? TestBlock__A_op10 : array_index_71102[2];
  assign array_update_71106[3] = literal_71103 == 32'h0000_0003 ? TestBlock__A_op10 : array_index_71102[3];
  assign array_update_71106[4] = literal_71103 == 32'h0000_0004 ? TestBlock__A_op10 : array_index_71102[4];
  assign array_update_71106[5] = literal_71103 == 32'h0000_0005 ? TestBlock__A_op10 : array_index_71102[5];
  assign array_update_71106[6] = literal_71103 == 32'h0000_0006 ? TestBlock__A_op10 : array_index_71102[6];
  assign array_update_71106[7] = literal_71103 == 32'h0000_0007 ? TestBlock__A_op10 : array_index_71102[7];
  assign array_update_71106[8] = literal_71103 == 32'h0000_0008 ? TestBlock__A_op10 : array_index_71102[8];
  assign array_update_71106[9] = literal_71103 == 32'h0000_0009 ? TestBlock__A_op10 : array_index_71102[9];
  assign array_update_71107[0] = literal_71105 == 32'h0000_0000 ? TestBlock__B_op10 : array_index_71104[0];
  assign array_update_71107[1] = literal_71105 == 32'h0000_0001 ? TestBlock__B_op10 : array_index_71104[1];
  assign array_update_71107[2] = literal_71105 == 32'h0000_0002 ? TestBlock__B_op10 : array_index_71104[2];
  assign array_update_71107[3] = literal_71105 == 32'h0000_0003 ? TestBlock__B_op10 : array_index_71104[3];
  assign array_update_71107[4] = literal_71105 == 32'h0000_0004 ? TestBlock__B_op10 : array_index_71104[4];
  assign array_update_71107[5] = literal_71105 == 32'h0000_0005 ? TestBlock__B_op10 : array_index_71104[5];
  assign array_update_71107[6] = literal_71105 == 32'h0000_0006 ? TestBlock__B_op10 : array_index_71104[6];
  assign array_update_71107[7] = literal_71105 == 32'h0000_0007 ? TestBlock__B_op10 : array_index_71104[7];
  assign array_update_71107[8] = literal_71105 == 32'h0000_0008 ? TestBlock__B_op10 : array_index_71104[8];
  assign array_update_71107[9] = literal_71105 == 32'h0000_0009 ? TestBlock__B_op10 : array_index_71104[9];
  assign array_update_71108[0] = add_71099 == 32'h0000_0000 ? array_update_71106 : array_update_71098[0];
  assign array_update_71108[1] = add_71099 == 32'h0000_0001 ? array_update_71106 : array_update_71098[1];
  assign array_update_71108[2] = add_71099 == 32'h0000_0002 ? array_update_71106 : array_update_71098[2];
  assign array_update_71108[3] = add_71099 == 32'h0000_0003 ? array_update_71106 : array_update_71098[3];
  assign array_update_71108[4] = add_71099 == 32'h0000_0004 ? array_update_71106 : array_update_71098[4];
  assign array_update_71108[5] = add_71099 == 32'h0000_0005 ? array_update_71106 : array_update_71098[5];
  assign array_update_71108[6] = add_71099 == 32'h0000_0006 ? array_update_71106 : array_update_71098[6];
  assign array_update_71108[7] = add_71099 == 32'h0000_0007 ? array_update_71106 : array_update_71098[7];
  assign array_update_71108[8] = add_71099 == 32'h0000_0008 ? array_update_71106 : array_update_71098[8];
  assign array_update_71108[9] = add_71099 == 32'h0000_0009 ? array_update_71106 : array_update_71098[9];
  assign array_update_71110[0] = add_71101 == 32'h0000_0000 ? array_update_71107 : array_update_71100[0];
  assign array_update_71110[1] = add_71101 == 32'h0000_0001 ? array_update_71107 : array_update_71100[1];
  assign array_update_71110[2] = add_71101 == 32'h0000_0002 ? array_update_71107 : array_update_71100[2];
  assign array_update_71110[3] = add_71101 == 32'h0000_0003 ? array_update_71107 : array_update_71100[3];
  assign array_update_71110[4] = add_71101 == 32'h0000_0004 ? array_update_71107 : array_update_71100[4];
  assign array_update_71110[5] = add_71101 == 32'h0000_0005 ? array_update_71107 : array_update_71100[5];
  assign array_update_71110[6] = add_71101 == 32'h0000_0006 ? array_update_71107 : array_update_71100[6];
  assign array_update_71110[7] = add_71101 == 32'h0000_0007 ? array_update_71107 : array_update_71100[7];
  assign array_update_71110[8] = add_71101 == 32'h0000_0008 ? array_update_71107 : array_update_71100[8];
  assign array_update_71110[9] = add_71101 == 32'h0000_0009 ? array_update_71107 : array_update_71100[9];
  assign array_index_71112 = array_update_71108[add_71099 > 32'h0000_0009 ? 4'h9 : add_71099[3:0]];
  assign add_71113 = literal_71103 + 32'h0000_0001;
  assign array_index_71114 = array_update_71110[add_71101 > 32'h0000_0009 ? 4'h9 : add_71101[3:0]];
  assign add_71115 = literal_71105 + 32'h0000_0001;
  assign array_update_71116[0] = add_71113 == 32'h0000_0000 ? TestBlock__A_op11 : array_index_71112[0];
  assign array_update_71116[1] = add_71113 == 32'h0000_0001 ? TestBlock__A_op11 : array_index_71112[1];
  assign array_update_71116[2] = add_71113 == 32'h0000_0002 ? TestBlock__A_op11 : array_index_71112[2];
  assign array_update_71116[3] = add_71113 == 32'h0000_0003 ? TestBlock__A_op11 : array_index_71112[3];
  assign array_update_71116[4] = add_71113 == 32'h0000_0004 ? TestBlock__A_op11 : array_index_71112[4];
  assign array_update_71116[5] = add_71113 == 32'h0000_0005 ? TestBlock__A_op11 : array_index_71112[5];
  assign array_update_71116[6] = add_71113 == 32'h0000_0006 ? TestBlock__A_op11 : array_index_71112[6];
  assign array_update_71116[7] = add_71113 == 32'h0000_0007 ? TestBlock__A_op11 : array_index_71112[7];
  assign array_update_71116[8] = add_71113 == 32'h0000_0008 ? TestBlock__A_op11 : array_index_71112[8];
  assign array_update_71116[9] = add_71113 == 32'h0000_0009 ? TestBlock__A_op11 : array_index_71112[9];
  assign array_update_71117[0] = add_71115 == 32'h0000_0000 ? TestBlock__B_op11 : array_index_71114[0];
  assign array_update_71117[1] = add_71115 == 32'h0000_0001 ? TestBlock__B_op11 : array_index_71114[1];
  assign array_update_71117[2] = add_71115 == 32'h0000_0002 ? TestBlock__B_op11 : array_index_71114[2];
  assign array_update_71117[3] = add_71115 == 32'h0000_0003 ? TestBlock__B_op11 : array_index_71114[3];
  assign array_update_71117[4] = add_71115 == 32'h0000_0004 ? TestBlock__B_op11 : array_index_71114[4];
  assign array_update_71117[5] = add_71115 == 32'h0000_0005 ? TestBlock__B_op11 : array_index_71114[5];
  assign array_update_71117[6] = add_71115 == 32'h0000_0006 ? TestBlock__B_op11 : array_index_71114[6];
  assign array_update_71117[7] = add_71115 == 32'h0000_0007 ? TestBlock__B_op11 : array_index_71114[7];
  assign array_update_71117[8] = add_71115 == 32'h0000_0008 ? TestBlock__B_op11 : array_index_71114[8];
  assign array_update_71117[9] = add_71115 == 32'h0000_0009 ? TestBlock__B_op11 : array_index_71114[9];
  assign array_update_71118[0] = add_71099 == 32'h0000_0000 ? array_update_71116 : array_update_71108[0];
  assign array_update_71118[1] = add_71099 == 32'h0000_0001 ? array_update_71116 : array_update_71108[1];
  assign array_update_71118[2] = add_71099 == 32'h0000_0002 ? array_update_71116 : array_update_71108[2];
  assign array_update_71118[3] = add_71099 == 32'h0000_0003 ? array_update_71116 : array_update_71108[3];
  assign array_update_71118[4] = add_71099 == 32'h0000_0004 ? array_update_71116 : array_update_71108[4];
  assign array_update_71118[5] = add_71099 == 32'h0000_0005 ? array_update_71116 : array_update_71108[5];
  assign array_update_71118[6] = add_71099 == 32'h0000_0006 ? array_update_71116 : array_update_71108[6];
  assign array_update_71118[7] = add_71099 == 32'h0000_0007 ? array_update_71116 : array_update_71108[7];
  assign array_update_71118[8] = add_71099 == 32'h0000_0008 ? array_update_71116 : array_update_71108[8];
  assign array_update_71118[9] = add_71099 == 32'h0000_0009 ? array_update_71116 : array_update_71108[9];
  assign array_update_71120[0] = add_71101 == 32'h0000_0000 ? array_update_71117 : array_update_71110[0];
  assign array_update_71120[1] = add_71101 == 32'h0000_0001 ? array_update_71117 : array_update_71110[1];
  assign array_update_71120[2] = add_71101 == 32'h0000_0002 ? array_update_71117 : array_update_71110[2];
  assign array_update_71120[3] = add_71101 == 32'h0000_0003 ? array_update_71117 : array_update_71110[3];
  assign array_update_71120[4] = add_71101 == 32'h0000_0004 ? array_update_71117 : array_update_71110[4];
  assign array_update_71120[5] = add_71101 == 32'h0000_0005 ? array_update_71117 : array_update_71110[5];
  assign array_update_71120[6] = add_71101 == 32'h0000_0006 ? array_update_71117 : array_update_71110[6];
  assign array_update_71120[7] = add_71101 == 32'h0000_0007 ? array_update_71117 : array_update_71110[7];
  assign array_update_71120[8] = add_71101 == 32'h0000_0008 ? array_update_71117 : array_update_71110[8];
  assign array_update_71120[9] = add_71101 == 32'h0000_0009 ? array_update_71117 : array_update_71110[9];
  assign array_index_71122 = array_update_71118[add_71099 > 32'h0000_0009 ? 4'h9 : add_71099[3:0]];
  assign add_71123 = add_71113 + 32'h0000_0001;
  assign array_index_71124 = array_update_71120[add_71101 > 32'h0000_0009 ? 4'h9 : add_71101[3:0]];
  assign add_71125 = add_71115 + 32'h0000_0001;
  assign array_update_71126[0] = add_71123 == 32'h0000_0000 ? TestBlock__A_op12 : array_index_71122[0];
  assign array_update_71126[1] = add_71123 == 32'h0000_0001 ? TestBlock__A_op12 : array_index_71122[1];
  assign array_update_71126[2] = add_71123 == 32'h0000_0002 ? TestBlock__A_op12 : array_index_71122[2];
  assign array_update_71126[3] = add_71123 == 32'h0000_0003 ? TestBlock__A_op12 : array_index_71122[3];
  assign array_update_71126[4] = add_71123 == 32'h0000_0004 ? TestBlock__A_op12 : array_index_71122[4];
  assign array_update_71126[5] = add_71123 == 32'h0000_0005 ? TestBlock__A_op12 : array_index_71122[5];
  assign array_update_71126[6] = add_71123 == 32'h0000_0006 ? TestBlock__A_op12 : array_index_71122[6];
  assign array_update_71126[7] = add_71123 == 32'h0000_0007 ? TestBlock__A_op12 : array_index_71122[7];
  assign array_update_71126[8] = add_71123 == 32'h0000_0008 ? TestBlock__A_op12 : array_index_71122[8];
  assign array_update_71126[9] = add_71123 == 32'h0000_0009 ? TestBlock__A_op12 : array_index_71122[9];
  assign array_update_71127[0] = add_71125 == 32'h0000_0000 ? TestBlock__B_op12 : array_index_71124[0];
  assign array_update_71127[1] = add_71125 == 32'h0000_0001 ? TestBlock__B_op12 : array_index_71124[1];
  assign array_update_71127[2] = add_71125 == 32'h0000_0002 ? TestBlock__B_op12 : array_index_71124[2];
  assign array_update_71127[3] = add_71125 == 32'h0000_0003 ? TestBlock__B_op12 : array_index_71124[3];
  assign array_update_71127[4] = add_71125 == 32'h0000_0004 ? TestBlock__B_op12 : array_index_71124[4];
  assign array_update_71127[5] = add_71125 == 32'h0000_0005 ? TestBlock__B_op12 : array_index_71124[5];
  assign array_update_71127[6] = add_71125 == 32'h0000_0006 ? TestBlock__B_op12 : array_index_71124[6];
  assign array_update_71127[7] = add_71125 == 32'h0000_0007 ? TestBlock__B_op12 : array_index_71124[7];
  assign array_update_71127[8] = add_71125 == 32'h0000_0008 ? TestBlock__B_op12 : array_index_71124[8];
  assign array_update_71127[9] = add_71125 == 32'h0000_0009 ? TestBlock__B_op12 : array_index_71124[9];
  assign array_update_71128[0] = add_71099 == 32'h0000_0000 ? array_update_71126 : array_update_71118[0];
  assign array_update_71128[1] = add_71099 == 32'h0000_0001 ? array_update_71126 : array_update_71118[1];
  assign array_update_71128[2] = add_71099 == 32'h0000_0002 ? array_update_71126 : array_update_71118[2];
  assign array_update_71128[3] = add_71099 == 32'h0000_0003 ? array_update_71126 : array_update_71118[3];
  assign array_update_71128[4] = add_71099 == 32'h0000_0004 ? array_update_71126 : array_update_71118[4];
  assign array_update_71128[5] = add_71099 == 32'h0000_0005 ? array_update_71126 : array_update_71118[5];
  assign array_update_71128[6] = add_71099 == 32'h0000_0006 ? array_update_71126 : array_update_71118[6];
  assign array_update_71128[7] = add_71099 == 32'h0000_0007 ? array_update_71126 : array_update_71118[7];
  assign array_update_71128[8] = add_71099 == 32'h0000_0008 ? array_update_71126 : array_update_71118[8];
  assign array_update_71128[9] = add_71099 == 32'h0000_0009 ? array_update_71126 : array_update_71118[9];
  assign array_update_71130[0] = add_71101 == 32'h0000_0000 ? array_update_71127 : array_update_71120[0];
  assign array_update_71130[1] = add_71101 == 32'h0000_0001 ? array_update_71127 : array_update_71120[1];
  assign array_update_71130[2] = add_71101 == 32'h0000_0002 ? array_update_71127 : array_update_71120[2];
  assign array_update_71130[3] = add_71101 == 32'h0000_0003 ? array_update_71127 : array_update_71120[3];
  assign array_update_71130[4] = add_71101 == 32'h0000_0004 ? array_update_71127 : array_update_71120[4];
  assign array_update_71130[5] = add_71101 == 32'h0000_0005 ? array_update_71127 : array_update_71120[5];
  assign array_update_71130[6] = add_71101 == 32'h0000_0006 ? array_update_71127 : array_update_71120[6];
  assign array_update_71130[7] = add_71101 == 32'h0000_0007 ? array_update_71127 : array_update_71120[7];
  assign array_update_71130[8] = add_71101 == 32'h0000_0008 ? array_update_71127 : array_update_71120[8];
  assign array_update_71130[9] = add_71101 == 32'h0000_0009 ? array_update_71127 : array_update_71120[9];
  assign array_index_71132 = array_update_71128[add_71099 > 32'h0000_0009 ? 4'h9 : add_71099[3:0]];
  assign add_71133 = add_71123 + 32'h0000_0001;
  assign array_index_71134 = array_update_71130[add_71101 > 32'h0000_0009 ? 4'h9 : add_71101[3:0]];
  assign add_71135 = add_71125 + 32'h0000_0001;
  assign array_update_71136[0] = add_71133 == 32'h0000_0000 ? TestBlock__A_op13 : array_index_71132[0];
  assign array_update_71136[1] = add_71133 == 32'h0000_0001 ? TestBlock__A_op13 : array_index_71132[1];
  assign array_update_71136[2] = add_71133 == 32'h0000_0002 ? TestBlock__A_op13 : array_index_71132[2];
  assign array_update_71136[3] = add_71133 == 32'h0000_0003 ? TestBlock__A_op13 : array_index_71132[3];
  assign array_update_71136[4] = add_71133 == 32'h0000_0004 ? TestBlock__A_op13 : array_index_71132[4];
  assign array_update_71136[5] = add_71133 == 32'h0000_0005 ? TestBlock__A_op13 : array_index_71132[5];
  assign array_update_71136[6] = add_71133 == 32'h0000_0006 ? TestBlock__A_op13 : array_index_71132[6];
  assign array_update_71136[7] = add_71133 == 32'h0000_0007 ? TestBlock__A_op13 : array_index_71132[7];
  assign array_update_71136[8] = add_71133 == 32'h0000_0008 ? TestBlock__A_op13 : array_index_71132[8];
  assign array_update_71136[9] = add_71133 == 32'h0000_0009 ? TestBlock__A_op13 : array_index_71132[9];
  assign array_update_71137[0] = add_71135 == 32'h0000_0000 ? TestBlock__B_op13 : array_index_71134[0];
  assign array_update_71137[1] = add_71135 == 32'h0000_0001 ? TestBlock__B_op13 : array_index_71134[1];
  assign array_update_71137[2] = add_71135 == 32'h0000_0002 ? TestBlock__B_op13 : array_index_71134[2];
  assign array_update_71137[3] = add_71135 == 32'h0000_0003 ? TestBlock__B_op13 : array_index_71134[3];
  assign array_update_71137[4] = add_71135 == 32'h0000_0004 ? TestBlock__B_op13 : array_index_71134[4];
  assign array_update_71137[5] = add_71135 == 32'h0000_0005 ? TestBlock__B_op13 : array_index_71134[5];
  assign array_update_71137[6] = add_71135 == 32'h0000_0006 ? TestBlock__B_op13 : array_index_71134[6];
  assign array_update_71137[7] = add_71135 == 32'h0000_0007 ? TestBlock__B_op13 : array_index_71134[7];
  assign array_update_71137[8] = add_71135 == 32'h0000_0008 ? TestBlock__B_op13 : array_index_71134[8];
  assign array_update_71137[9] = add_71135 == 32'h0000_0009 ? TestBlock__B_op13 : array_index_71134[9];
  assign array_update_71138[0] = add_71099 == 32'h0000_0000 ? array_update_71136 : array_update_71128[0];
  assign array_update_71138[1] = add_71099 == 32'h0000_0001 ? array_update_71136 : array_update_71128[1];
  assign array_update_71138[2] = add_71099 == 32'h0000_0002 ? array_update_71136 : array_update_71128[2];
  assign array_update_71138[3] = add_71099 == 32'h0000_0003 ? array_update_71136 : array_update_71128[3];
  assign array_update_71138[4] = add_71099 == 32'h0000_0004 ? array_update_71136 : array_update_71128[4];
  assign array_update_71138[5] = add_71099 == 32'h0000_0005 ? array_update_71136 : array_update_71128[5];
  assign array_update_71138[6] = add_71099 == 32'h0000_0006 ? array_update_71136 : array_update_71128[6];
  assign array_update_71138[7] = add_71099 == 32'h0000_0007 ? array_update_71136 : array_update_71128[7];
  assign array_update_71138[8] = add_71099 == 32'h0000_0008 ? array_update_71136 : array_update_71128[8];
  assign array_update_71138[9] = add_71099 == 32'h0000_0009 ? array_update_71136 : array_update_71128[9];
  assign array_update_71140[0] = add_71101 == 32'h0000_0000 ? array_update_71137 : array_update_71130[0];
  assign array_update_71140[1] = add_71101 == 32'h0000_0001 ? array_update_71137 : array_update_71130[1];
  assign array_update_71140[2] = add_71101 == 32'h0000_0002 ? array_update_71137 : array_update_71130[2];
  assign array_update_71140[3] = add_71101 == 32'h0000_0003 ? array_update_71137 : array_update_71130[3];
  assign array_update_71140[4] = add_71101 == 32'h0000_0004 ? array_update_71137 : array_update_71130[4];
  assign array_update_71140[5] = add_71101 == 32'h0000_0005 ? array_update_71137 : array_update_71130[5];
  assign array_update_71140[6] = add_71101 == 32'h0000_0006 ? array_update_71137 : array_update_71130[6];
  assign array_update_71140[7] = add_71101 == 32'h0000_0007 ? array_update_71137 : array_update_71130[7];
  assign array_update_71140[8] = add_71101 == 32'h0000_0008 ? array_update_71137 : array_update_71130[8];
  assign array_update_71140[9] = add_71101 == 32'h0000_0009 ? array_update_71137 : array_update_71130[9];
  assign array_index_71142 = array_update_71138[add_71099 > 32'h0000_0009 ? 4'h9 : add_71099[3:0]];
  assign add_71143 = add_71133 + 32'h0000_0001;
  assign array_index_71144 = array_update_71140[add_71101 > 32'h0000_0009 ? 4'h9 : add_71101[3:0]];
  assign add_71145 = add_71135 + 32'h0000_0001;
  assign array_update_71146[0] = add_71143 == 32'h0000_0000 ? TestBlock__A_op14 : array_index_71142[0];
  assign array_update_71146[1] = add_71143 == 32'h0000_0001 ? TestBlock__A_op14 : array_index_71142[1];
  assign array_update_71146[2] = add_71143 == 32'h0000_0002 ? TestBlock__A_op14 : array_index_71142[2];
  assign array_update_71146[3] = add_71143 == 32'h0000_0003 ? TestBlock__A_op14 : array_index_71142[3];
  assign array_update_71146[4] = add_71143 == 32'h0000_0004 ? TestBlock__A_op14 : array_index_71142[4];
  assign array_update_71146[5] = add_71143 == 32'h0000_0005 ? TestBlock__A_op14 : array_index_71142[5];
  assign array_update_71146[6] = add_71143 == 32'h0000_0006 ? TestBlock__A_op14 : array_index_71142[6];
  assign array_update_71146[7] = add_71143 == 32'h0000_0007 ? TestBlock__A_op14 : array_index_71142[7];
  assign array_update_71146[8] = add_71143 == 32'h0000_0008 ? TestBlock__A_op14 : array_index_71142[8];
  assign array_update_71146[9] = add_71143 == 32'h0000_0009 ? TestBlock__A_op14 : array_index_71142[9];
  assign array_update_71147[0] = add_71145 == 32'h0000_0000 ? TestBlock__B_op14 : array_index_71144[0];
  assign array_update_71147[1] = add_71145 == 32'h0000_0001 ? TestBlock__B_op14 : array_index_71144[1];
  assign array_update_71147[2] = add_71145 == 32'h0000_0002 ? TestBlock__B_op14 : array_index_71144[2];
  assign array_update_71147[3] = add_71145 == 32'h0000_0003 ? TestBlock__B_op14 : array_index_71144[3];
  assign array_update_71147[4] = add_71145 == 32'h0000_0004 ? TestBlock__B_op14 : array_index_71144[4];
  assign array_update_71147[5] = add_71145 == 32'h0000_0005 ? TestBlock__B_op14 : array_index_71144[5];
  assign array_update_71147[6] = add_71145 == 32'h0000_0006 ? TestBlock__B_op14 : array_index_71144[6];
  assign array_update_71147[7] = add_71145 == 32'h0000_0007 ? TestBlock__B_op14 : array_index_71144[7];
  assign array_update_71147[8] = add_71145 == 32'h0000_0008 ? TestBlock__B_op14 : array_index_71144[8];
  assign array_update_71147[9] = add_71145 == 32'h0000_0009 ? TestBlock__B_op14 : array_index_71144[9];
  assign array_update_71148[0] = add_71099 == 32'h0000_0000 ? array_update_71146 : array_update_71138[0];
  assign array_update_71148[1] = add_71099 == 32'h0000_0001 ? array_update_71146 : array_update_71138[1];
  assign array_update_71148[2] = add_71099 == 32'h0000_0002 ? array_update_71146 : array_update_71138[2];
  assign array_update_71148[3] = add_71099 == 32'h0000_0003 ? array_update_71146 : array_update_71138[3];
  assign array_update_71148[4] = add_71099 == 32'h0000_0004 ? array_update_71146 : array_update_71138[4];
  assign array_update_71148[5] = add_71099 == 32'h0000_0005 ? array_update_71146 : array_update_71138[5];
  assign array_update_71148[6] = add_71099 == 32'h0000_0006 ? array_update_71146 : array_update_71138[6];
  assign array_update_71148[7] = add_71099 == 32'h0000_0007 ? array_update_71146 : array_update_71138[7];
  assign array_update_71148[8] = add_71099 == 32'h0000_0008 ? array_update_71146 : array_update_71138[8];
  assign array_update_71148[9] = add_71099 == 32'h0000_0009 ? array_update_71146 : array_update_71138[9];
  assign array_update_71150[0] = add_71101 == 32'h0000_0000 ? array_update_71147 : array_update_71140[0];
  assign array_update_71150[1] = add_71101 == 32'h0000_0001 ? array_update_71147 : array_update_71140[1];
  assign array_update_71150[2] = add_71101 == 32'h0000_0002 ? array_update_71147 : array_update_71140[2];
  assign array_update_71150[3] = add_71101 == 32'h0000_0003 ? array_update_71147 : array_update_71140[3];
  assign array_update_71150[4] = add_71101 == 32'h0000_0004 ? array_update_71147 : array_update_71140[4];
  assign array_update_71150[5] = add_71101 == 32'h0000_0005 ? array_update_71147 : array_update_71140[5];
  assign array_update_71150[6] = add_71101 == 32'h0000_0006 ? array_update_71147 : array_update_71140[6];
  assign array_update_71150[7] = add_71101 == 32'h0000_0007 ? array_update_71147 : array_update_71140[7];
  assign array_update_71150[8] = add_71101 == 32'h0000_0008 ? array_update_71147 : array_update_71140[8];
  assign array_update_71150[9] = add_71101 == 32'h0000_0009 ? array_update_71147 : array_update_71140[9];
  assign array_index_71152 = array_update_71148[add_71099 > 32'h0000_0009 ? 4'h9 : add_71099[3:0]];
  assign add_71153 = add_71143 + 32'h0000_0001;
  assign array_index_71154 = array_update_71150[add_71101 > 32'h0000_0009 ? 4'h9 : add_71101[3:0]];
  assign add_71155 = add_71145 + 32'h0000_0001;
  assign array_update_71156[0] = add_71153 == 32'h0000_0000 ? TestBlock__A_op15 : array_index_71152[0];
  assign array_update_71156[1] = add_71153 == 32'h0000_0001 ? TestBlock__A_op15 : array_index_71152[1];
  assign array_update_71156[2] = add_71153 == 32'h0000_0002 ? TestBlock__A_op15 : array_index_71152[2];
  assign array_update_71156[3] = add_71153 == 32'h0000_0003 ? TestBlock__A_op15 : array_index_71152[3];
  assign array_update_71156[4] = add_71153 == 32'h0000_0004 ? TestBlock__A_op15 : array_index_71152[4];
  assign array_update_71156[5] = add_71153 == 32'h0000_0005 ? TestBlock__A_op15 : array_index_71152[5];
  assign array_update_71156[6] = add_71153 == 32'h0000_0006 ? TestBlock__A_op15 : array_index_71152[6];
  assign array_update_71156[7] = add_71153 == 32'h0000_0007 ? TestBlock__A_op15 : array_index_71152[7];
  assign array_update_71156[8] = add_71153 == 32'h0000_0008 ? TestBlock__A_op15 : array_index_71152[8];
  assign array_update_71156[9] = add_71153 == 32'h0000_0009 ? TestBlock__A_op15 : array_index_71152[9];
  assign array_update_71157[0] = add_71155 == 32'h0000_0000 ? TestBlock__B_op15 : array_index_71154[0];
  assign array_update_71157[1] = add_71155 == 32'h0000_0001 ? TestBlock__B_op15 : array_index_71154[1];
  assign array_update_71157[2] = add_71155 == 32'h0000_0002 ? TestBlock__B_op15 : array_index_71154[2];
  assign array_update_71157[3] = add_71155 == 32'h0000_0003 ? TestBlock__B_op15 : array_index_71154[3];
  assign array_update_71157[4] = add_71155 == 32'h0000_0004 ? TestBlock__B_op15 : array_index_71154[4];
  assign array_update_71157[5] = add_71155 == 32'h0000_0005 ? TestBlock__B_op15 : array_index_71154[5];
  assign array_update_71157[6] = add_71155 == 32'h0000_0006 ? TestBlock__B_op15 : array_index_71154[6];
  assign array_update_71157[7] = add_71155 == 32'h0000_0007 ? TestBlock__B_op15 : array_index_71154[7];
  assign array_update_71157[8] = add_71155 == 32'h0000_0008 ? TestBlock__B_op15 : array_index_71154[8];
  assign array_update_71157[9] = add_71155 == 32'h0000_0009 ? TestBlock__B_op15 : array_index_71154[9];
  assign array_update_71158[0] = add_71099 == 32'h0000_0000 ? array_update_71156 : array_update_71148[0];
  assign array_update_71158[1] = add_71099 == 32'h0000_0001 ? array_update_71156 : array_update_71148[1];
  assign array_update_71158[2] = add_71099 == 32'h0000_0002 ? array_update_71156 : array_update_71148[2];
  assign array_update_71158[3] = add_71099 == 32'h0000_0003 ? array_update_71156 : array_update_71148[3];
  assign array_update_71158[4] = add_71099 == 32'h0000_0004 ? array_update_71156 : array_update_71148[4];
  assign array_update_71158[5] = add_71099 == 32'h0000_0005 ? array_update_71156 : array_update_71148[5];
  assign array_update_71158[6] = add_71099 == 32'h0000_0006 ? array_update_71156 : array_update_71148[6];
  assign array_update_71158[7] = add_71099 == 32'h0000_0007 ? array_update_71156 : array_update_71148[7];
  assign array_update_71158[8] = add_71099 == 32'h0000_0008 ? array_update_71156 : array_update_71148[8];
  assign array_update_71158[9] = add_71099 == 32'h0000_0009 ? array_update_71156 : array_update_71148[9];
  assign array_update_71160[0] = add_71101 == 32'h0000_0000 ? array_update_71157 : array_update_71150[0];
  assign array_update_71160[1] = add_71101 == 32'h0000_0001 ? array_update_71157 : array_update_71150[1];
  assign array_update_71160[2] = add_71101 == 32'h0000_0002 ? array_update_71157 : array_update_71150[2];
  assign array_update_71160[3] = add_71101 == 32'h0000_0003 ? array_update_71157 : array_update_71150[3];
  assign array_update_71160[4] = add_71101 == 32'h0000_0004 ? array_update_71157 : array_update_71150[4];
  assign array_update_71160[5] = add_71101 == 32'h0000_0005 ? array_update_71157 : array_update_71150[5];
  assign array_update_71160[6] = add_71101 == 32'h0000_0006 ? array_update_71157 : array_update_71150[6];
  assign array_update_71160[7] = add_71101 == 32'h0000_0007 ? array_update_71157 : array_update_71150[7];
  assign array_update_71160[8] = add_71101 == 32'h0000_0008 ? array_update_71157 : array_update_71150[8];
  assign array_update_71160[9] = add_71101 == 32'h0000_0009 ? array_update_71157 : array_update_71150[9];
  assign array_index_71162 = array_update_71158[add_71099 > 32'h0000_0009 ? 4'h9 : add_71099[3:0]];
  assign add_71163 = add_71153 + 32'h0000_0001;
  assign array_index_71164 = array_update_71160[add_71101 > 32'h0000_0009 ? 4'h9 : add_71101[3:0]];
  assign add_71165 = add_71155 + 32'h0000_0001;
  assign array_update_71166[0] = add_71163 == 32'h0000_0000 ? TestBlock__A_op16 : array_index_71162[0];
  assign array_update_71166[1] = add_71163 == 32'h0000_0001 ? TestBlock__A_op16 : array_index_71162[1];
  assign array_update_71166[2] = add_71163 == 32'h0000_0002 ? TestBlock__A_op16 : array_index_71162[2];
  assign array_update_71166[3] = add_71163 == 32'h0000_0003 ? TestBlock__A_op16 : array_index_71162[3];
  assign array_update_71166[4] = add_71163 == 32'h0000_0004 ? TestBlock__A_op16 : array_index_71162[4];
  assign array_update_71166[5] = add_71163 == 32'h0000_0005 ? TestBlock__A_op16 : array_index_71162[5];
  assign array_update_71166[6] = add_71163 == 32'h0000_0006 ? TestBlock__A_op16 : array_index_71162[6];
  assign array_update_71166[7] = add_71163 == 32'h0000_0007 ? TestBlock__A_op16 : array_index_71162[7];
  assign array_update_71166[8] = add_71163 == 32'h0000_0008 ? TestBlock__A_op16 : array_index_71162[8];
  assign array_update_71166[9] = add_71163 == 32'h0000_0009 ? TestBlock__A_op16 : array_index_71162[9];
  assign array_update_71167[0] = add_71165 == 32'h0000_0000 ? TestBlock__B_op16 : array_index_71164[0];
  assign array_update_71167[1] = add_71165 == 32'h0000_0001 ? TestBlock__B_op16 : array_index_71164[1];
  assign array_update_71167[2] = add_71165 == 32'h0000_0002 ? TestBlock__B_op16 : array_index_71164[2];
  assign array_update_71167[3] = add_71165 == 32'h0000_0003 ? TestBlock__B_op16 : array_index_71164[3];
  assign array_update_71167[4] = add_71165 == 32'h0000_0004 ? TestBlock__B_op16 : array_index_71164[4];
  assign array_update_71167[5] = add_71165 == 32'h0000_0005 ? TestBlock__B_op16 : array_index_71164[5];
  assign array_update_71167[6] = add_71165 == 32'h0000_0006 ? TestBlock__B_op16 : array_index_71164[6];
  assign array_update_71167[7] = add_71165 == 32'h0000_0007 ? TestBlock__B_op16 : array_index_71164[7];
  assign array_update_71167[8] = add_71165 == 32'h0000_0008 ? TestBlock__B_op16 : array_index_71164[8];
  assign array_update_71167[9] = add_71165 == 32'h0000_0009 ? TestBlock__B_op16 : array_index_71164[9];
  assign array_update_71168[0] = add_71099 == 32'h0000_0000 ? array_update_71166 : array_update_71158[0];
  assign array_update_71168[1] = add_71099 == 32'h0000_0001 ? array_update_71166 : array_update_71158[1];
  assign array_update_71168[2] = add_71099 == 32'h0000_0002 ? array_update_71166 : array_update_71158[2];
  assign array_update_71168[3] = add_71099 == 32'h0000_0003 ? array_update_71166 : array_update_71158[3];
  assign array_update_71168[4] = add_71099 == 32'h0000_0004 ? array_update_71166 : array_update_71158[4];
  assign array_update_71168[5] = add_71099 == 32'h0000_0005 ? array_update_71166 : array_update_71158[5];
  assign array_update_71168[6] = add_71099 == 32'h0000_0006 ? array_update_71166 : array_update_71158[6];
  assign array_update_71168[7] = add_71099 == 32'h0000_0007 ? array_update_71166 : array_update_71158[7];
  assign array_update_71168[8] = add_71099 == 32'h0000_0008 ? array_update_71166 : array_update_71158[8];
  assign array_update_71168[9] = add_71099 == 32'h0000_0009 ? array_update_71166 : array_update_71158[9];
  assign array_update_71170[0] = add_71101 == 32'h0000_0000 ? array_update_71167 : array_update_71160[0];
  assign array_update_71170[1] = add_71101 == 32'h0000_0001 ? array_update_71167 : array_update_71160[1];
  assign array_update_71170[2] = add_71101 == 32'h0000_0002 ? array_update_71167 : array_update_71160[2];
  assign array_update_71170[3] = add_71101 == 32'h0000_0003 ? array_update_71167 : array_update_71160[3];
  assign array_update_71170[4] = add_71101 == 32'h0000_0004 ? array_update_71167 : array_update_71160[4];
  assign array_update_71170[5] = add_71101 == 32'h0000_0005 ? array_update_71167 : array_update_71160[5];
  assign array_update_71170[6] = add_71101 == 32'h0000_0006 ? array_update_71167 : array_update_71160[6];
  assign array_update_71170[7] = add_71101 == 32'h0000_0007 ? array_update_71167 : array_update_71160[7];
  assign array_update_71170[8] = add_71101 == 32'h0000_0008 ? array_update_71167 : array_update_71160[8];
  assign array_update_71170[9] = add_71101 == 32'h0000_0009 ? array_update_71167 : array_update_71160[9];
  assign array_index_71172 = array_update_71168[add_71099 > 32'h0000_0009 ? 4'h9 : add_71099[3:0]];
  assign add_71173 = add_71163 + 32'h0000_0001;
  assign array_index_71174 = array_update_71170[add_71101 > 32'h0000_0009 ? 4'h9 : add_71101[3:0]];
  assign add_71175 = add_71165 + 32'h0000_0001;
  assign array_update_71176[0] = add_71173 == 32'h0000_0000 ? TestBlock__A_op17 : array_index_71172[0];
  assign array_update_71176[1] = add_71173 == 32'h0000_0001 ? TestBlock__A_op17 : array_index_71172[1];
  assign array_update_71176[2] = add_71173 == 32'h0000_0002 ? TestBlock__A_op17 : array_index_71172[2];
  assign array_update_71176[3] = add_71173 == 32'h0000_0003 ? TestBlock__A_op17 : array_index_71172[3];
  assign array_update_71176[4] = add_71173 == 32'h0000_0004 ? TestBlock__A_op17 : array_index_71172[4];
  assign array_update_71176[5] = add_71173 == 32'h0000_0005 ? TestBlock__A_op17 : array_index_71172[5];
  assign array_update_71176[6] = add_71173 == 32'h0000_0006 ? TestBlock__A_op17 : array_index_71172[6];
  assign array_update_71176[7] = add_71173 == 32'h0000_0007 ? TestBlock__A_op17 : array_index_71172[7];
  assign array_update_71176[8] = add_71173 == 32'h0000_0008 ? TestBlock__A_op17 : array_index_71172[8];
  assign array_update_71176[9] = add_71173 == 32'h0000_0009 ? TestBlock__A_op17 : array_index_71172[9];
  assign array_update_71177[0] = add_71175 == 32'h0000_0000 ? TestBlock__B_op17 : array_index_71174[0];
  assign array_update_71177[1] = add_71175 == 32'h0000_0001 ? TestBlock__B_op17 : array_index_71174[1];
  assign array_update_71177[2] = add_71175 == 32'h0000_0002 ? TestBlock__B_op17 : array_index_71174[2];
  assign array_update_71177[3] = add_71175 == 32'h0000_0003 ? TestBlock__B_op17 : array_index_71174[3];
  assign array_update_71177[4] = add_71175 == 32'h0000_0004 ? TestBlock__B_op17 : array_index_71174[4];
  assign array_update_71177[5] = add_71175 == 32'h0000_0005 ? TestBlock__B_op17 : array_index_71174[5];
  assign array_update_71177[6] = add_71175 == 32'h0000_0006 ? TestBlock__B_op17 : array_index_71174[6];
  assign array_update_71177[7] = add_71175 == 32'h0000_0007 ? TestBlock__B_op17 : array_index_71174[7];
  assign array_update_71177[8] = add_71175 == 32'h0000_0008 ? TestBlock__B_op17 : array_index_71174[8];
  assign array_update_71177[9] = add_71175 == 32'h0000_0009 ? TestBlock__B_op17 : array_index_71174[9];
  assign array_update_71178[0] = add_71099 == 32'h0000_0000 ? array_update_71176 : array_update_71168[0];
  assign array_update_71178[1] = add_71099 == 32'h0000_0001 ? array_update_71176 : array_update_71168[1];
  assign array_update_71178[2] = add_71099 == 32'h0000_0002 ? array_update_71176 : array_update_71168[2];
  assign array_update_71178[3] = add_71099 == 32'h0000_0003 ? array_update_71176 : array_update_71168[3];
  assign array_update_71178[4] = add_71099 == 32'h0000_0004 ? array_update_71176 : array_update_71168[4];
  assign array_update_71178[5] = add_71099 == 32'h0000_0005 ? array_update_71176 : array_update_71168[5];
  assign array_update_71178[6] = add_71099 == 32'h0000_0006 ? array_update_71176 : array_update_71168[6];
  assign array_update_71178[7] = add_71099 == 32'h0000_0007 ? array_update_71176 : array_update_71168[7];
  assign array_update_71178[8] = add_71099 == 32'h0000_0008 ? array_update_71176 : array_update_71168[8];
  assign array_update_71178[9] = add_71099 == 32'h0000_0009 ? array_update_71176 : array_update_71168[9];
  assign array_update_71180[0] = add_71101 == 32'h0000_0000 ? array_update_71177 : array_update_71170[0];
  assign array_update_71180[1] = add_71101 == 32'h0000_0001 ? array_update_71177 : array_update_71170[1];
  assign array_update_71180[2] = add_71101 == 32'h0000_0002 ? array_update_71177 : array_update_71170[2];
  assign array_update_71180[3] = add_71101 == 32'h0000_0003 ? array_update_71177 : array_update_71170[3];
  assign array_update_71180[4] = add_71101 == 32'h0000_0004 ? array_update_71177 : array_update_71170[4];
  assign array_update_71180[5] = add_71101 == 32'h0000_0005 ? array_update_71177 : array_update_71170[5];
  assign array_update_71180[6] = add_71101 == 32'h0000_0006 ? array_update_71177 : array_update_71170[6];
  assign array_update_71180[7] = add_71101 == 32'h0000_0007 ? array_update_71177 : array_update_71170[7];
  assign array_update_71180[8] = add_71101 == 32'h0000_0008 ? array_update_71177 : array_update_71170[8];
  assign array_update_71180[9] = add_71101 == 32'h0000_0009 ? array_update_71177 : array_update_71170[9];
  assign array_index_71182 = array_update_71178[add_71099 > 32'h0000_0009 ? 4'h9 : add_71099[3:0]];
  assign add_71183 = add_71173 + 32'h0000_0001;
  assign array_index_71184 = array_update_71180[add_71101 > 32'h0000_0009 ? 4'h9 : add_71101[3:0]];
  assign add_71185 = add_71175 + 32'h0000_0001;
  assign array_update_71186[0] = add_71183 == 32'h0000_0000 ? TestBlock__A_op18 : array_index_71182[0];
  assign array_update_71186[1] = add_71183 == 32'h0000_0001 ? TestBlock__A_op18 : array_index_71182[1];
  assign array_update_71186[2] = add_71183 == 32'h0000_0002 ? TestBlock__A_op18 : array_index_71182[2];
  assign array_update_71186[3] = add_71183 == 32'h0000_0003 ? TestBlock__A_op18 : array_index_71182[3];
  assign array_update_71186[4] = add_71183 == 32'h0000_0004 ? TestBlock__A_op18 : array_index_71182[4];
  assign array_update_71186[5] = add_71183 == 32'h0000_0005 ? TestBlock__A_op18 : array_index_71182[5];
  assign array_update_71186[6] = add_71183 == 32'h0000_0006 ? TestBlock__A_op18 : array_index_71182[6];
  assign array_update_71186[7] = add_71183 == 32'h0000_0007 ? TestBlock__A_op18 : array_index_71182[7];
  assign array_update_71186[8] = add_71183 == 32'h0000_0008 ? TestBlock__A_op18 : array_index_71182[8];
  assign array_update_71186[9] = add_71183 == 32'h0000_0009 ? TestBlock__A_op18 : array_index_71182[9];
  assign array_update_71187[0] = add_71185 == 32'h0000_0000 ? TestBlock__B_op18 : array_index_71184[0];
  assign array_update_71187[1] = add_71185 == 32'h0000_0001 ? TestBlock__B_op18 : array_index_71184[1];
  assign array_update_71187[2] = add_71185 == 32'h0000_0002 ? TestBlock__B_op18 : array_index_71184[2];
  assign array_update_71187[3] = add_71185 == 32'h0000_0003 ? TestBlock__B_op18 : array_index_71184[3];
  assign array_update_71187[4] = add_71185 == 32'h0000_0004 ? TestBlock__B_op18 : array_index_71184[4];
  assign array_update_71187[5] = add_71185 == 32'h0000_0005 ? TestBlock__B_op18 : array_index_71184[5];
  assign array_update_71187[6] = add_71185 == 32'h0000_0006 ? TestBlock__B_op18 : array_index_71184[6];
  assign array_update_71187[7] = add_71185 == 32'h0000_0007 ? TestBlock__B_op18 : array_index_71184[7];
  assign array_update_71187[8] = add_71185 == 32'h0000_0008 ? TestBlock__B_op18 : array_index_71184[8];
  assign array_update_71187[9] = add_71185 == 32'h0000_0009 ? TestBlock__B_op18 : array_index_71184[9];
  assign array_update_71188[0] = add_71099 == 32'h0000_0000 ? array_update_71186 : array_update_71178[0];
  assign array_update_71188[1] = add_71099 == 32'h0000_0001 ? array_update_71186 : array_update_71178[1];
  assign array_update_71188[2] = add_71099 == 32'h0000_0002 ? array_update_71186 : array_update_71178[2];
  assign array_update_71188[3] = add_71099 == 32'h0000_0003 ? array_update_71186 : array_update_71178[3];
  assign array_update_71188[4] = add_71099 == 32'h0000_0004 ? array_update_71186 : array_update_71178[4];
  assign array_update_71188[5] = add_71099 == 32'h0000_0005 ? array_update_71186 : array_update_71178[5];
  assign array_update_71188[6] = add_71099 == 32'h0000_0006 ? array_update_71186 : array_update_71178[6];
  assign array_update_71188[7] = add_71099 == 32'h0000_0007 ? array_update_71186 : array_update_71178[7];
  assign array_update_71188[8] = add_71099 == 32'h0000_0008 ? array_update_71186 : array_update_71178[8];
  assign array_update_71188[9] = add_71099 == 32'h0000_0009 ? array_update_71186 : array_update_71178[9];
  assign array_update_71190[0] = add_71101 == 32'h0000_0000 ? array_update_71187 : array_update_71180[0];
  assign array_update_71190[1] = add_71101 == 32'h0000_0001 ? array_update_71187 : array_update_71180[1];
  assign array_update_71190[2] = add_71101 == 32'h0000_0002 ? array_update_71187 : array_update_71180[2];
  assign array_update_71190[3] = add_71101 == 32'h0000_0003 ? array_update_71187 : array_update_71180[3];
  assign array_update_71190[4] = add_71101 == 32'h0000_0004 ? array_update_71187 : array_update_71180[4];
  assign array_update_71190[5] = add_71101 == 32'h0000_0005 ? array_update_71187 : array_update_71180[5];
  assign array_update_71190[6] = add_71101 == 32'h0000_0006 ? array_update_71187 : array_update_71180[6];
  assign array_update_71190[7] = add_71101 == 32'h0000_0007 ? array_update_71187 : array_update_71180[7];
  assign array_update_71190[8] = add_71101 == 32'h0000_0008 ? array_update_71187 : array_update_71180[8];
  assign array_update_71190[9] = add_71101 == 32'h0000_0009 ? array_update_71187 : array_update_71180[9];
  assign array_index_71192 = array_update_71188[add_71099 > 32'h0000_0009 ? 4'h9 : add_71099[3:0]];
  assign add_71193 = add_71183 + 32'h0000_0001;
  assign array_index_71194 = array_update_71190[add_71101 > 32'h0000_0009 ? 4'h9 : add_71101[3:0]];
  assign add_71195 = add_71185 + 32'h0000_0001;
  assign array_update_71196[0] = add_71193 == 32'h0000_0000 ? TestBlock__A_op19 : array_index_71192[0];
  assign array_update_71196[1] = add_71193 == 32'h0000_0001 ? TestBlock__A_op19 : array_index_71192[1];
  assign array_update_71196[2] = add_71193 == 32'h0000_0002 ? TestBlock__A_op19 : array_index_71192[2];
  assign array_update_71196[3] = add_71193 == 32'h0000_0003 ? TestBlock__A_op19 : array_index_71192[3];
  assign array_update_71196[4] = add_71193 == 32'h0000_0004 ? TestBlock__A_op19 : array_index_71192[4];
  assign array_update_71196[5] = add_71193 == 32'h0000_0005 ? TestBlock__A_op19 : array_index_71192[5];
  assign array_update_71196[6] = add_71193 == 32'h0000_0006 ? TestBlock__A_op19 : array_index_71192[6];
  assign array_update_71196[7] = add_71193 == 32'h0000_0007 ? TestBlock__A_op19 : array_index_71192[7];
  assign array_update_71196[8] = add_71193 == 32'h0000_0008 ? TestBlock__A_op19 : array_index_71192[8];
  assign array_update_71196[9] = add_71193 == 32'h0000_0009 ? TestBlock__A_op19 : array_index_71192[9];
  assign array_update_71198[0] = add_71195 == 32'h0000_0000 ? TestBlock__B_op19 : array_index_71194[0];
  assign array_update_71198[1] = add_71195 == 32'h0000_0001 ? TestBlock__B_op19 : array_index_71194[1];
  assign array_update_71198[2] = add_71195 == 32'h0000_0002 ? TestBlock__B_op19 : array_index_71194[2];
  assign array_update_71198[3] = add_71195 == 32'h0000_0003 ? TestBlock__B_op19 : array_index_71194[3];
  assign array_update_71198[4] = add_71195 == 32'h0000_0004 ? TestBlock__B_op19 : array_index_71194[4];
  assign array_update_71198[5] = add_71195 == 32'h0000_0005 ? TestBlock__B_op19 : array_index_71194[5];
  assign array_update_71198[6] = add_71195 == 32'h0000_0006 ? TestBlock__B_op19 : array_index_71194[6];
  assign array_update_71198[7] = add_71195 == 32'h0000_0007 ? TestBlock__B_op19 : array_index_71194[7];
  assign array_update_71198[8] = add_71195 == 32'h0000_0008 ? TestBlock__B_op19 : array_index_71194[8];
  assign array_update_71198[9] = add_71195 == 32'h0000_0009 ? TestBlock__B_op19 : array_index_71194[9];
  assign array_update_71200[0] = add_71099 == 32'h0000_0000 ? array_update_71196 : array_update_71188[0];
  assign array_update_71200[1] = add_71099 == 32'h0000_0001 ? array_update_71196 : array_update_71188[1];
  assign array_update_71200[2] = add_71099 == 32'h0000_0002 ? array_update_71196 : array_update_71188[2];
  assign array_update_71200[3] = add_71099 == 32'h0000_0003 ? array_update_71196 : array_update_71188[3];
  assign array_update_71200[4] = add_71099 == 32'h0000_0004 ? array_update_71196 : array_update_71188[4];
  assign array_update_71200[5] = add_71099 == 32'h0000_0005 ? array_update_71196 : array_update_71188[5];
  assign array_update_71200[6] = add_71099 == 32'h0000_0006 ? array_update_71196 : array_update_71188[6];
  assign array_update_71200[7] = add_71099 == 32'h0000_0007 ? array_update_71196 : array_update_71188[7];
  assign array_update_71200[8] = add_71099 == 32'h0000_0008 ? array_update_71196 : array_update_71188[8];
  assign array_update_71200[9] = add_71099 == 32'h0000_0009 ? array_update_71196 : array_update_71188[9];
  assign add_71201 = add_71099 + 32'h0000_0001;
  assign array_update_71202[0] = add_71101 == 32'h0000_0000 ? array_update_71198 : array_update_71190[0];
  assign array_update_71202[1] = add_71101 == 32'h0000_0001 ? array_update_71198 : array_update_71190[1];
  assign array_update_71202[2] = add_71101 == 32'h0000_0002 ? array_update_71198 : array_update_71190[2];
  assign array_update_71202[3] = add_71101 == 32'h0000_0003 ? array_update_71198 : array_update_71190[3];
  assign array_update_71202[4] = add_71101 == 32'h0000_0004 ? array_update_71198 : array_update_71190[4];
  assign array_update_71202[5] = add_71101 == 32'h0000_0005 ? array_update_71198 : array_update_71190[5];
  assign array_update_71202[6] = add_71101 == 32'h0000_0006 ? array_update_71198 : array_update_71190[6];
  assign array_update_71202[7] = add_71101 == 32'h0000_0007 ? array_update_71198 : array_update_71190[7];
  assign array_update_71202[8] = add_71101 == 32'h0000_0008 ? array_update_71198 : array_update_71190[8];
  assign array_update_71202[9] = add_71101 == 32'h0000_0009 ? array_update_71198 : array_update_71190[9];
  assign add_71203 = add_71101 + 32'h0000_0001;
  assign array_index_71204 = array_update_71200[add_71201 > 32'h0000_0009 ? 4'h9 : add_71201[3:0]];
  assign literal_71205 = 32'h0000_0000;
  assign array_index_71206 = array_update_71202[add_71203 > 32'h0000_0009 ? 4'h9 : add_71203[3:0]];
  assign literal_71207 = 32'h0000_0000;
  assign array_update_71208[0] = literal_71205 == 32'h0000_0000 ? TestBlock__A_op20 : array_index_71204[0];
  assign array_update_71208[1] = literal_71205 == 32'h0000_0001 ? TestBlock__A_op20 : array_index_71204[1];
  assign array_update_71208[2] = literal_71205 == 32'h0000_0002 ? TestBlock__A_op20 : array_index_71204[2];
  assign array_update_71208[3] = literal_71205 == 32'h0000_0003 ? TestBlock__A_op20 : array_index_71204[3];
  assign array_update_71208[4] = literal_71205 == 32'h0000_0004 ? TestBlock__A_op20 : array_index_71204[4];
  assign array_update_71208[5] = literal_71205 == 32'h0000_0005 ? TestBlock__A_op20 : array_index_71204[5];
  assign array_update_71208[6] = literal_71205 == 32'h0000_0006 ? TestBlock__A_op20 : array_index_71204[6];
  assign array_update_71208[7] = literal_71205 == 32'h0000_0007 ? TestBlock__A_op20 : array_index_71204[7];
  assign array_update_71208[8] = literal_71205 == 32'h0000_0008 ? TestBlock__A_op20 : array_index_71204[8];
  assign array_update_71208[9] = literal_71205 == 32'h0000_0009 ? TestBlock__A_op20 : array_index_71204[9];
  assign array_update_71209[0] = literal_71207 == 32'h0000_0000 ? TestBlock__B_op20 : array_index_71206[0];
  assign array_update_71209[1] = literal_71207 == 32'h0000_0001 ? TestBlock__B_op20 : array_index_71206[1];
  assign array_update_71209[2] = literal_71207 == 32'h0000_0002 ? TestBlock__B_op20 : array_index_71206[2];
  assign array_update_71209[3] = literal_71207 == 32'h0000_0003 ? TestBlock__B_op20 : array_index_71206[3];
  assign array_update_71209[4] = literal_71207 == 32'h0000_0004 ? TestBlock__B_op20 : array_index_71206[4];
  assign array_update_71209[5] = literal_71207 == 32'h0000_0005 ? TestBlock__B_op20 : array_index_71206[5];
  assign array_update_71209[6] = literal_71207 == 32'h0000_0006 ? TestBlock__B_op20 : array_index_71206[6];
  assign array_update_71209[7] = literal_71207 == 32'h0000_0007 ? TestBlock__B_op20 : array_index_71206[7];
  assign array_update_71209[8] = literal_71207 == 32'h0000_0008 ? TestBlock__B_op20 : array_index_71206[8];
  assign array_update_71209[9] = literal_71207 == 32'h0000_0009 ? TestBlock__B_op20 : array_index_71206[9];
  assign array_update_71210[0] = add_71201 == 32'h0000_0000 ? array_update_71208 : array_update_71200[0];
  assign array_update_71210[1] = add_71201 == 32'h0000_0001 ? array_update_71208 : array_update_71200[1];
  assign array_update_71210[2] = add_71201 == 32'h0000_0002 ? array_update_71208 : array_update_71200[2];
  assign array_update_71210[3] = add_71201 == 32'h0000_0003 ? array_update_71208 : array_update_71200[3];
  assign array_update_71210[4] = add_71201 == 32'h0000_0004 ? array_update_71208 : array_update_71200[4];
  assign array_update_71210[5] = add_71201 == 32'h0000_0005 ? array_update_71208 : array_update_71200[5];
  assign array_update_71210[6] = add_71201 == 32'h0000_0006 ? array_update_71208 : array_update_71200[6];
  assign array_update_71210[7] = add_71201 == 32'h0000_0007 ? array_update_71208 : array_update_71200[7];
  assign array_update_71210[8] = add_71201 == 32'h0000_0008 ? array_update_71208 : array_update_71200[8];
  assign array_update_71210[9] = add_71201 == 32'h0000_0009 ? array_update_71208 : array_update_71200[9];
  assign array_update_71212[0] = add_71203 == 32'h0000_0000 ? array_update_71209 : array_update_71202[0];
  assign array_update_71212[1] = add_71203 == 32'h0000_0001 ? array_update_71209 : array_update_71202[1];
  assign array_update_71212[2] = add_71203 == 32'h0000_0002 ? array_update_71209 : array_update_71202[2];
  assign array_update_71212[3] = add_71203 == 32'h0000_0003 ? array_update_71209 : array_update_71202[3];
  assign array_update_71212[4] = add_71203 == 32'h0000_0004 ? array_update_71209 : array_update_71202[4];
  assign array_update_71212[5] = add_71203 == 32'h0000_0005 ? array_update_71209 : array_update_71202[5];
  assign array_update_71212[6] = add_71203 == 32'h0000_0006 ? array_update_71209 : array_update_71202[6];
  assign array_update_71212[7] = add_71203 == 32'h0000_0007 ? array_update_71209 : array_update_71202[7];
  assign array_update_71212[8] = add_71203 == 32'h0000_0008 ? array_update_71209 : array_update_71202[8];
  assign array_update_71212[9] = add_71203 == 32'h0000_0009 ? array_update_71209 : array_update_71202[9];
  assign array_index_71214 = array_update_71210[add_71201 > 32'h0000_0009 ? 4'h9 : add_71201[3:0]];
  assign add_71215 = literal_71205 + 32'h0000_0001;
  assign array_index_71216 = array_update_71212[add_71203 > 32'h0000_0009 ? 4'h9 : add_71203[3:0]];
  assign add_71217 = literal_71207 + 32'h0000_0001;
  assign array_update_71218[0] = add_71215 == 32'h0000_0000 ? TestBlock__A_op21 : array_index_71214[0];
  assign array_update_71218[1] = add_71215 == 32'h0000_0001 ? TestBlock__A_op21 : array_index_71214[1];
  assign array_update_71218[2] = add_71215 == 32'h0000_0002 ? TestBlock__A_op21 : array_index_71214[2];
  assign array_update_71218[3] = add_71215 == 32'h0000_0003 ? TestBlock__A_op21 : array_index_71214[3];
  assign array_update_71218[4] = add_71215 == 32'h0000_0004 ? TestBlock__A_op21 : array_index_71214[4];
  assign array_update_71218[5] = add_71215 == 32'h0000_0005 ? TestBlock__A_op21 : array_index_71214[5];
  assign array_update_71218[6] = add_71215 == 32'h0000_0006 ? TestBlock__A_op21 : array_index_71214[6];
  assign array_update_71218[7] = add_71215 == 32'h0000_0007 ? TestBlock__A_op21 : array_index_71214[7];
  assign array_update_71218[8] = add_71215 == 32'h0000_0008 ? TestBlock__A_op21 : array_index_71214[8];
  assign array_update_71218[9] = add_71215 == 32'h0000_0009 ? TestBlock__A_op21 : array_index_71214[9];
  assign array_update_71219[0] = add_71217 == 32'h0000_0000 ? TestBlock__B_op21 : array_index_71216[0];
  assign array_update_71219[1] = add_71217 == 32'h0000_0001 ? TestBlock__B_op21 : array_index_71216[1];
  assign array_update_71219[2] = add_71217 == 32'h0000_0002 ? TestBlock__B_op21 : array_index_71216[2];
  assign array_update_71219[3] = add_71217 == 32'h0000_0003 ? TestBlock__B_op21 : array_index_71216[3];
  assign array_update_71219[4] = add_71217 == 32'h0000_0004 ? TestBlock__B_op21 : array_index_71216[4];
  assign array_update_71219[5] = add_71217 == 32'h0000_0005 ? TestBlock__B_op21 : array_index_71216[5];
  assign array_update_71219[6] = add_71217 == 32'h0000_0006 ? TestBlock__B_op21 : array_index_71216[6];
  assign array_update_71219[7] = add_71217 == 32'h0000_0007 ? TestBlock__B_op21 : array_index_71216[7];
  assign array_update_71219[8] = add_71217 == 32'h0000_0008 ? TestBlock__B_op21 : array_index_71216[8];
  assign array_update_71219[9] = add_71217 == 32'h0000_0009 ? TestBlock__B_op21 : array_index_71216[9];
  assign array_update_71220[0] = add_71201 == 32'h0000_0000 ? array_update_71218 : array_update_71210[0];
  assign array_update_71220[1] = add_71201 == 32'h0000_0001 ? array_update_71218 : array_update_71210[1];
  assign array_update_71220[2] = add_71201 == 32'h0000_0002 ? array_update_71218 : array_update_71210[2];
  assign array_update_71220[3] = add_71201 == 32'h0000_0003 ? array_update_71218 : array_update_71210[3];
  assign array_update_71220[4] = add_71201 == 32'h0000_0004 ? array_update_71218 : array_update_71210[4];
  assign array_update_71220[5] = add_71201 == 32'h0000_0005 ? array_update_71218 : array_update_71210[5];
  assign array_update_71220[6] = add_71201 == 32'h0000_0006 ? array_update_71218 : array_update_71210[6];
  assign array_update_71220[7] = add_71201 == 32'h0000_0007 ? array_update_71218 : array_update_71210[7];
  assign array_update_71220[8] = add_71201 == 32'h0000_0008 ? array_update_71218 : array_update_71210[8];
  assign array_update_71220[9] = add_71201 == 32'h0000_0009 ? array_update_71218 : array_update_71210[9];
  assign array_update_71222[0] = add_71203 == 32'h0000_0000 ? array_update_71219 : array_update_71212[0];
  assign array_update_71222[1] = add_71203 == 32'h0000_0001 ? array_update_71219 : array_update_71212[1];
  assign array_update_71222[2] = add_71203 == 32'h0000_0002 ? array_update_71219 : array_update_71212[2];
  assign array_update_71222[3] = add_71203 == 32'h0000_0003 ? array_update_71219 : array_update_71212[3];
  assign array_update_71222[4] = add_71203 == 32'h0000_0004 ? array_update_71219 : array_update_71212[4];
  assign array_update_71222[5] = add_71203 == 32'h0000_0005 ? array_update_71219 : array_update_71212[5];
  assign array_update_71222[6] = add_71203 == 32'h0000_0006 ? array_update_71219 : array_update_71212[6];
  assign array_update_71222[7] = add_71203 == 32'h0000_0007 ? array_update_71219 : array_update_71212[7];
  assign array_update_71222[8] = add_71203 == 32'h0000_0008 ? array_update_71219 : array_update_71212[8];
  assign array_update_71222[9] = add_71203 == 32'h0000_0009 ? array_update_71219 : array_update_71212[9];
  assign array_index_71224 = array_update_71220[add_71201 > 32'h0000_0009 ? 4'h9 : add_71201[3:0]];
  assign add_71225 = add_71215 + 32'h0000_0001;
  assign array_index_71226 = array_update_71222[add_71203 > 32'h0000_0009 ? 4'h9 : add_71203[3:0]];
  assign add_71227 = add_71217 + 32'h0000_0001;
  assign array_update_71228[0] = add_71225 == 32'h0000_0000 ? TestBlock__A_op22 : array_index_71224[0];
  assign array_update_71228[1] = add_71225 == 32'h0000_0001 ? TestBlock__A_op22 : array_index_71224[1];
  assign array_update_71228[2] = add_71225 == 32'h0000_0002 ? TestBlock__A_op22 : array_index_71224[2];
  assign array_update_71228[3] = add_71225 == 32'h0000_0003 ? TestBlock__A_op22 : array_index_71224[3];
  assign array_update_71228[4] = add_71225 == 32'h0000_0004 ? TestBlock__A_op22 : array_index_71224[4];
  assign array_update_71228[5] = add_71225 == 32'h0000_0005 ? TestBlock__A_op22 : array_index_71224[5];
  assign array_update_71228[6] = add_71225 == 32'h0000_0006 ? TestBlock__A_op22 : array_index_71224[6];
  assign array_update_71228[7] = add_71225 == 32'h0000_0007 ? TestBlock__A_op22 : array_index_71224[7];
  assign array_update_71228[8] = add_71225 == 32'h0000_0008 ? TestBlock__A_op22 : array_index_71224[8];
  assign array_update_71228[9] = add_71225 == 32'h0000_0009 ? TestBlock__A_op22 : array_index_71224[9];
  assign array_update_71229[0] = add_71227 == 32'h0000_0000 ? TestBlock__B_op22 : array_index_71226[0];
  assign array_update_71229[1] = add_71227 == 32'h0000_0001 ? TestBlock__B_op22 : array_index_71226[1];
  assign array_update_71229[2] = add_71227 == 32'h0000_0002 ? TestBlock__B_op22 : array_index_71226[2];
  assign array_update_71229[3] = add_71227 == 32'h0000_0003 ? TestBlock__B_op22 : array_index_71226[3];
  assign array_update_71229[4] = add_71227 == 32'h0000_0004 ? TestBlock__B_op22 : array_index_71226[4];
  assign array_update_71229[5] = add_71227 == 32'h0000_0005 ? TestBlock__B_op22 : array_index_71226[5];
  assign array_update_71229[6] = add_71227 == 32'h0000_0006 ? TestBlock__B_op22 : array_index_71226[6];
  assign array_update_71229[7] = add_71227 == 32'h0000_0007 ? TestBlock__B_op22 : array_index_71226[7];
  assign array_update_71229[8] = add_71227 == 32'h0000_0008 ? TestBlock__B_op22 : array_index_71226[8];
  assign array_update_71229[9] = add_71227 == 32'h0000_0009 ? TestBlock__B_op22 : array_index_71226[9];
  assign array_update_71230[0] = add_71201 == 32'h0000_0000 ? array_update_71228 : array_update_71220[0];
  assign array_update_71230[1] = add_71201 == 32'h0000_0001 ? array_update_71228 : array_update_71220[1];
  assign array_update_71230[2] = add_71201 == 32'h0000_0002 ? array_update_71228 : array_update_71220[2];
  assign array_update_71230[3] = add_71201 == 32'h0000_0003 ? array_update_71228 : array_update_71220[3];
  assign array_update_71230[4] = add_71201 == 32'h0000_0004 ? array_update_71228 : array_update_71220[4];
  assign array_update_71230[5] = add_71201 == 32'h0000_0005 ? array_update_71228 : array_update_71220[5];
  assign array_update_71230[6] = add_71201 == 32'h0000_0006 ? array_update_71228 : array_update_71220[6];
  assign array_update_71230[7] = add_71201 == 32'h0000_0007 ? array_update_71228 : array_update_71220[7];
  assign array_update_71230[8] = add_71201 == 32'h0000_0008 ? array_update_71228 : array_update_71220[8];
  assign array_update_71230[9] = add_71201 == 32'h0000_0009 ? array_update_71228 : array_update_71220[9];
  assign array_update_71232[0] = add_71203 == 32'h0000_0000 ? array_update_71229 : array_update_71222[0];
  assign array_update_71232[1] = add_71203 == 32'h0000_0001 ? array_update_71229 : array_update_71222[1];
  assign array_update_71232[2] = add_71203 == 32'h0000_0002 ? array_update_71229 : array_update_71222[2];
  assign array_update_71232[3] = add_71203 == 32'h0000_0003 ? array_update_71229 : array_update_71222[3];
  assign array_update_71232[4] = add_71203 == 32'h0000_0004 ? array_update_71229 : array_update_71222[4];
  assign array_update_71232[5] = add_71203 == 32'h0000_0005 ? array_update_71229 : array_update_71222[5];
  assign array_update_71232[6] = add_71203 == 32'h0000_0006 ? array_update_71229 : array_update_71222[6];
  assign array_update_71232[7] = add_71203 == 32'h0000_0007 ? array_update_71229 : array_update_71222[7];
  assign array_update_71232[8] = add_71203 == 32'h0000_0008 ? array_update_71229 : array_update_71222[8];
  assign array_update_71232[9] = add_71203 == 32'h0000_0009 ? array_update_71229 : array_update_71222[9];
  assign array_index_71234 = array_update_71230[add_71201 > 32'h0000_0009 ? 4'h9 : add_71201[3:0]];
  assign add_71235 = add_71225 + 32'h0000_0001;
  assign array_index_71236 = array_update_71232[add_71203 > 32'h0000_0009 ? 4'h9 : add_71203[3:0]];
  assign add_71237 = add_71227 + 32'h0000_0001;
  assign array_update_71238[0] = add_71235 == 32'h0000_0000 ? TestBlock__A_op23 : array_index_71234[0];
  assign array_update_71238[1] = add_71235 == 32'h0000_0001 ? TestBlock__A_op23 : array_index_71234[1];
  assign array_update_71238[2] = add_71235 == 32'h0000_0002 ? TestBlock__A_op23 : array_index_71234[2];
  assign array_update_71238[3] = add_71235 == 32'h0000_0003 ? TestBlock__A_op23 : array_index_71234[3];
  assign array_update_71238[4] = add_71235 == 32'h0000_0004 ? TestBlock__A_op23 : array_index_71234[4];
  assign array_update_71238[5] = add_71235 == 32'h0000_0005 ? TestBlock__A_op23 : array_index_71234[5];
  assign array_update_71238[6] = add_71235 == 32'h0000_0006 ? TestBlock__A_op23 : array_index_71234[6];
  assign array_update_71238[7] = add_71235 == 32'h0000_0007 ? TestBlock__A_op23 : array_index_71234[7];
  assign array_update_71238[8] = add_71235 == 32'h0000_0008 ? TestBlock__A_op23 : array_index_71234[8];
  assign array_update_71238[9] = add_71235 == 32'h0000_0009 ? TestBlock__A_op23 : array_index_71234[9];
  assign array_update_71239[0] = add_71237 == 32'h0000_0000 ? TestBlock__B_op23 : array_index_71236[0];
  assign array_update_71239[1] = add_71237 == 32'h0000_0001 ? TestBlock__B_op23 : array_index_71236[1];
  assign array_update_71239[2] = add_71237 == 32'h0000_0002 ? TestBlock__B_op23 : array_index_71236[2];
  assign array_update_71239[3] = add_71237 == 32'h0000_0003 ? TestBlock__B_op23 : array_index_71236[3];
  assign array_update_71239[4] = add_71237 == 32'h0000_0004 ? TestBlock__B_op23 : array_index_71236[4];
  assign array_update_71239[5] = add_71237 == 32'h0000_0005 ? TestBlock__B_op23 : array_index_71236[5];
  assign array_update_71239[6] = add_71237 == 32'h0000_0006 ? TestBlock__B_op23 : array_index_71236[6];
  assign array_update_71239[7] = add_71237 == 32'h0000_0007 ? TestBlock__B_op23 : array_index_71236[7];
  assign array_update_71239[8] = add_71237 == 32'h0000_0008 ? TestBlock__B_op23 : array_index_71236[8];
  assign array_update_71239[9] = add_71237 == 32'h0000_0009 ? TestBlock__B_op23 : array_index_71236[9];
  assign array_update_71240[0] = add_71201 == 32'h0000_0000 ? array_update_71238 : array_update_71230[0];
  assign array_update_71240[1] = add_71201 == 32'h0000_0001 ? array_update_71238 : array_update_71230[1];
  assign array_update_71240[2] = add_71201 == 32'h0000_0002 ? array_update_71238 : array_update_71230[2];
  assign array_update_71240[3] = add_71201 == 32'h0000_0003 ? array_update_71238 : array_update_71230[3];
  assign array_update_71240[4] = add_71201 == 32'h0000_0004 ? array_update_71238 : array_update_71230[4];
  assign array_update_71240[5] = add_71201 == 32'h0000_0005 ? array_update_71238 : array_update_71230[5];
  assign array_update_71240[6] = add_71201 == 32'h0000_0006 ? array_update_71238 : array_update_71230[6];
  assign array_update_71240[7] = add_71201 == 32'h0000_0007 ? array_update_71238 : array_update_71230[7];
  assign array_update_71240[8] = add_71201 == 32'h0000_0008 ? array_update_71238 : array_update_71230[8];
  assign array_update_71240[9] = add_71201 == 32'h0000_0009 ? array_update_71238 : array_update_71230[9];
  assign array_update_71242[0] = add_71203 == 32'h0000_0000 ? array_update_71239 : array_update_71232[0];
  assign array_update_71242[1] = add_71203 == 32'h0000_0001 ? array_update_71239 : array_update_71232[1];
  assign array_update_71242[2] = add_71203 == 32'h0000_0002 ? array_update_71239 : array_update_71232[2];
  assign array_update_71242[3] = add_71203 == 32'h0000_0003 ? array_update_71239 : array_update_71232[3];
  assign array_update_71242[4] = add_71203 == 32'h0000_0004 ? array_update_71239 : array_update_71232[4];
  assign array_update_71242[5] = add_71203 == 32'h0000_0005 ? array_update_71239 : array_update_71232[5];
  assign array_update_71242[6] = add_71203 == 32'h0000_0006 ? array_update_71239 : array_update_71232[6];
  assign array_update_71242[7] = add_71203 == 32'h0000_0007 ? array_update_71239 : array_update_71232[7];
  assign array_update_71242[8] = add_71203 == 32'h0000_0008 ? array_update_71239 : array_update_71232[8];
  assign array_update_71242[9] = add_71203 == 32'h0000_0009 ? array_update_71239 : array_update_71232[9];
  assign array_index_71244 = array_update_71240[add_71201 > 32'h0000_0009 ? 4'h9 : add_71201[3:0]];
  assign add_71245 = add_71235 + 32'h0000_0001;
  assign array_index_71246 = array_update_71242[add_71203 > 32'h0000_0009 ? 4'h9 : add_71203[3:0]];
  assign add_71247 = add_71237 + 32'h0000_0001;
  assign array_update_71248[0] = add_71245 == 32'h0000_0000 ? TestBlock__A_op24 : array_index_71244[0];
  assign array_update_71248[1] = add_71245 == 32'h0000_0001 ? TestBlock__A_op24 : array_index_71244[1];
  assign array_update_71248[2] = add_71245 == 32'h0000_0002 ? TestBlock__A_op24 : array_index_71244[2];
  assign array_update_71248[3] = add_71245 == 32'h0000_0003 ? TestBlock__A_op24 : array_index_71244[3];
  assign array_update_71248[4] = add_71245 == 32'h0000_0004 ? TestBlock__A_op24 : array_index_71244[4];
  assign array_update_71248[5] = add_71245 == 32'h0000_0005 ? TestBlock__A_op24 : array_index_71244[5];
  assign array_update_71248[6] = add_71245 == 32'h0000_0006 ? TestBlock__A_op24 : array_index_71244[6];
  assign array_update_71248[7] = add_71245 == 32'h0000_0007 ? TestBlock__A_op24 : array_index_71244[7];
  assign array_update_71248[8] = add_71245 == 32'h0000_0008 ? TestBlock__A_op24 : array_index_71244[8];
  assign array_update_71248[9] = add_71245 == 32'h0000_0009 ? TestBlock__A_op24 : array_index_71244[9];
  assign array_update_71249[0] = add_71247 == 32'h0000_0000 ? TestBlock__B_op24 : array_index_71246[0];
  assign array_update_71249[1] = add_71247 == 32'h0000_0001 ? TestBlock__B_op24 : array_index_71246[1];
  assign array_update_71249[2] = add_71247 == 32'h0000_0002 ? TestBlock__B_op24 : array_index_71246[2];
  assign array_update_71249[3] = add_71247 == 32'h0000_0003 ? TestBlock__B_op24 : array_index_71246[3];
  assign array_update_71249[4] = add_71247 == 32'h0000_0004 ? TestBlock__B_op24 : array_index_71246[4];
  assign array_update_71249[5] = add_71247 == 32'h0000_0005 ? TestBlock__B_op24 : array_index_71246[5];
  assign array_update_71249[6] = add_71247 == 32'h0000_0006 ? TestBlock__B_op24 : array_index_71246[6];
  assign array_update_71249[7] = add_71247 == 32'h0000_0007 ? TestBlock__B_op24 : array_index_71246[7];
  assign array_update_71249[8] = add_71247 == 32'h0000_0008 ? TestBlock__B_op24 : array_index_71246[8];
  assign array_update_71249[9] = add_71247 == 32'h0000_0009 ? TestBlock__B_op24 : array_index_71246[9];
  assign array_update_71250[0] = add_71201 == 32'h0000_0000 ? array_update_71248 : array_update_71240[0];
  assign array_update_71250[1] = add_71201 == 32'h0000_0001 ? array_update_71248 : array_update_71240[1];
  assign array_update_71250[2] = add_71201 == 32'h0000_0002 ? array_update_71248 : array_update_71240[2];
  assign array_update_71250[3] = add_71201 == 32'h0000_0003 ? array_update_71248 : array_update_71240[3];
  assign array_update_71250[4] = add_71201 == 32'h0000_0004 ? array_update_71248 : array_update_71240[4];
  assign array_update_71250[5] = add_71201 == 32'h0000_0005 ? array_update_71248 : array_update_71240[5];
  assign array_update_71250[6] = add_71201 == 32'h0000_0006 ? array_update_71248 : array_update_71240[6];
  assign array_update_71250[7] = add_71201 == 32'h0000_0007 ? array_update_71248 : array_update_71240[7];
  assign array_update_71250[8] = add_71201 == 32'h0000_0008 ? array_update_71248 : array_update_71240[8];
  assign array_update_71250[9] = add_71201 == 32'h0000_0009 ? array_update_71248 : array_update_71240[9];
  assign array_update_71252[0] = add_71203 == 32'h0000_0000 ? array_update_71249 : array_update_71242[0];
  assign array_update_71252[1] = add_71203 == 32'h0000_0001 ? array_update_71249 : array_update_71242[1];
  assign array_update_71252[2] = add_71203 == 32'h0000_0002 ? array_update_71249 : array_update_71242[2];
  assign array_update_71252[3] = add_71203 == 32'h0000_0003 ? array_update_71249 : array_update_71242[3];
  assign array_update_71252[4] = add_71203 == 32'h0000_0004 ? array_update_71249 : array_update_71242[4];
  assign array_update_71252[5] = add_71203 == 32'h0000_0005 ? array_update_71249 : array_update_71242[5];
  assign array_update_71252[6] = add_71203 == 32'h0000_0006 ? array_update_71249 : array_update_71242[6];
  assign array_update_71252[7] = add_71203 == 32'h0000_0007 ? array_update_71249 : array_update_71242[7];
  assign array_update_71252[8] = add_71203 == 32'h0000_0008 ? array_update_71249 : array_update_71242[8];
  assign array_update_71252[9] = add_71203 == 32'h0000_0009 ? array_update_71249 : array_update_71242[9];
  assign array_index_71254 = array_update_71250[add_71201 > 32'h0000_0009 ? 4'h9 : add_71201[3:0]];
  assign add_71255 = add_71245 + 32'h0000_0001;
  assign array_index_71256 = array_update_71252[add_71203 > 32'h0000_0009 ? 4'h9 : add_71203[3:0]];
  assign add_71257 = add_71247 + 32'h0000_0001;
  assign array_update_71258[0] = add_71255 == 32'h0000_0000 ? TestBlock__A_op25 : array_index_71254[0];
  assign array_update_71258[1] = add_71255 == 32'h0000_0001 ? TestBlock__A_op25 : array_index_71254[1];
  assign array_update_71258[2] = add_71255 == 32'h0000_0002 ? TestBlock__A_op25 : array_index_71254[2];
  assign array_update_71258[3] = add_71255 == 32'h0000_0003 ? TestBlock__A_op25 : array_index_71254[3];
  assign array_update_71258[4] = add_71255 == 32'h0000_0004 ? TestBlock__A_op25 : array_index_71254[4];
  assign array_update_71258[5] = add_71255 == 32'h0000_0005 ? TestBlock__A_op25 : array_index_71254[5];
  assign array_update_71258[6] = add_71255 == 32'h0000_0006 ? TestBlock__A_op25 : array_index_71254[6];
  assign array_update_71258[7] = add_71255 == 32'h0000_0007 ? TestBlock__A_op25 : array_index_71254[7];
  assign array_update_71258[8] = add_71255 == 32'h0000_0008 ? TestBlock__A_op25 : array_index_71254[8];
  assign array_update_71258[9] = add_71255 == 32'h0000_0009 ? TestBlock__A_op25 : array_index_71254[9];
  assign array_update_71259[0] = add_71257 == 32'h0000_0000 ? TestBlock__B_op25 : array_index_71256[0];
  assign array_update_71259[1] = add_71257 == 32'h0000_0001 ? TestBlock__B_op25 : array_index_71256[1];
  assign array_update_71259[2] = add_71257 == 32'h0000_0002 ? TestBlock__B_op25 : array_index_71256[2];
  assign array_update_71259[3] = add_71257 == 32'h0000_0003 ? TestBlock__B_op25 : array_index_71256[3];
  assign array_update_71259[4] = add_71257 == 32'h0000_0004 ? TestBlock__B_op25 : array_index_71256[4];
  assign array_update_71259[5] = add_71257 == 32'h0000_0005 ? TestBlock__B_op25 : array_index_71256[5];
  assign array_update_71259[6] = add_71257 == 32'h0000_0006 ? TestBlock__B_op25 : array_index_71256[6];
  assign array_update_71259[7] = add_71257 == 32'h0000_0007 ? TestBlock__B_op25 : array_index_71256[7];
  assign array_update_71259[8] = add_71257 == 32'h0000_0008 ? TestBlock__B_op25 : array_index_71256[8];
  assign array_update_71259[9] = add_71257 == 32'h0000_0009 ? TestBlock__B_op25 : array_index_71256[9];
  assign array_update_71260[0] = add_71201 == 32'h0000_0000 ? array_update_71258 : array_update_71250[0];
  assign array_update_71260[1] = add_71201 == 32'h0000_0001 ? array_update_71258 : array_update_71250[1];
  assign array_update_71260[2] = add_71201 == 32'h0000_0002 ? array_update_71258 : array_update_71250[2];
  assign array_update_71260[3] = add_71201 == 32'h0000_0003 ? array_update_71258 : array_update_71250[3];
  assign array_update_71260[4] = add_71201 == 32'h0000_0004 ? array_update_71258 : array_update_71250[4];
  assign array_update_71260[5] = add_71201 == 32'h0000_0005 ? array_update_71258 : array_update_71250[5];
  assign array_update_71260[6] = add_71201 == 32'h0000_0006 ? array_update_71258 : array_update_71250[6];
  assign array_update_71260[7] = add_71201 == 32'h0000_0007 ? array_update_71258 : array_update_71250[7];
  assign array_update_71260[8] = add_71201 == 32'h0000_0008 ? array_update_71258 : array_update_71250[8];
  assign array_update_71260[9] = add_71201 == 32'h0000_0009 ? array_update_71258 : array_update_71250[9];
  assign array_update_71262[0] = add_71203 == 32'h0000_0000 ? array_update_71259 : array_update_71252[0];
  assign array_update_71262[1] = add_71203 == 32'h0000_0001 ? array_update_71259 : array_update_71252[1];
  assign array_update_71262[2] = add_71203 == 32'h0000_0002 ? array_update_71259 : array_update_71252[2];
  assign array_update_71262[3] = add_71203 == 32'h0000_0003 ? array_update_71259 : array_update_71252[3];
  assign array_update_71262[4] = add_71203 == 32'h0000_0004 ? array_update_71259 : array_update_71252[4];
  assign array_update_71262[5] = add_71203 == 32'h0000_0005 ? array_update_71259 : array_update_71252[5];
  assign array_update_71262[6] = add_71203 == 32'h0000_0006 ? array_update_71259 : array_update_71252[6];
  assign array_update_71262[7] = add_71203 == 32'h0000_0007 ? array_update_71259 : array_update_71252[7];
  assign array_update_71262[8] = add_71203 == 32'h0000_0008 ? array_update_71259 : array_update_71252[8];
  assign array_update_71262[9] = add_71203 == 32'h0000_0009 ? array_update_71259 : array_update_71252[9];
  assign array_index_71264 = array_update_71260[add_71201 > 32'h0000_0009 ? 4'h9 : add_71201[3:0]];
  assign add_71265 = add_71255 + 32'h0000_0001;
  assign array_index_71266 = array_update_71262[add_71203 > 32'h0000_0009 ? 4'h9 : add_71203[3:0]];
  assign add_71267 = add_71257 + 32'h0000_0001;
  assign array_update_71268[0] = add_71265 == 32'h0000_0000 ? TestBlock__A_op26 : array_index_71264[0];
  assign array_update_71268[1] = add_71265 == 32'h0000_0001 ? TestBlock__A_op26 : array_index_71264[1];
  assign array_update_71268[2] = add_71265 == 32'h0000_0002 ? TestBlock__A_op26 : array_index_71264[2];
  assign array_update_71268[3] = add_71265 == 32'h0000_0003 ? TestBlock__A_op26 : array_index_71264[3];
  assign array_update_71268[4] = add_71265 == 32'h0000_0004 ? TestBlock__A_op26 : array_index_71264[4];
  assign array_update_71268[5] = add_71265 == 32'h0000_0005 ? TestBlock__A_op26 : array_index_71264[5];
  assign array_update_71268[6] = add_71265 == 32'h0000_0006 ? TestBlock__A_op26 : array_index_71264[6];
  assign array_update_71268[7] = add_71265 == 32'h0000_0007 ? TestBlock__A_op26 : array_index_71264[7];
  assign array_update_71268[8] = add_71265 == 32'h0000_0008 ? TestBlock__A_op26 : array_index_71264[8];
  assign array_update_71268[9] = add_71265 == 32'h0000_0009 ? TestBlock__A_op26 : array_index_71264[9];
  assign array_update_71269[0] = add_71267 == 32'h0000_0000 ? TestBlock__B_op26 : array_index_71266[0];
  assign array_update_71269[1] = add_71267 == 32'h0000_0001 ? TestBlock__B_op26 : array_index_71266[1];
  assign array_update_71269[2] = add_71267 == 32'h0000_0002 ? TestBlock__B_op26 : array_index_71266[2];
  assign array_update_71269[3] = add_71267 == 32'h0000_0003 ? TestBlock__B_op26 : array_index_71266[3];
  assign array_update_71269[4] = add_71267 == 32'h0000_0004 ? TestBlock__B_op26 : array_index_71266[4];
  assign array_update_71269[5] = add_71267 == 32'h0000_0005 ? TestBlock__B_op26 : array_index_71266[5];
  assign array_update_71269[6] = add_71267 == 32'h0000_0006 ? TestBlock__B_op26 : array_index_71266[6];
  assign array_update_71269[7] = add_71267 == 32'h0000_0007 ? TestBlock__B_op26 : array_index_71266[7];
  assign array_update_71269[8] = add_71267 == 32'h0000_0008 ? TestBlock__B_op26 : array_index_71266[8];
  assign array_update_71269[9] = add_71267 == 32'h0000_0009 ? TestBlock__B_op26 : array_index_71266[9];
  assign array_update_71270[0] = add_71201 == 32'h0000_0000 ? array_update_71268 : array_update_71260[0];
  assign array_update_71270[1] = add_71201 == 32'h0000_0001 ? array_update_71268 : array_update_71260[1];
  assign array_update_71270[2] = add_71201 == 32'h0000_0002 ? array_update_71268 : array_update_71260[2];
  assign array_update_71270[3] = add_71201 == 32'h0000_0003 ? array_update_71268 : array_update_71260[3];
  assign array_update_71270[4] = add_71201 == 32'h0000_0004 ? array_update_71268 : array_update_71260[4];
  assign array_update_71270[5] = add_71201 == 32'h0000_0005 ? array_update_71268 : array_update_71260[5];
  assign array_update_71270[6] = add_71201 == 32'h0000_0006 ? array_update_71268 : array_update_71260[6];
  assign array_update_71270[7] = add_71201 == 32'h0000_0007 ? array_update_71268 : array_update_71260[7];
  assign array_update_71270[8] = add_71201 == 32'h0000_0008 ? array_update_71268 : array_update_71260[8];
  assign array_update_71270[9] = add_71201 == 32'h0000_0009 ? array_update_71268 : array_update_71260[9];
  assign array_update_71272[0] = add_71203 == 32'h0000_0000 ? array_update_71269 : array_update_71262[0];
  assign array_update_71272[1] = add_71203 == 32'h0000_0001 ? array_update_71269 : array_update_71262[1];
  assign array_update_71272[2] = add_71203 == 32'h0000_0002 ? array_update_71269 : array_update_71262[2];
  assign array_update_71272[3] = add_71203 == 32'h0000_0003 ? array_update_71269 : array_update_71262[3];
  assign array_update_71272[4] = add_71203 == 32'h0000_0004 ? array_update_71269 : array_update_71262[4];
  assign array_update_71272[5] = add_71203 == 32'h0000_0005 ? array_update_71269 : array_update_71262[5];
  assign array_update_71272[6] = add_71203 == 32'h0000_0006 ? array_update_71269 : array_update_71262[6];
  assign array_update_71272[7] = add_71203 == 32'h0000_0007 ? array_update_71269 : array_update_71262[7];
  assign array_update_71272[8] = add_71203 == 32'h0000_0008 ? array_update_71269 : array_update_71262[8];
  assign array_update_71272[9] = add_71203 == 32'h0000_0009 ? array_update_71269 : array_update_71262[9];
  assign array_index_71274 = array_update_71270[add_71201 > 32'h0000_0009 ? 4'h9 : add_71201[3:0]];
  assign add_71275 = add_71265 + 32'h0000_0001;
  assign array_index_71276 = array_update_71272[add_71203 > 32'h0000_0009 ? 4'h9 : add_71203[3:0]];
  assign add_71277 = add_71267 + 32'h0000_0001;
  assign array_update_71278[0] = add_71275 == 32'h0000_0000 ? TestBlock__A_op27 : array_index_71274[0];
  assign array_update_71278[1] = add_71275 == 32'h0000_0001 ? TestBlock__A_op27 : array_index_71274[1];
  assign array_update_71278[2] = add_71275 == 32'h0000_0002 ? TestBlock__A_op27 : array_index_71274[2];
  assign array_update_71278[3] = add_71275 == 32'h0000_0003 ? TestBlock__A_op27 : array_index_71274[3];
  assign array_update_71278[4] = add_71275 == 32'h0000_0004 ? TestBlock__A_op27 : array_index_71274[4];
  assign array_update_71278[5] = add_71275 == 32'h0000_0005 ? TestBlock__A_op27 : array_index_71274[5];
  assign array_update_71278[6] = add_71275 == 32'h0000_0006 ? TestBlock__A_op27 : array_index_71274[6];
  assign array_update_71278[7] = add_71275 == 32'h0000_0007 ? TestBlock__A_op27 : array_index_71274[7];
  assign array_update_71278[8] = add_71275 == 32'h0000_0008 ? TestBlock__A_op27 : array_index_71274[8];
  assign array_update_71278[9] = add_71275 == 32'h0000_0009 ? TestBlock__A_op27 : array_index_71274[9];
  assign array_update_71279[0] = add_71277 == 32'h0000_0000 ? TestBlock__B_op27 : array_index_71276[0];
  assign array_update_71279[1] = add_71277 == 32'h0000_0001 ? TestBlock__B_op27 : array_index_71276[1];
  assign array_update_71279[2] = add_71277 == 32'h0000_0002 ? TestBlock__B_op27 : array_index_71276[2];
  assign array_update_71279[3] = add_71277 == 32'h0000_0003 ? TestBlock__B_op27 : array_index_71276[3];
  assign array_update_71279[4] = add_71277 == 32'h0000_0004 ? TestBlock__B_op27 : array_index_71276[4];
  assign array_update_71279[5] = add_71277 == 32'h0000_0005 ? TestBlock__B_op27 : array_index_71276[5];
  assign array_update_71279[6] = add_71277 == 32'h0000_0006 ? TestBlock__B_op27 : array_index_71276[6];
  assign array_update_71279[7] = add_71277 == 32'h0000_0007 ? TestBlock__B_op27 : array_index_71276[7];
  assign array_update_71279[8] = add_71277 == 32'h0000_0008 ? TestBlock__B_op27 : array_index_71276[8];
  assign array_update_71279[9] = add_71277 == 32'h0000_0009 ? TestBlock__B_op27 : array_index_71276[9];
  assign array_update_71280[0] = add_71201 == 32'h0000_0000 ? array_update_71278 : array_update_71270[0];
  assign array_update_71280[1] = add_71201 == 32'h0000_0001 ? array_update_71278 : array_update_71270[1];
  assign array_update_71280[2] = add_71201 == 32'h0000_0002 ? array_update_71278 : array_update_71270[2];
  assign array_update_71280[3] = add_71201 == 32'h0000_0003 ? array_update_71278 : array_update_71270[3];
  assign array_update_71280[4] = add_71201 == 32'h0000_0004 ? array_update_71278 : array_update_71270[4];
  assign array_update_71280[5] = add_71201 == 32'h0000_0005 ? array_update_71278 : array_update_71270[5];
  assign array_update_71280[6] = add_71201 == 32'h0000_0006 ? array_update_71278 : array_update_71270[6];
  assign array_update_71280[7] = add_71201 == 32'h0000_0007 ? array_update_71278 : array_update_71270[7];
  assign array_update_71280[8] = add_71201 == 32'h0000_0008 ? array_update_71278 : array_update_71270[8];
  assign array_update_71280[9] = add_71201 == 32'h0000_0009 ? array_update_71278 : array_update_71270[9];
  assign array_update_71282[0] = add_71203 == 32'h0000_0000 ? array_update_71279 : array_update_71272[0];
  assign array_update_71282[1] = add_71203 == 32'h0000_0001 ? array_update_71279 : array_update_71272[1];
  assign array_update_71282[2] = add_71203 == 32'h0000_0002 ? array_update_71279 : array_update_71272[2];
  assign array_update_71282[3] = add_71203 == 32'h0000_0003 ? array_update_71279 : array_update_71272[3];
  assign array_update_71282[4] = add_71203 == 32'h0000_0004 ? array_update_71279 : array_update_71272[4];
  assign array_update_71282[5] = add_71203 == 32'h0000_0005 ? array_update_71279 : array_update_71272[5];
  assign array_update_71282[6] = add_71203 == 32'h0000_0006 ? array_update_71279 : array_update_71272[6];
  assign array_update_71282[7] = add_71203 == 32'h0000_0007 ? array_update_71279 : array_update_71272[7];
  assign array_update_71282[8] = add_71203 == 32'h0000_0008 ? array_update_71279 : array_update_71272[8];
  assign array_update_71282[9] = add_71203 == 32'h0000_0009 ? array_update_71279 : array_update_71272[9];
  assign array_index_71284 = array_update_71280[add_71201 > 32'h0000_0009 ? 4'h9 : add_71201[3:0]];
  assign add_71285 = add_71275 + 32'h0000_0001;
  assign array_index_71286 = array_update_71282[add_71203 > 32'h0000_0009 ? 4'h9 : add_71203[3:0]];
  assign add_71287 = add_71277 + 32'h0000_0001;
  assign array_update_71288[0] = add_71285 == 32'h0000_0000 ? TestBlock__A_op28 : array_index_71284[0];
  assign array_update_71288[1] = add_71285 == 32'h0000_0001 ? TestBlock__A_op28 : array_index_71284[1];
  assign array_update_71288[2] = add_71285 == 32'h0000_0002 ? TestBlock__A_op28 : array_index_71284[2];
  assign array_update_71288[3] = add_71285 == 32'h0000_0003 ? TestBlock__A_op28 : array_index_71284[3];
  assign array_update_71288[4] = add_71285 == 32'h0000_0004 ? TestBlock__A_op28 : array_index_71284[4];
  assign array_update_71288[5] = add_71285 == 32'h0000_0005 ? TestBlock__A_op28 : array_index_71284[5];
  assign array_update_71288[6] = add_71285 == 32'h0000_0006 ? TestBlock__A_op28 : array_index_71284[6];
  assign array_update_71288[7] = add_71285 == 32'h0000_0007 ? TestBlock__A_op28 : array_index_71284[7];
  assign array_update_71288[8] = add_71285 == 32'h0000_0008 ? TestBlock__A_op28 : array_index_71284[8];
  assign array_update_71288[9] = add_71285 == 32'h0000_0009 ? TestBlock__A_op28 : array_index_71284[9];
  assign array_update_71289[0] = add_71287 == 32'h0000_0000 ? TestBlock__B_op28 : array_index_71286[0];
  assign array_update_71289[1] = add_71287 == 32'h0000_0001 ? TestBlock__B_op28 : array_index_71286[1];
  assign array_update_71289[2] = add_71287 == 32'h0000_0002 ? TestBlock__B_op28 : array_index_71286[2];
  assign array_update_71289[3] = add_71287 == 32'h0000_0003 ? TestBlock__B_op28 : array_index_71286[3];
  assign array_update_71289[4] = add_71287 == 32'h0000_0004 ? TestBlock__B_op28 : array_index_71286[4];
  assign array_update_71289[5] = add_71287 == 32'h0000_0005 ? TestBlock__B_op28 : array_index_71286[5];
  assign array_update_71289[6] = add_71287 == 32'h0000_0006 ? TestBlock__B_op28 : array_index_71286[6];
  assign array_update_71289[7] = add_71287 == 32'h0000_0007 ? TestBlock__B_op28 : array_index_71286[7];
  assign array_update_71289[8] = add_71287 == 32'h0000_0008 ? TestBlock__B_op28 : array_index_71286[8];
  assign array_update_71289[9] = add_71287 == 32'h0000_0009 ? TestBlock__B_op28 : array_index_71286[9];
  assign array_update_71290[0] = add_71201 == 32'h0000_0000 ? array_update_71288 : array_update_71280[0];
  assign array_update_71290[1] = add_71201 == 32'h0000_0001 ? array_update_71288 : array_update_71280[1];
  assign array_update_71290[2] = add_71201 == 32'h0000_0002 ? array_update_71288 : array_update_71280[2];
  assign array_update_71290[3] = add_71201 == 32'h0000_0003 ? array_update_71288 : array_update_71280[3];
  assign array_update_71290[4] = add_71201 == 32'h0000_0004 ? array_update_71288 : array_update_71280[4];
  assign array_update_71290[5] = add_71201 == 32'h0000_0005 ? array_update_71288 : array_update_71280[5];
  assign array_update_71290[6] = add_71201 == 32'h0000_0006 ? array_update_71288 : array_update_71280[6];
  assign array_update_71290[7] = add_71201 == 32'h0000_0007 ? array_update_71288 : array_update_71280[7];
  assign array_update_71290[8] = add_71201 == 32'h0000_0008 ? array_update_71288 : array_update_71280[8];
  assign array_update_71290[9] = add_71201 == 32'h0000_0009 ? array_update_71288 : array_update_71280[9];
  assign array_update_71292[0] = add_71203 == 32'h0000_0000 ? array_update_71289 : array_update_71282[0];
  assign array_update_71292[1] = add_71203 == 32'h0000_0001 ? array_update_71289 : array_update_71282[1];
  assign array_update_71292[2] = add_71203 == 32'h0000_0002 ? array_update_71289 : array_update_71282[2];
  assign array_update_71292[3] = add_71203 == 32'h0000_0003 ? array_update_71289 : array_update_71282[3];
  assign array_update_71292[4] = add_71203 == 32'h0000_0004 ? array_update_71289 : array_update_71282[4];
  assign array_update_71292[5] = add_71203 == 32'h0000_0005 ? array_update_71289 : array_update_71282[5];
  assign array_update_71292[6] = add_71203 == 32'h0000_0006 ? array_update_71289 : array_update_71282[6];
  assign array_update_71292[7] = add_71203 == 32'h0000_0007 ? array_update_71289 : array_update_71282[7];
  assign array_update_71292[8] = add_71203 == 32'h0000_0008 ? array_update_71289 : array_update_71282[8];
  assign array_update_71292[9] = add_71203 == 32'h0000_0009 ? array_update_71289 : array_update_71282[9];
  assign array_index_71294 = array_update_71290[add_71201 > 32'h0000_0009 ? 4'h9 : add_71201[3:0]];
  assign add_71295 = add_71285 + 32'h0000_0001;
  assign array_index_71296 = array_update_71292[add_71203 > 32'h0000_0009 ? 4'h9 : add_71203[3:0]];
  assign add_71297 = add_71287 + 32'h0000_0001;
  assign array_update_71298[0] = add_71295 == 32'h0000_0000 ? TestBlock__A_op29 : array_index_71294[0];
  assign array_update_71298[1] = add_71295 == 32'h0000_0001 ? TestBlock__A_op29 : array_index_71294[1];
  assign array_update_71298[2] = add_71295 == 32'h0000_0002 ? TestBlock__A_op29 : array_index_71294[2];
  assign array_update_71298[3] = add_71295 == 32'h0000_0003 ? TestBlock__A_op29 : array_index_71294[3];
  assign array_update_71298[4] = add_71295 == 32'h0000_0004 ? TestBlock__A_op29 : array_index_71294[4];
  assign array_update_71298[5] = add_71295 == 32'h0000_0005 ? TestBlock__A_op29 : array_index_71294[5];
  assign array_update_71298[6] = add_71295 == 32'h0000_0006 ? TestBlock__A_op29 : array_index_71294[6];
  assign array_update_71298[7] = add_71295 == 32'h0000_0007 ? TestBlock__A_op29 : array_index_71294[7];
  assign array_update_71298[8] = add_71295 == 32'h0000_0008 ? TestBlock__A_op29 : array_index_71294[8];
  assign array_update_71298[9] = add_71295 == 32'h0000_0009 ? TestBlock__A_op29 : array_index_71294[9];
  assign array_update_71300[0] = add_71297 == 32'h0000_0000 ? TestBlock__B_op29 : array_index_71296[0];
  assign array_update_71300[1] = add_71297 == 32'h0000_0001 ? TestBlock__B_op29 : array_index_71296[1];
  assign array_update_71300[2] = add_71297 == 32'h0000_0002 ? TestBlock__B_op29 : array_index_71296[2];
  assign array_update_71300[3] = add_71297 == 32'h0000_0003 ? TestBlock__B_op29 : array_index_71296[3];
  assign array_update_71300[4] = add_71297 == 32'h0000_0004 ? TestBlock__B_op29 : array_index_71296[4];
  assign array_update_71300[5] = add_71297 == 32'h0000_0005 ? TestBlock__B_op29 : array_index_71296[5];
  assign array_update_71300[6] = add_71297 == 32'h0000_0006 ? TestBlock__B_op29 : array_index_71296[6];
  assign array_update_71300[7] = add_71297 == 32'h0000_0007 ? TestBlock__B_op29 : array_index_71296[7];
  assign array_update_71300[8] = add_71297 == 32'h0000_0008 ? TestBlock__B_op29 : array_index_71296[8];
  assign array_update_71300[9] = add_71297 == 32'h0000_0009 ? TestBlock__B_op29 : array_index_71296[9];
  assign array_update_71302[0] = add_71201 == 32'h0000_0000 ? array_update_71298 : array_update_71290[0];
  assign array_update_71302[1] = add_71201 == 32'h0000_0001 ? array_update_71298 : array_update_71290[1];
  assign array_update_71302[2] = add_71201 == 32'h0000_0002 ? array_update_71298 : array_update_71290[2];
  assign array_update_71302[3] = add_71201 == 32'h0000_0003 ? array_update_71298 : array_update_71290[3];
  assign array_update_71302[4] = add_71201 == 32'h0000_0004 ? array_update_71298 : array_update_71290[4];
  assign array_update_71302[5] = add_71201 == 32'h0000_0005 ? array_update_71298 : array_update_71290[5];
  assign array_update_71302[6] = add_71201 == 32'h0000_0006 ? array_update_71298 : array_update_71290[6];
  assign array_update_71302[7] = add_71201 == 32'h0000_0007 ? array_update_71298 : array_update_71290[7];
  assign array_update_71302[8] = add_71201 == 32'h0000_0008 ? array_update_71298 : array_update_71290[8];
  assign array_update_71302[9] = add_71201 == 32'h0000_0009 ? array_update_71298 : array_update_71290[9];
  assign add_71303 = add_71201 + 32'h0000_0001;
  assign array_update_71304[0] = add_71203 == 32'h0000_0000 ? array_update_71300 : array_update_71292[0];
  assign array_update_71304[1] = add_71203 == 32'h0000_0001 ? array_update_71300 : array_update_71292[1];
  assign array_update_71304[2] = add_71203 == 32'h0000_0002 ? array_update_71300 : array_update_71292[2];
  assign array_update_71304[3] = add_71203 == 32'h0000_0003 ? array_update_71300 : array_update_71292[3];
  assign array_update_71304[4] = add_71203 == 32'h0000_0004 ? array_update_71300 : array_update_71292[4];
  assign array_update_71304[5] = add_71203 == 32'h0000_0005 ? array_update_71300 : array_update_71292[5];
  assign array_update_71304[6] = add_71203 == 32'h0000_0006 ? array_update_71300 : array_update_71292[6];
  assign array_update_71304[7] = add_71203 == 32'h0000_0007 ? array_update_71300 : array_update_71292[7];
  assign array_update_71304[8] = add_71203 == 32'h0000_0008 ? array_update_71300 : array_update_71292[8];
  assign array_update_71304[9] = add_71203 == 32'h0000_0009 ? array_update_71300 : array_update_71292[9];
  assign add_71305 = add_71203 + 32'h0000_0001;
  assign array_index_71306 = array_update_71302[add_71303 > 32'h0000_0009 ? 4'h9 : add_71303[3:0]];
  assign literal_71307 = 32'h0000_0000;
  assign array_index_71308 = array_update_71304[add_71305 > 32'h0000_0009 ? 4'h9 : add_71305[3:0]];
  assign literal_71309 = 32'h0000_0000;
  assign array_update_71310[0] = literal_71307 == 32'h0000_0000 ? TestBlock__A_op30 : array_index_71306[0];
  assign array_update_71310[1] = literal_71307 == 32'h0000_0001 ? TestBlock__A_op30 : array_index_71306[1];
  assign array_update_71310[2] = literal_71307 == 32'h0000_0002 ? TestBlock__A_op30 : array_index_71306[2];
  assign array_update_71310[3] = literal_71307 == 32'h0000_0003 ? TestBlock__A_op30 : array_index_71306[3];
  assign array_update_71310[4] = literal_71307 == 32'h0000_0004 ? TestBlock__A_op30 : array_index_71306[4];
  assign array_update_71310[5] = literal_71307 == 32'h0000_0005 ? TestBlock__A_op30 : array_index_71306[5];
  assign array_update_71310[6] = literal_71307 == 32'h0000_0006 ? TestBlock__A_op30 : array_index_71306[6];
  assign array_update_71310[7] = literal_71307 == 32'h0000_0007 ? TestBlock__A_op30 : array_index_71306[7];
  assign array_update_71310[8] = literal_71307 == 32'h0000_0008 ? TestBlock__A_op30 : array_index_71306[8];
  assign array_update_71310[9] = literal_71307 == 32'h0000_0009 ? TestBlock__A_op30 : array_index_71306[9];
  assign array_update_71311[0] = literal_71309 == 32'h0000_0000 ? TestBlock__B_op30 : array_index_71308[0];
  assign array_update_71311[1] = literal_71309 == 32'h0000_0001 ? TestBlock__B_op30 : array_index_71308[1];
  assign array_update_71311[2] = literal_71309 == 32'h0000_0002 ? TestBlock__B_op30 : array_index_71308[2];
  assign array_update_71311[3] = literal_71309 == 32'h0000_0003 ? TestBlock__B_op30 : array_index_71308[3];
  assign array_update_71311[4] = literal_71309 == 32'h0000_0004 ? TestBlock__B_op30 : array_index_71308[4];
  assign array_update_71311[5] = literal_71309 == 32'h0000_0005 ? TestBlock__B_op30 : array_index_71308[5];
  assign array_update_71311[6] = literal_71309 == 32'h0000_0006 ? TestBlock__B_op30 : array_index_71308[6];
  assign array_update_71311[7] = literal_71309 == 32'h0000_0007 ? TestBlock__B_op30 : array_index_71308[7];
  assign array_update_71311[8] = literal_71309 == 32'h0000_0008 ? TestBlock__B_op30 : array_index_71308[8];
  assign array_update_71311[9] = literal_71309 == 32'h0000_0009 ? TestBlock__B_op30 : array_index_71308[9];
  assign array_update_71312[0] = add_71303 == 32'h0000_0000 ? array_update_71310 : array_update_71302[0];
  assign array_update_71312[1] = add_71303 == 32'h0000_0001 ? array_update_71310 : array_update_71302[1];
  assign array_update_71312[2] = add_71303 == 32'h0000_0002 ? array_update_71310 : array_update_71302[2];
  assign array_update_71312[3] = add_71303 == 32'h0000_0003 ? array_update_71310 : array_update_71302[3];
  assign array_update_71312[4] = add_71303 == 32'h0000_0004 ? array_update_71310 : array_update_71302[4];
  assign array_update_71312[5] = add_71303 == 32'h0000_0005 ? array_update_71310 : array_update_71302[5];
  assign array_update_71312[6] = add_71303 == 32'h0000_0006 ? array_update_71310 : array_update_71302[6];
  assign array_update_71312[7] = add_71303 == 32'h0000_0007 ? array_update_71310 : array_update_71302[7];
  assign array_update_71312[8] = add_71303 == 32'h0000_0008 ? array_update_71310 : array_update_71302[8];
  assign array_update_71312[9] = add_71303 == 32'h0000_0009 ? array_update_71310 : array_update_71302[9];
  assign array_update_71314[0] = add_71305 == 32'h0000_0000 ? array_update_71311 : array_update_71304[0];
  assign array_update_71314[1] = add_71305 == 32'h0000_0001 ? array_update_71311 : array_update_71304[1];
  assign array_update_71314[2] = add_71305 == 32'h0000_0002 ? array_update_71311 : array_update_71304[2];
  assign array_update_71314[3] = add_71305 == 32'h0000_0003 ? array_update_71311 : array_update_71304[3];
  assign array_update_71314[4] = add_71305 == 32'h0000_0004 ? array_update_71311 : array_update_71304[4];
  assign array_update_71314[5] = add_71305 == 32'h0000_0005 ? array_update_71311 : array_update_71304[5];
  assign array_update_71314[6] = add_71305 == 32'h0000_0006 ? array_update_71311 : array_update_71304[6];
  assign array_update_71314[7] = add_71305 == 32'h0000_0007 ? array_update_71311 : array_update_71304[7];
  assign array_update_71314[8] = add_71305 == 32'h0000_0008 ? array_update_71311 : array_update_71304[8];
  assign array_update_71314[9] = add_71305 == 32'h0000_0009 ? array_update_71311 : array_update_71304[9];
  assign array_index_71316 = array_update_71312[add_71303 > 32'h0000_0009 ? 4'h9 : add_71303[3:0]];
  assign add_71317 = literal_71307 + 32'h0000_0001;
  assign array_index_71318 = array_update_71314[add_71305 > 32'h0000_0009 ? 4'h9 : add_71305[3:0]];
  assign add_71319 = literal_71309 + 32'h0000_0001;
  assign array_update_71320[0] = add_71317 == 32'h0000_0000 ? TestBlock__A_op31 : array_index_71316[0];
  assign array_update_71320[1] = add_71317 == 32'h0000_0001 ? TestBlock__A_op31 : array_index_71316[1];
  assign array_update_71320[2] = add_71317 == 32'h0000_0002 ? TestBlock__A_op31 : array_index_71316[2];
  assign array_update_71320[3] = add_71317 == 32'h0000_0003 ? TestBlock__A_op31 : array_index_71316[3];
  assign array_update_71320[4] = add_71317 == 32'h0000_0004 ? TestBlock__A_op31 : array_index_71316[4];
  assign array_update_71320[5] = add_71317 == 32'h0000_0005 ? TestBlock__A_op31 : array_index_71316[5];
  assign array_update_71320[6] = add_71317 == 32'h0000_0006 ? TestBlock__A_op31 : array_index_71316[6];
  assign array_update_71320[7] = add_71317 == 32'h0000_0007 ? TestBlock__A_op31 : array_index_71316[7];
  assign array_update_71320[8] = add_71317 == 32'h0000_0008 ? TestBlock__A_op31 : array_index_71316[8];
  assign array_update_71320[9] = add_71317 == 32'h0000_0009 ? TestBlock__A_op31 : array_index_71316[9];
  assign array_update_71321[0] = add_71319 == 32'h0000_0000 ? TestBlock__B_op31 : array_index_71318[0];
  assign array_update_71321[1] = add_71319 == 32'h0000_0001 ? TestBlock__B_op31 : array_index_71318[1];
  assign array_update_71321[2] = add_71319 == 32'h0000_0002 ? TestBlock__B_op31 : array_index_71318[2];
  assign array_update_71321[3] = add_71319 == 32'h0000_0003 ? TestBlock__B_op31 : array_index_71318[3];
  assign array_update_71321[4] = add_71319 == 32'h0000_0004 ? TestBlock__B_op31 : array_index_71318[4];
  assign array_update_71321[5] = add_71319 == 32'h0000_0005 ? TestBlock__B_op31 : array_index_71318[5];
  assign array_update_71321[6] = add_71319 == 32'h0000_0006 ? TestBlock__B_op31 : array_index_71318[6];
  assign array_update_71321[7] = add_71319 == 32'h0000_0007 ? TestBlock__B_op31 : array_index_71318[7];
  assign array_update_71321[8] = add_71319 == 32'h0000_0008 ? TestBlock__B_op31 : array_index_71318[8];
  assign array_update_71321[9] = add_71319 == 32'h0000_0009 ? TestBlock__B_op31 : array_index_71318[9];
  assign array_update_71322[0] = add_71303 == 32'h0000_0000 ? array_update_71320 : array_update_71312[0];
  assign array_update_71322[1] = add_71303 == 32'h0000_0001 ? array_update_71320 : array_update_71312[1];
  assign array_update_71322[2] = add_71303 == 32'h0000_0002 ? array_update_71320 : array_update_71312[2];
  assign array_update_71322[3] = add_71303 == 32'h0000_0003 ? array_update_71320 : array_update_71312[3];
  assign array_update_71322[4] = add_71303 == 32'h0000_0004 ? array_update_71320 : array_update_71312[4];
  assign array_update_71322[5] = add_71303 == 32'h0000_0005 ? array_update_71320 : array_update_71312[5];
  assign array_update_71322[6] = add_71303 == 32'h0000_0006 ? array_update_71320 : array_update_71312[6];
  assign array_update_71322[7] = add_71303 == 32'h0000_0007 ? array_update_71320 : array_update_71312[7];
  assign array_update_71322[8] = add_71303 == 32'h0000_0008 ? array_update_71320 : array_update_71312[8];
  assign array_update_71322[9] = add_71303 == 32'h0000_0009 ? array_update_71320 : array_update_71312[9];
  assign array_update_71324[0] = add_71305 == 32'h0000_0000 ? array_update_71321 : array_update_71314[0];
  assign array_update_71324[1] = add_71305 == 32'h0000_0001 ? array_update_71321 : array_update_71314[1];
  assign array_update_71324[2] = add_71305 == 32'h0000_0002 ? array_update_71321 : array_update_71314[2];
  assign array_update_71324[3] = add_71305 == 32'h0000_0003 ? array_update_71321 : array_update_71314[3];
  assign array_update_71324[4] = add_71305 == 32'h0000_0004 ? array_update_71321 : array_update_71314[4];
  assign array_update_71324[5] = add_71305 == 32'h0000_0005 ? array_update_71321 : array_update_71314[5];
  assign array_update_71324[6] = add_71305 == 32'h0000_0006 ? array_update_71321 : array_update_71314[6];
  assign array_update_71324[7] = add_71305 == 32'h0000_0007 ? array_update_71321 : array_update_71314[7];
  assign array_update_71324[8] = add_71305 == 32'h0000_0008 ? array_update_71321 : array_update_71314[8];
  assign array_update_71324[9] = add_71305 == 32'h0000_0009 ? array_update_71321 : array_update_71314[9];
  assign array_index_71326 = array_update_71322[add_71303 > 32'h0000_0009 ? 4'h9 : add_71303[3:0]];
  assign add_71327 = add_71317 + 32'h0000_0001;
  assign array_index_71328 = array_update_71324[add_71305 > 32'h0000_0009 ? 4'h9 : add_71305[3:0]];
  assign add_71329 = add_71319 + 32'h0000_0001;
  assign array_update_71330[0] = add_71327 == 32'h0000_0000 ? TestBlock__A_op32 : array_index_71326[0];
  assign array_update_71330[1] = add_71327 == 32'h0000_0001 ? TestBlock__A_op32 : array_index_71326[1];
  assign array_update_71330[2] = add_71327 == 32'h0000_0002 ? TestBlock__A_op32 : array_index_71326[2];
  assign array_update_71330[3] = add_71327 == 32'h0000_0003 ? TestBlock__A_op32 : array_index_71326[3];
  assign array_update_71330[4] = add_71327 == 32'h0000_0004 ? TestBlock__A_op32 : array_index_71326[4];
  assign array_update_71330[5] = add_71327 == 32'h0000_0005 ? TestBlock__A_op32 : array_index_71326[5];
  assign array_update_71330[6] = add_71327 == 32'h0000_0006 ? TestBlock__A_op32 : array_index_71326[6];
  assign array_update_71330[7] = add_71327 == 32'h0000_0007 ? TestBlock__A_op32 : array_index_71326[7];
  assign array_update_71330[8] = add_71327 == 32'h0000_0008 ? TestBlock__A_op32 : array_index_71326[8];
  assign array_update_71330[9] = add_71327 == 32'h0000_0009 ? TestBlock__A_op32 : array_index_71326[9];
  assign array_update_71331[0] = add_71329 == 32'h0000_0000 ? TestBlock__B_op32 : array_index_71328[0];
  assign array_update_71331[1] = add_71329 == 32'h0000_0001 ? TestBlock__B_op32 : array_index_71328[1];
  assign array_update_71331[2] = add_71329 == 32'h0000_0002 ? TestBlock__B_op32 : array_index_71328[2];
  assign array_update_71331[3] = add_71329 == 32'h0000_0003 ? TestBlock__B_op32 : array_index_71328[3];
  assign array_update_71331[4] = add_71329 == 32'h0000_0004 ? TestBlock__B_op32 : array_index_71328[4];
  assign array_update_71331[5] = add_71329 == 32'h0000_0005 ? TestBlock__B_op32 : array_index_71328[5];
  assign array_update_71331[6] = add_71329 == 32'h0000_0006 ? TestBlock__B_op32 : array_index_71328[6];
  assign array_update_71331[7] = add_71329 == 32'h0000_0007 ? TestBlock__B_op32 : array_index_71328[7];
  assign array_update_71331[8] = add_71329 == 32'h0000_0008 ? TestBlock__B_op32 : array_index_71328[8];
  assign array_update_71331[9] = add_71329 == 32'h0000_0009 ? TestBlock__B_op32 : array_index_71328[9];
  assign array_update_71332[0] = add_71303 == 32'h0000_0000 ? array_update_71330 : array_update_71322[0];
  assign array_update_71332[1] = add_71303 == 32'h0000_0001 ? array_update_71330 : array_update_71322[1];
  assign array_update_71332[2] = add_71303 == 32'h0000_0002 ? array_update_71330 : array_update_71322[2];
  assign array_update_71332[3] = add_71303 == 32'h0000_0003 ? array_update_71330 : array_update_71322[3];
  assign array_update_71332[4] = add_71303 == 32'h0000_0004 ? array_update_71330 : array_update_71322[4];
  assign array_update_71332[5] = add_71303 == 32'h0000_0005 ? array_update_71330 : array_update_71322[5];
  assign array_update_71332[6] = add_71303 == 32'h0000_0006 ? array_update_71330 : array_update_71322[6];
  assign array_update_71332[7] = add_71303 == 32'h0000_0007 ? array_update_71330 : array_update_71322[7];
  assign array_update_71332[8] = add_71303 == 32'h0000_0008 ? array_update_71330 : array_update_71322[8];
  assign array_update_71332[9] = add_71303 == 32'h0000_0009 ? array_update_71330 : array_update_71322[9];
  assign array_update_71334[0] = add_71305 == 32'h0000_0000 ? array_update_71331 : array_update_71324[0];
  assign array_update_71334[1] = add_71305 == 32'h0000_0001 ? array_update_71331 : array_update_71324[1];
  assign array_update_71334[2] = add_71305 == 32'h0000_0002 ? array_update_71331 : array_update_71324[2];
  assign array_update_71334[3] = add_71305 == 32'h0000_0003 ? array_update_71331 : array_update_71324[3];
  assign array_update_71334[4] = add_71305 == 32'h0000_0004 ? array_update_71331 : array_update_71324[4];
  assign array_update_71334[5] = add_71305 == 32'h0000_0005 ? array_update_71331 : array_update_71324[5];
  assign array_update_71334[6] = add_71305 == 32'h0000_0006 ? array_update_71331 : array_update_71324[6];
  assign array_update_71334[7] = add_71305 == 32'h0000_0007 ? array_update_71331 : array_update_71324[7];
  assign array_update_71334[8] = add_71305 == 32'h0000_0008 ? array_update_71331 : array_update_71324[8];
  assign array_update_71334[9] = add_71305 == 32'h0000_0009 ? array_update_71331 : array_update_71324[9];
  assign array_index_71336 = array_update_71332[add_71303 > 32'h0000_0009 ? 4'h9 : add_71303[3:0]];
  assign add_71337 = add_71327 + 32'h0000_0001;
  assign array_index_71338 = array_update_71334[add_71305 > 32'h0000_0009 ? 4'h9 : add_71305[3:0]];
  assign add_71339 = add_71329 + 32'h0000_0001;
  assign array_update_71340[0] = add_71337 == 32'h0000_0000 ? TestBlock__A_op33 : array_index_71336[0];
  assign array_update_71340[1] = add_71337 == 32'h0000_0001 ? TestBlock__A_op33 : array_index_71336[1];
  assign array_update_71340[2] = add_71337 == 32'h0000_0002 ? TestBlock__A_op33 : array_index_71336[2];
  assign array_update_71340[3] = add_71337 == 32'h0000_0003 ? TestBlock__A_op33 : array_index_71336[3];
  assign array_update_71340[4] = add_71337 == 32'h0000_0004 ? TestBlock__A_op33 : array_index_71336[4];
  assign array_update_71340[5] = add_71337 == 32'h0000_0005 ? TestBlock__A_op33 : array_index_71336[5];
  assign array_update_71340[6] = add_71337 == 32'h0000_0006 ? TestBlock__A_op33 : array_index_71336[6];
  assign array_update_71340[7] = add_71337 == 32'h0000_0007 ? TestBlock__A_op33 : array_index_71336[7];
  assign array_update_71340[8] = add_71337 == 32'h0000_0008 ? TestBlock__A_op33 : array_index_71336[8];
  assign array_update_71340[9] = add_71337 == 32'h0000_0009 ? TestBlock__A_op33 : array_index_71336[9];
  assign array_update_71341[0] = add_71339 == 32'h0000_0000 ? TestBlock__B_op33 : array_index_71338[0];
  assign array_update_71341[1] = add_71339 == 32'h0000_0001 ? TestBlock__B_op33 : array_index_71338[1];
  assign array_update_71341[2] = add_71339 == 32'h0000_0002 ? TestBlock__B_op33 : array_index_71338[2];
  assign array_update_71341[3] = add_71339 == 32'h0000_0003 ? TestBlock__B_op33 : array_index_71338[3];
  assign array_update_71341[4] = add_71339 == 32'h0000_0004 ? TestBlock__B_op33 : array_index_71338[4];
  assign array_update_71341[5] = add_71339 == 32'h0000_0005 ? TestBlock__B_op33 : array_index_71338[5];
  assign array_update_71341[6] = add_71339 == 32'h0000_0006 ? TestBlock__B_op33 : array_index_71338[6];
  assign array_update_71341[7] = add_71339 == 32'h0000_0007 ? TestBlock__B_op33 : array_index_71338[7];
  assign array_update_71341[8] = add_71339 == 32'h0000_0008 ? TestBlock__B_op33 : array_index_71338[8];
  assign array_update_71341[9] = add_71339 == 32'h0000_0009 ? TestBlock__B_op33 : array_index_71338[9];
  assign array_update_71342[0] = add_71303 == 32'h0000_0000 ? array_update_71340 : array_update_71332[0];
  assign array_update_71342[1] = add_71303 == 32'h0000_0001 ? array_update_71340 : array_update_71332[1];
  assign array_update_71342[2] = add_71303 == 32'h0000_0002 ? array_update_71340 : array_update_71332[2];
  assign array_update_71342[3] = add_71303 == 32'h0000_0003 ? array_update_71340 : array_update_71332[3];
  assign array_update_71342[4] = add_71303 == 32'h0000_0004 ? array_update_71340 : array_update_71332[4];
  assign array_update_71342[5] = add_71303 == 32'h0000_0005 ? array_update_71340 : array_update_71332[5];
  assign array_update_71342[6] = add_71303 == 32'h0000_0006 ? array_update_71340 : array_update_71332[6];
  assign array_update_71342[7] = add_71303 == 32'h0000_0007 ? array_update_71340 : array_update_71332[7];
  assign array_update_71342[8] = add_71303 == 32'h0000_0008 ? array_update_71340 : array_update_71332[8];
  assign array_update_71342[9] = add_71303 == 32'h0000_0009 ? array_update_71340 : array_update_71332[9];
  assign array_update_71344[0] = add_71305 == 32'h0000_0000 ? array_update_71341 : array_update_71334[0];
  assign array_update_71344[1] = add_71305 == 32'h0000_0001 ? array_update_71341 : array_update_71334[1];
  assign array_update_71344[2] = add_71305 == 32'h0000_0002 ? array_update_71341 : array_update_71334[2];
  assign array_update_71344[3] = add_71305 == 32'h0000_0003 ? array_update_71341 : array_update_71334[3];
  assign array_update_71344[4] = add_71305 == 32'h0000_0004 ? array_update_71341 : array_update_71334[4];
  assign array_update_71344[5] = add_71305 == 32'h0000_0005 ? array_update_71341 : array_update_71334[5];
  assign array_update_71344[6] = add_71305 == 32'h0000_0006 ? array_update_71341 : array_update_71334[6];
  assign array_update_71344[7] = add_71305 == 32'h0000_0007 ? array_update_71341 : array_update_71334[7];
  assign array_update_71344[8] = add_71305 == 32'h0000_0008 ? array_update_71341 : array_update_71334[8];
  assign array_update_71344[9] = add_71305 == 32'h0000_0009 ? array_update_71341 : array_update_71334[9];
  assign array_index_71346 = array_update_71342[add_71303 > 32'h0000_0009 ? 4'h9 : add_71303[3:0]];
  assign add_71347 = add_71337 + 32'h0000_0001;
  assign array_index_71348 = array_update_71344[add_71305 > 32'h0000_0009 ? 4'h9 : add_71305[3:0]];
  assign add_71349 = add_71339 + 32'h0000_0001;
  assign array_update_71350[0] = add_71347 == 32'h0000_0000 ? TestBlock__A_op34 : array_index_71346[0];
  assign array_update_71350[1] = add_71347 == 32'h0000_0001 ? TestBlock__A_op34 : array_index_71346[1];
  assign array_update_71350[2] = add_71347 == 32'h0000_0002 ? TestBlock__A_op34 : array_index_71346[2];
  assign array_update_71350[3] = add_71347 == 32'h0000_0003 ? TestBlock__A_op34 : array_index_71346[3];
  assign array_update_71350[4] = add_71347 == 32'h0000_0004 ? TestBlock__A_op34 : array_index_71346[4];
  assign array_update_71350[5] = add_71347 == 32'h0000_0005 ? TestBlock__A_op34 : array_index_71346[5];
  assign array_update_71350[6] = add_71347 == 32'h0000_0006 ? TestBlock__A_op34 : array_index_71346[6];
  assign array_update_71350[7] = add_71347 == 32'h0000_0007 ? TestBlock__A_op34 : array_index_71346[7];
  assign array_update_71350[8] = add_71347 == 32'h0000_0008 ? TestBlock__A_op34 : array_index_71346[8];
  assign array_update_71350[9] = add_71347 == 32'h0000_0009 ? TestBlock__A_op34 : array_index_71346[9];
  assign array_update_71351[0] = add_71349 == 32'h0000_0000 ? TestBlock__B_op34 : array_index_71348[0];
  assign array_update_71351[1] = add_71349 == 32'h0000_0001 ? TestBlock__B_op34 : array_index_71348[1];
  assign array_update_71351[2] = add_71349 == 32'h0000_0002 ? TestBlock__B_op34 : array_index_71348[2];
  assign array_update_71351[3] = add_71349 == 32'h0000_0003 ? TestBlock__B_op34 : array_index_71348[3];
  assign array_update_71351[4] = add_71349 == 32'h0000_0004 ? TestBlock__B_op34 : array_index_71348[4];
  assign array_update_71351[5] = add_71349 == 32'h0000_0005 ? TestBlock__B_op34 : array_index_71348[5];
  assign array_update_71351[6] = add_71349 == 32'h0000_0006 ? TestBlock__B_op34 : array_index_71348[6];
  assign array_update_71351[7] = add_71349 == 32'h0000_0007 ? TestBlock__B_op34 : array_index_71348[7];
  assign array_update_71351[8] = add_71349 == 32'h0000_0008 ? TestBlock__B_op34 : array_index_71348[8];
  assign array_update_71351[9] = add_71349 == 32'h0000_0009 ? TestBlock__B_op34 : array_index_71348[9];
  assign array_update_71352[0] = add_71303 == 32'h0000_0000 ? array_update_71350 : array_update_71342[0];
  assign array_update_71352[1] = add_71303 == 32'h0000_0001 ? array_update_71350 : array_update_71342[1];
  assign array_update_71352[2] = add_71303 == 32'h0000_0002 ? array_update_71350 : array_update_71342[2];
  assign array_update_71352[3] = add_71303 == 32'h0000_0003 ? array_update_71350 : array_update_71342[3];
  assign array_update_71352[4] = add_71303 == 32'h0000_0004 ? array_update_71350 : array_update_71342[4];
  assign array_update_71352[5] = add_71303 == 32'h0000_0005 ? array_update_71350 : array_update_71342[5];
  assign array_update_71352[6] = add_71303 == 32'h0000_0006 ? array_update_71350 : array_update_71342[6];
  assign array_update_71352[7] = add_71303 == 32'h0000_0007 ? array_update_71350 : array_update_71342[7];
  assign array_update_71352[8] = add_71303 == 32'h0000_0008 ? array_update_71350 : array_update_71342[8];
  assign array_update_71352[9] = add_71303 == 32'h0000_0009 ? array_update_71350 : array_update_71342[9];
  assign array_update_71354[0] = add_71305 == 32'h0000_0000 ? array_update_71351 : array_update_71344[0];
  assign array_update_71354[1] = add_71305 == 32'h0000_0001 ? array_update_71351 : array_update_71344[1];
  assign array_update_71354[2] = add_71305 == 32'h0000_0002 ? array_update_71351 : array_update_71344[2];
  assign array_update_71354[3] = add_71305 == 32'h0000_0003 ? array_update_71351 : array_update_71344[3];
  assign array_update_71354[4] = add_71305 == 32'h0000_0004 ? array_update_71351 : array_update_71344[4];
  assign array_update_71354[5] = add_71305 == 32'h0000_0005 ? array_update_71351 : array_update_71344[5];
  assign array_update_71354[6] = add_71305 == 32'h0000_0006 ? array_update_71351 : array_update_71344[6];
  assign array_update_71354[7] = add_71305 == 32'h0000_0007 ? array_update_71351 : array_update_71344[7];
  assign array_update_71354[8] = add_71305 == 32'h0000_0008 ? array_update_71351 : array_update_71344[8];
  assign array_update_71354[9] = add_71305 == 32'h0000_0009 ? array_update_71351 : array_update_71344[9];
  assign array_index_71356 = array_update_71352[add_71303 > 32'h0000_0009 ? 4'h9 : add_71303[3:0]];
  assign add_71357 = add_71347 + 32'h0000_0001;
  assign array_index_71358 = array_update_71354[add_71305 > 32'h0000_0009 ? 4'h9 : add_71305[3:0]];
  assign add_71359 = add_71349 + 32'h0000_0001;
  assign array_update_71360[0] = add_71357 == 32'h0000_0000 ? TestBlock__A_op35 : array_index_71356[0];
  assign array_update_71360[1] = add_71357 == 32'h0000_0001 ? TestBlock__A_op35 : array_index_71356[1];
  assign array_update_71360[2] = add_71357 == 32'h0000_0002 ? TestBlock__A_op35 : array_index_71356[2];
  assign array_update_71360[3] = add_71357 == 32'h0000_0003 ? TestBlock__A_op35 : array_index_71356[3];
  assign array_update_71360[4] = add_71357 == 32'h0000_0004 ? TestBlock__A_op35 : array_index_71356[4];
  assign array_update_71360[5] = add_71357 == 32'h0000_0005 ? TestBlock__A_op35 : array_index_71356[5];
  assign array_update_71360[6] = add_71357 == 32'h0000_0006 ? TestBlock__A_op35 : array_index_71356[6];
  assign array_update_71360[7] = add_71357 == 32'h0000_0007 ? TestBlock__A_op35 : array_index_71356[7];
  assign array_update_71360[8] = add_71357 == 32'h0000_0008 ? TestBlock__A_op35 : array_index_71356[8];
  assign array_update_71360[9] = add_71357 == 32'h0000_0009 ? TestBlock__A_op35 : array_index_71356[9];
  assign array_update_71361[0] = add_71359 == 32'h0000_0000 ? TestBlock__B_op35 : array_index_71358[0];
  assign array_update_71361[1] = add_71359 == 32'h0000_0001 ? TestBlock__B_op35 : array_index_71358[1];
  assign array_update_71361[2] = add_71359 == 32'h0000_0002 ? TestBlock__B_op35 : array_index_71358[2];
  assign array_update_71361[3] = add_71359 == 32'h0000_0003 ? TestBlock__B_op35 : array_index_71358[3];
  assign array_update_71361[4] = add_71359 == 32'h0000_0004 ? TestBlock__B_op35 : array_index_71358[4];
  assign array_update_71361[5] = add_71359 == 32'h0000_0005 ? TestBlock__B_op35 : array_index_71358[5];
  assign array_update_71361[6] = add_71359 == 32'h0000_0006 ? TestBlock__B_op35 : array_index_71358[6];
  assign array_update_71361[7] = add_71359 == 32'h0000_0007 ? TestBlock__B_op35 : array_index_71358[7];
  assign array_update_71361[8] = add_71359 == 32'h0000_0008 ? TestBlock__B_op35 : array_index_71358[8];
  assign array_update_71361[9] = add_71359 == 32'h0000_0009 ? TestBlock__B_op35 : array_index_71358[9];
  assign array_update_71362[0] = add_71303 == 32'h0000_0000 ? array_update_71360 : array_update_71352[0];
  assign array_update_71362[1] = add_71303 == 32'h0000_0001 ? array_update_71360 : array_update_71352[1];
  assign array_update_71362[2] = add_71303 == 32'h0000_0002 ? array_update_71360 : array_update_71352[2];
  assign array_update_71362[3] = add_71303 == 32'h0000_0003 ? array_update_71360 : array_update_71352[3];
  assign array_update_71362[4] = add_71303 == 32'h0000_0004 ? array_update_71360 : array_update_71352[4];
  assign array_update_71362[5] = add_71303 == 32'h0000_0005 ? array_update_71360 : array_update_71352[5];
  assign array_update_71362[6] = add_71303 == 32'h0000_0006 ? array_update_71360 : array_update_71352[6];
  assign array_update_71362[7] = add_71303 == 32'h0000_0007 ? array_update_71360 : array_update_71352[7];
  assign array_update_71362[8] = add_71303 == 32'h0000_0008 ? array_update_71360 : array_update_71352[8];
  assign array_update_71362[9] = add_71303 == 32'h0000_0009 ? array_update_71360 : array_update_71352[9];
  assign array_update_71364[0] = add_71305 == 32'h0000_0000 ? array_update_71361 : array_update_71354[0];
  assign array_update_71364[1] = add_71305 == 32'h0000_0001 ? array_update_71361 : array_update_71354[1];
  assign array_update_71364[2] = add_71305 == 32'h0000_0002 ? array_update_71361 : array_update_71354[2];
  assign array_update_71364[3] = add_71305 == 32'h0000_0003 ? array_update_71361 : array_update_71354[3];
  assign array_update_71364[4] = add_71305 == 32'h0000_0004 ? array_update_71361 : array_update_71354[4];
  assign array_update_71364[5] = add_71305 == 32'h0000_0005 ? array_update_71361 : array_update_71354[5];
  assign array_update_71364[6] = add_71305 == 32'h0000_0006 ? array_update_71361 : array_update_71354[6];
  assign array_update_71364[7] = add_71305 == 32'h0000_0007 ? array_update_71361 : array_update_71354[7];
  assign array_update_71364[8] = add_71305 == 32'h0000_0008 ? array_update_71361 : array_update_71354[8];
  assign array_update_71364[9] = add_71305 == 32'h0000_0009 ? array_update_71361 : array_update_71354[9];
  assign array_index_71366 = array_update_71362[add_71303 > 32'h0000_0009 ? 4'h9 : add_71303[3:0]];
  assign add_71367 = add_71357 + 32'h0000_0001;
  assign array_index_71368 = array_update_71364[add_71305 > 32'h0000_0009 ? 4'h9 : add_71305[3:0]];
  assign add_71369 = add_71359 + 32'h0000_0001;
  assign array_update_71370[0] = add_71367 == 32'h0000_0000 ? TestBlock__A_op36 : array_index_71366[0];
  assign array_update_71370[1] = add_71367 == 32'h0000_0001 ? TestBlock__A_op36 : array_index_71366[1];
  assign array_update_71370[2] = add_71367 == 32'h0000_0002 ? TestBlock__A_op36 : array_index_71366[2];
  assign array_update_71370[3] = add_71367 == 32'h0000_0003 ? TestBlock__A_op36 : array_index_71366[3];
  assign array_update_71370[4] = add_71367 == 32'h0000_0004 ? TestBlock__A_op36 : array_index_71366[4];
  assign array_update_71370[5] = add_71367 == 32'h0000_0005 ? TestBlock__A_op36 : array_index_71366[5];
  assign array_update_71370[6] = add_71367 == 32'h0000_0006 ? TestBlock__A_op36 : array_index_71366[6];
  assign array_update_71370[7] = add_71367 == 32'h0000_0007 ? TestBlock__A_op36 : array_index_71366[7];
  assign array_update_71370[8] = add_71367 == 32'h0000_0008 ? TestBlock__A_op36 : array_index_71366[8];
  assign array_update_71370[9] = add_71367 == 32'h0000_0009 ? TestBlock__A_op36 : array_index_71366[9];
  assign array_update_71371[0] = add_71369 == 32'h0000_0000 ? TestBlock__B_op36 : array_index_71368[0];
  assign array_update_71371[1] = add_71369 == 32'h0000_0001 ? TestBlock__B_op36 : array_index_71368[1];
  assign array_update_71371[2] = add_71369 == 32'h0000_0002 ? TestBlock__B_op36 : array_index_71368[2];
  assign array_update_71371[3] = add_71369 == 32'h0000_0003 ? TestBlock__B_op36 : array_index_71368[3];
  assign array_update_71371[4] = add_71369 == 32'h0000_0004 ? TestBlock__B_op36 : array_index_71368[4];
  assign array_update_71371[5] = add_71369 == 32'h0000_0005 ? TestBlock__B_op36 : array_index_71368[5];
  assign array_update_71371[6] = add_71369 == 32'h0000_0006 ? TestBlock__B_op36 : array_index_71368[6];
  assign array_update_71371[7] = add_71369 == 32'h0000_0007 ? TestBlock__B_op36 : array_index_71368[7];
  assign array_update_71371[8] = add_71369 == 32'h0000_0008 ? TestBlock__B_op36 : array_index_71368[8];
  assign array_update_71371[9] = add_71369 == 32'h0000_0009 ? TestBlock__B_op36 : array_index_71368[9];
  assign array_update_71372[0] = add_71303 == 32'h0000_0000 ? array_update_71370 : array_update_71362[0];
  assign array_update_71372[1] = add_71303 == 32'h0000_0001 ? array_update_71370 : array_update_71362[1];
  assign array_update_71372[2] = add_71303 == 32'h0000_0002 ? array_update_71370 : array_update_71362[2];
  assign array_update_71372[3] = add_71303 == 32'h0000_0003 ? array_update_71370 : array_update_71362[3];
  assign array_update_71372[4] = add_71303 == 32'h0000_0004 ? array_update_71370 : array_update_71362[4];
  assign array_update_71372[5] = add_71303 == 32'h0000_0005 ? array_update_71370 : array_update_71362[5];
  assign array_update_71372[6] = add_71303 == 32'h0000_0006 ? array_update_71370 : array_update_71362[6];
  assign array_update_71372[7] = add_71303 == 32'h0000_0007 ? array_update_71370 : array_update_71362[7];
  assign array_update_71372[8] = add_71303 == 32'h0000_0008 ? array_update_71370 : array_update_71362[8];
  assign array_update_71372[9] = add_71303 == 32'h0000_0009 ? array_update_71370 : array_update_71362[9];
  assign array_update_71374[0] = add_71305 == 32'h0000_0000 ? array_update_71371 : array_update_71364[0];
  assign array_update_71374[1] = add_71305 == 32'h0000_0001 ? array_update_71371 : array_update_71364[1];
  assign array_update_71374[2] = add_71305 == 32'h0000_0002 ? array_update_71371 : array_update_71364[2];
  assign array_update_71374[3] = add_71305 == 32'h0000_0003 ? array_update_71371 : array_update_71364[3];
  assign array_update_71374[4] = add_71305 == 32'h0000_0004 ? array_update_71371 : array_update_71364[4];
  assign array_update_71374[5] = add_71305 == 32'h0000_0005 ? array_update_71371 : array_update_71364[5];
  assign array_update_71374[6] = add_71305 == 32'h0000_0006 ? array_update_71371 : array_update_71364[6];
  assign array_update_71374[7] = add_71305 == 32'h0000_0007 ? array_update_71371 : array_update_71364[7];
  assign array_update_71374[8] = add_71305 == 32'h0000_0008 ? array_update_71371 : array_update_71364[8];
  assign array_update_71374[9] = add_71305 == 32'h0000_0009 ? array_update_71371 : array_update_71364[9];
  assign array_index_71376 = array_update_71372[add_71303 > 32'h0000_0009 ? 4'h9 : add_71303[3:0]];
  assign add_71377 = add_71367 + 32'h0000_0001;
  assign array_index_71378 = array_update_71374[add_71305 > 32'h0000_0009 ? 4'h9 : add_71305[3:0]];
  assign add_71379 = add_71369 + 32'h0000_0001;
  assign array_update_71380[0] = add_71377 == 32'h0000_0000 ? TestBlock__A_op37 : array_index_71376[0];
  assign array_update_71380[1] = add_71377 == 32'h0000_0001 ? TestBlock__A_op37 : array_index_71376[1];
  assign array_update_71380[2] = add_71377 == 32'h0000_0002 ? TestBlock__A_op37 : array_index_71376[2];
  assign array_update_71380[3] = add_71377 == 32'h0000_0003 ? TestBlock__A_op37 : array_index_71376[3];
  assign array_update_71380[4] = add_71377 == 32'h0000_0004 ? TestBlock__A_op37 : array_index_71376[4];
  assign array_update_71380[5] = add_71377 == 32'h0000_0005 ? TestBlock__A_op37 : array_index_71376[5];
  assign array_update_71380[6] = add_71377 == 32'h0000_0006 ? TestBlock__A_op37 : array_index_71376[6];
  assign array_update_71380[7] = add_71377 == 32'h0000_0007 ? TestBlock__A_op37 : array_index_71376[7];
  assign array_update_71380[8] = add_71377 == 32'h0000_0008 ? TestBlock__A_op37 : array_index_71376[8];
  assign array_update_71380[9] = add_71377 == 32'h0000_0009 ? TestBlock__A_op37 : array_index_71376[9];
  assign array_update_71381[0] = add_71379 == 32'h0000_0000 ? TestBlock__B_op37 : array_index_71378[0];
  assign array_update_71381[1] = add_71379 == 32'h0000_0001 ? TestBlock__B_op37 : array_index_71378[1];
  assign array_update_71381[2] = add_71379 == 32'h0000_0002 ? TestBlock__B_op37 : array_index_71378[2];
  assign array_update_71381[3] = add_71379 == 32'h0000_0003 ? TestBlock__B_op37 : array_index_71378[3];
  assign array_update_71381[4] = add_71379 == 32'h0000_0004 ? TestBlock__B_op37 : array_index_71378[4];
  assign array_update_71381[5] = add_71379 == 32'h0000_0005 ? TestBlock__B_op37 : array_index_71378[5];
  assign array_update_71381[6] = add_71379 == 32'h0000_0006 ? TestBlock__B_op37 : array_index_71378[6];
  assign array_update_71381[7] = add_71379 == 32'h0000_0007 ? TestBlock__B_op37 : array_index_71378[7];
  assign array_update_71381[8] = add_71379 == 32'h0000_0008 ? TestBlock__B_op37 : array_index_71378[8];
  assign array_update_71381[9] = add_71379 == 32'h0000_0009 ? TestBlock__B_op37 : array_index_71378[9];
  assign array_update_71382[0] = add_71303 == 32'h0000_0000 ? array_update_71380 : array_update_71372[0];
  assign array_update_71382[1] = add_71303 == 32'h0000_0001 ? array_update_71380 : array_update_71372[1];
  assign array_update_71382[2] = add_71303 == 32'h0000_0002 ? array_update_71380 : array_update_71372[2];
  assign array_update_71382[3] = add_71303 == 32'h0000_0003 ? array_update_71380 : array_update_71372[3];
  assign array_update_71382[4] = add_71303 == 32'h0000_0004 ? array_update_71380 : array_update_71372[4];
  assign array_update_71382[5] = add_71303 == 32'h0000_0005 ? array_update_71380 : array_update_71372[5];
  assign array_update_71382[6] = add_71303 == 32'h0000_0006 ? array_update_71380 : array_update_71372[6];
  assign array_update_71382[7] = add_71303 == 32'h0000_0007 ? array_update_71380 : array_update_71372[7];
  assign array_update_71382[8] = add_71303 == 32'h0000_0008 ? array_update_71380 : array_update_71372[8];
  assign array_update_71382[9] = add_71303 == 32'h0000_0009 ? array_update_71380 : array_update_71372[9];
  assign array_update_71384[0] = add_71305 == 32'h0000_0000 ? array_update_71381 : array_update_71374[0];
  assign array_update_71384[1] = add_71305 == 32'h0000_0001 ? array_update_71381 : array_update_71374[1];
  assign array_update_71384[2] = add_71305 == 32'h0000_0002 ? array_update_71381 : array_update_71374[2];
  assign array_update_71384[3] = add_71305 == 32'h0000_0003 ? array_update_71381 : array_update_71374[3];
  assign array_update_71384[4] = add_71305 == 32'h0000_0004 ? array_update_71381 : array_update_71374[4];
  assign array_update_71384[5] = add_71305 == 32'h0000_0005 ? array_update_71381 : array_update_71374[5];
  assign array_update_71384[6] = add_71305 == 32'h0000_0006 ? array_update_71381 : array_update_71374[6];
  assign array_update_71384[7] = add_71305 == 32'h0000_0007 ? array_update_71381 : array_update_71374[7];
  assign array_update_71384[8] = add_71305 == 32'h0000_0008 ? array_update_71381 : array_update_71374[8];
  assign array_update_71384[9] = add_71305 == 32'h0000_0009 ? array_update_71381 : array_update_71374[9];
  assign array_index_71386 = array_update_71382[add_71303 > 32'h0000_0009 ? 4'h9 : add_71303[3:0]];
  assign add_71387 = add_71377 + 32'h0000_0001;
  assign array_index_71388 = array_update_71384[add_71305 > 32'h0000_0009 ? 4'h9 : add_71305[3:0]];
  assign add_71389 = add_71379 + 32'h0000_0001;
  assign array_update_71390[0] = add_71387 == 32'h0000_0000 ? TestBlock__A_op38 : array_index_71386[0];
  assign array_update_71390[1] = add_71387 == 32'h0000_0001 ? TestBlock__A_op38 : array_index_71386[1];
  assign array_update_71390[2] = add_71387 == 32'h0000_0002 ? TestBlock__A_op38 : array_index_71386[2];
  assign array_update_71390[3] = add_71387 == 32'h0000_0003 ? TestBlock__A_op38 : array_index_71386[3];
  assign array_update_71390[4] = add_71387 == 32'h0000_0004 ? TestBlock__A_op38 : array_index_71386[4];
  assign array_update_71390[5] = add_71387 == 32'h0000_0005 ? TestBlock__A_op38 : array_index_71386[5];
  assign array_update_71390[6] = add_71387 == 32'h0000_0006 ? TestBlock__A_op38 : array_index_71386[6];
  assign array_update_71390[7] = add_71387 == 32'h0000_0007 ? TestBlock__A_op38 : array_index_71386[7];
  assign array_update_71390[8] = add_71387 == 32'h0000_0008 ? TestBlock__A_op38 : array_index_71386[8];
  assign array_update_71390[9] = add_71387 == 32'h0000_0009 ? TestBlock__A_op38 : array_index_71386[9];
  assign array_update_71391[0] = add_71389 == 32'h0000_0000 ? TestBlock__B_op38 : array_index_71388[0];
  assign array_update_71391[1] = add_71389 == 32'h0000_0001 ? TestBlock__B_op38 : array_index_71388[1];
  assign array_update_71391[2] = add_71389 == 32'h0000_0002 ? TestBlock__B_op38 : array_index_71388[2];
  assign array_update_71391[3] = add_71389 == 32'h0000_0003 ? TestBlock__B_op38 : array_index_71388[3];
  assign array_update_71391[4] = add_71389 == 32'h0000_0004 ? TestBlock__B_op38 : array_index_71388[4];
  assign array_update_71391[5] = add_71389 == 32'h0000_0005 ? TestBlock__B_op38 : array_index_71388[5];
  assign array_update_71391[6] = add_71389 == 32'h0000_0006 ? TestBlock__B_op38 : array_index_71388[6];
  assign array_update_71391[7] = add_71389 == 32'h0000_0007 ? TestBlock__B_op38 : array_index_71388[7];
  assign array_update_71391[8] = add_71389 == 32'h0000_0008 ? TestBlock__B_op38 : array_index_71388[8];
  assign array_update_71391[9] = add_71389 == 32'h0000_0009 ? TestBlock__B_op38 : array_index_71388[9];
  assign array_update_71392[0] = add_71303 == 32'h0000_0000 ? array_update_71390 : array_update_71382[0];
  assign array_update_71392[1] = add_71303 == 32'h0000_0001 ? array_update_71390 : array_update_71382[1];
  assign array_update_71392[2] = add_71303 == 32'h0000_0002 ? array_update_71390 : array_update_71382[2];
  assign array_update_71392[3] = add_71303 == 32'h0000_0003 ? array_update_71390 : array_update_71382[3];
  assign array_update_71392[4] = add_71303 == 32'h0000_0004 ? array_update_71390 : array_update_71382[4];
  assign array_update_71392[5] = add_71303 == 32'h0000_0005 ? array_update_71390 : array_update_71382[5];
  assign array_update_71392[6] = add_71303 == 32'h0000_0006 ? array_update_71390 : array_update_71382[6];
  assign array_update_71392[7] = add_71303 == 32'h0000_0007 ? array_update_71390 : array_update_71382[7];
  assign array_update_71392[8] = add_71303 == 32'h0000_0008 ? array_update_71390 : array_update_71382[8];
  assign array_update_71392[9] = add_71303 == 32'h0000_0009 ? array_update_71390 : array_update_71382[9];
  assign array_update_71394[0] = add_71305 == 32'h0000_0000 ? array_update_71391 : array_update_71384[0];
  assign array_update_71394[1] = add_71305 == 32'h0000_0001 ? array_update_71391 : array_update_71384[1];
  assign array_update_71394[2] = add_71305 == 32'h0000_0002 ? array_update_71391 : array_update_71384[2];
  assign array_update_71394[3] = add_71305 == 32'h0000_0003 ? array_update_71391 : array_update_71384[3];
  assign array_update_71394[4] = add_71305 == 32'h0000_0004 ? array_update_71391 : array_update_71384[4];
  assign array_update_71394[5] = add_71305 == 32'h0000_0005 ? array_update_71391 : array_update_71384[5];
  assign array_update_71394[6] = add_71305 == 32'h0000_0006 ? array_update_71391 : array_update_71384[6];
  assign array_update_71394[7] = add_71305 == 32'h0000_0007 ? array_update_71391 : array_update_71384[7];
  assign array_update_71394[8] = add_71305 == 32'h0000_0008 ? array_update_71391 : array_update_71384[8];
  assign array_update_71394[9] = add_71305 == 32'h0000_0009 ? array_update_71391 : array_update_71384[9];
  assign array_index_71396 = array_update_71392[add_71303 > 32'h0000_0009 ? 4'h9 : add_71303[3:0]];
  assign add_71397 = add_71387 + 32'h0000_0001;
  assign array_index_71398 = array_update_71394[add_71305 > 32'h0000_0009 ? 4'h9 : add_71305[3:0]];
  assign add_71399 = add_71389 + 32'h0000_0001;
  assign array_update_71400[0] = add_71397 == 32'h0000_0000 ? TestBlock__A_op39 : array_index_71396[0];
  assign array_update_71400[1] = add_71397 == 32'h0000_0001 ? TestBlock__A_op39 : array_index_71396[1];
  assign array_update_71400[2] = add_71397 == 32'h0000_0002 ? TestBlock__A_op39 : array_index_71396[2];
  assign array_update_71400[3] = add_71397 == 32'h0000_0003 ? TestBlock__A_op39 : array_index_71396[3];
  assign array_update_71400[4] = add_71397 == 32'h0000_0004 ? TestBlock__A_op39 : array_index_71396[4];
  assign array_update_71400[5] = add_71397 == 32'h0000_0005 ? TestBlock__A_op39 : array_index_71396[5];
  assign array_update_71400[6] = add_71397 == 32'h0000_0006 ? TestBlock__A_op39 : array_index_71396[6];
  assign array_update_71400[7] = add_71397 == 32'h0000_0007 ? TestBlock__A_op39 : array_index_71396[7];
  assign array_update_71400[8] = add_71397 == 32'h0000_0008 ? TestBlock__A_op39 : array_index_71396[8];
  assign array_update_71400[9] = add_71397 == 32'h0000_0009 ? TestBlock__A_op39 : array_index_71396[9];
  assign array_update_71402[0] = add_71399 == 32'h0000_0000 ? TestBlock__B_op39 : array_index_71398[0];
  assign array_update_71402[1] = add_71399 == 32'h0000_0001 ? TestBlock__B_op39 : array_index_71398[1];
  assign array_update_71402[2] = add_71399 == 32'h0000_0002 ? TestBlock__B_op39 : array_index_71398[2];
  assign array_update_71402[3] = add_71399 == 32'h0000_0003 ? TestBlock__B_op39 : array_index_71398[3];
  assign array_update_71402[4] = add_71399 == 32'h0000_0004 ? TestBlock__B_op39 : array_index_71398[4];
  assign array_update_71402[5] = add_71399 == 32'h0000_0005 ? TestBlock__B_op39 : array_index_71398[5];
  assign array_update_71402[6] = add_71399 == 32'h0000_0006 ? TestBlock__B_op39 : array_index_71398[6];
  assign array_update_71402[7] = add_71399 == 32'h0000_0007 ? TestBlock__B_op39 : array_index_71398[7];
  assign array_update_71402[8] = add_71399 == 32'h0000_0008 ? TestBlock__B_op39 : array_index_71398[8];
  assign array_update_71402[9] = add_71399 == 32'h0000_0009 ? TestBlock__B_op39 : array_index_71398[9];
  assign array_update_71404[0] = add_71303 == 32'h0000_0000 ? array_update_71400 : array_update_71392[0];
  assign array_update_71404[1] = add_71303 == 32'h0000_0001 ? array_update_71400 : array_update_71392[1];
  assign array_update_71404[2] = add_71303 == 32'h0000_0002 ? array_update_71400 : array_update_71392[2];
  assign array_update_71404[3] = add_71303 == 32'h0000_0003 ? array_update_71400 : array_update_71392[3];
  assign array_update_71404[4] = add_71303 == 32'h0000_0004 ? array_update_71400 : array_update_71392[4];
  assign array_update_71404[5] = add_71303 == 32'h0000_0005 ? array_update_71400 : array_update_71392[5];
  assign array_update_71404[6] = add_71303 == 32'h0000_0006 ? array_update_71400 : array_update_71392[6];
  assign array_update_71404[7] = add_71303 == 32'h0000_0007 ? array_update_71400 : array_update_71392[7];
  assign array_update_71404[8] = add_71303 == 32'h0000_0008 ? array_update_71400 : array_update_71392[8];
  assign array_update_71404[9] = add_71303 == 32'h0000_0009 ? array_update_71400 : array_update_71392[9];
  assign add_71405 = add_71303 + 32'h0000_0001;
  assign array_update_71406[0] = add_71305 == 32'h0000_0000 ? array_update_71402 : array_update_71394[0];
  assign array_update_71406[1] = add_71305 == 32'h0000_0001 ? array_update_71402 : array_update_71394[1];
  assign array_update_71406[2] = add_71305 == 32'h0000_0002 ? array_update_71402 : array_update_71394[2];
  assign array_update_71406[3] = add_71305 == 32'h0000_0003 ? array_update_71402 : array_update_71394[3];
  assign array_update_71406[4] = add_71305 == 32'h0000_0004 ? array_update_71402 : array_update_71394[4];
  assign array_update_71406[5] = add_71305 == 32'h0000_0005 ? array_update_71402 : array_update_71394[5];
  assign array_update_71406[6] = add_71305 == 32'h0000_0006 ? array_update_71402 : array_update_71394[6];
  assign array_update_71406[7] = add_71305 == 32'h0000_0007 ? array_update_71402 : array_update_71394[7];
  assign array_update_71406[8] = add_71305 == 32'h0000_0008 ? array_update_71402 : array_update_71394[8];
  assign array_update_71406[9] = add_71305 == 32'h0000_0009 ? array_update_71402 : array_update_71394[9];
  assign add_71407 = add_71305 + 32'h0000_0001;
  assign array_index_71408 = array_update_71404[add_71405 > 32'h0000_0009 ? 4'h9 : add_71405[3:0]];
  assign literal_71409 = 32'h0000_0000;
  assign array_index_71410 = array_update_71406[add_71407 > 32'h0000_0009 ? 4'h9 : add_71407[3:0]];
  assign literal_71411 = 32'h0000_0000;
  assign array_update_71412[0] = literal_71409 == 32'h0000_0000 ? TestBlock__A_op40 : array_index_71408[0];
  assign array_update_71412[1] = literal_71409 == 32'h0000_0001 ? TestBlock__A_op40 : array_index_71408[1];
  assign array_update_71412[2] = literal_71409 == 32'h0000_0002 ? TestBlock__A_op40 : array_index_71408[2];
  assign array_update_71412[3] = literal_71409 == 32'h0000_0003 ? TestBlock__A_op40 : array_index_71408[3];
  assign array_update_71412[4] = literal_71409 == 32'h0000_0004 ? TestBlock__A_op40 : array_index_71408[4];
  assign array_update_71412[5] = literal_71409 == 32'h0000_0005 ? TestBlock__A_op40 : array_index_71408[5];
  assign array_update_71412[6] = literal_71409 == 32'h0000_0006 ? TestBlock__A_op40 : array_index_71408[6];
  assign array_update_71412[7] = literal_71409 == 32'h0000_0007 ? TestBlock__A_op40 : array_index_71408[7];
  assign array_update_71412[8] = literal_71409 == 32'h0000_0008 ? TestBlock__A_op40 : array_index_71408[8];
  assign array_update_71412[9] = literal_71409 == 32'h0000_0009 ? TestBlock__A_op40 : array_index_71408[9];
  assign array_update_71413[0] = literal_71411 == 32'h0000_0000 ? TestBlock__B_op40 : array_index_71410[0];
  assign array_update_71413[1] = literal_71411 == 32'h0000_0001 ? TestBlock__B_op40 : array_index_71410[1];
  assign array_update_71413[2] = literal_71411 == 32'h0000_0002 ? TestBlock__B_op40 : array_index_71410[2];
  assign array_update_71413[3] = literal_71411 == 32'h0000_0003 ? TestBlock__B_op40 : array_index_71410[3];
  assign array_update_71413[4] = literal_71411 == 32'h0000_0004 ? TestBlock__B_op40 : array_index_71410[4];
  assign array_update_71413[5] = literal_71411 == 32'h0000_0005 ? TestBlock__B_op40 : array_index_71410[5];
  assign array_update_71413[6] = literal_71411 == 32'h0000_0006 ? TestBlock__B_op40 : array_index_71410[6];
  assign array_update_71413[7] = literal_71411 == 32'h0000_0007 ? TestBlock__B_op40 : array_index_71410[7];
  assign array_update_71413[8] = literal_71411 == 32'h0000_0008 ? TestBlock__B_op40 : array_index_71410[8];
  assign array_update_71413[9] = literal_71411 == 32'h0000_0009 ? TestBlock__B_op40 : array_index_71410[9];
  assign array_update_71414[0] = add_71405 == 32'h0000_0000 ? array_update_71412 : array_update_71404[0];
  assign array_update_71414[1] = add_71405 == 32'h0000_0001 ? array_update_71412 : array_update_71404[1];
  assign array_update_71414[2] = add_71405 == 32'h0000_0002 ? array_update_71412 : array_update_71404[2];
  assign array_update_71414[3] = add_71405 == 32'h0000_0003 ? array_update_71412 : array_update_71404[3];
  assign array_update_71414[4] = add_71405 == 32'h0000_0004 ? array_update_71412 : array_update_71404[4];
  assign array_update_71414[5] = add_71405 == 32'h0000_0005 ? array_update_71412 : array_update_71404[5];
  assign array_update_71414[6] = add_71405 == 32'h0000_0006 ? array_update_71412 : array_update_71404[6];
  assign array_update_71414[7] = add_71405 == 32'h0000_0007 ? array_update_71412 : array_update_71404[7];
  assign array_update_71414[8] = add_71405 == 32'h0000_0008 ? array_update_71412 : array_update_71404[8];
  assign array_update_71414[9] = add_71405 == 32'h0000_0009 ? array_update_71412 : array_update_71404[9];
  assign array_update_71416[0] = add_71407 == 32'h0000_0000 ? array_update_71413 : array_update_71406[0];
  assign array_update_71416[1] = add_71407 == 32'h0000_0001 ? array_update_71413 : array_update_71406[1];
  assign array_update_71416[2] = add_71407 == 32'h0000_0002 ? array_update_71413 : array_update_71406[2];
  assign array_update_71416[3] = add_71407 == 32'h0000_0003 ? array_update_71413 : array_update_71406[3];
  assign array_update_71416[4] = add_71407 == 32'h0000_0004 ? array_update_71413 : array_update_71406[4];
  assign array_update_71416[5] = add_71407 == 32'h0000_0005 ? array_update_71413 : array_update_71406[5];
  assign array_update_71416[6] = add_71407 == 32'h0000_0006 ? array_update_71413 : array_update_71406[6];
  assign array_update_71416[7] = add_71407 == 32'h0000_0007 ? array_update_71413 : array_update_71406[7];
  assign array_update_71416[8] = add_71407 == 32'h0000_0008 ? array_update_71413 : array_update_71406[8];
  assign array_update_71416[9] = add_71407 == 32'h0000_0009 ? array_update_71413 : array_update_71406[9];
  assign array_index_71418 = array_update_71414[add_71405 > 32'h0000_0009 ? 4'h9 : add_71405[3:0]];
  assign add_71419 = literal_71409 + 32'h0000_0001;
  assign array_index_71420 = array_update_71416[add_71407 > 32'h0000_0009 ? 4'h9 : add_71407[3:0]];
  assign add_71421 = literal_71411 + 32'h0000_0001;
  assign array_update_71422[0] = add_71419 == 32'h0000_0000 ? TestBlock__A_op41 : array_index_71418[0];
  assign array_update_71422[1] = add_71419 == 32'h0000_0001 ? TestBlock__A_op41 : array_index_71418[1];
  assign array_update_71422[2] = add_71419 == 32'h0000_0002 ? TestBlock__A_op41 : array_index_71418[2];
  assign array_update_71422[3] = add_71419 == 32'h0000_0003 ? TestBlock__A_op41 : array_index_71418[3];
  assign array_update_71422[4] = add_71419 == 32'h0000_0004 ? TestBlock__A_op41 : array_index_71418[4];
  assign array_update_71422[5] = add_71419 == 32'h0000_0005 ? TestBlock__A_op41 : array_index_71418[5];
  assign array_update_71422[6] = add_71419 == 32'h0000_0006 ? TestBlock__A_op41 : array_index_71418[6];
  assign array_update_71422[7] = add_71419 == 32'h0000_0007 ? TestBlock__A_op41 : array_index_71418[7];
  assign array_update_71422[8] = add_71419 == 32'h0000_0008 ? TestBlock__A_op41 : array_index_71418[8];
  assign array_update_71422[9] = add_71419 == 32'h0000_0009 ? TestBlock__A_op41 : array_index_71418[9];
  assign array_update_71423[0] = add_71421 == 32'h0000_0000 ? TestBlock__B_op41 : array_index_71420[0];
  assign array_update_71423[1] = add_71421 == 32'h0000_0001 ? TestBlock__B_op41 : array_index_71420[1];
  assign array_update_71423[2] = add_71421 == 32'h0000_0002 ? TestBlock__B_op41 : array_index_71420[2];
  assign array_update_71423[3] = add_71421 == 32'h0000_0003 ? TestBlock__B_op41 : array_index_71420[3];
  assign array_update_71423[4] = add_71421 == 32'h0000_0004 ? TestBlock__B_op41 : array_index_71420[4];
  assign array_update_71423[5] = add_71421 == 32'h0000_0005 ? TestBlock__B_op41 : array_index_71420[5];
  assign array_update_71423[6] = add_71421 == 32'h0000_0006 ? TestBlock__B_op41 : array_index_71420[6];
  assign array_update_71423[7] = add_71421 == 32'h0000_0007 ? TestBlock__B_op41 : array_index_71420[7];
  assign array_update_71423[8] = add_71421 == 32'h0000_0008 ? TestBlock__B_op41 : array_index_71420[8];
  assign array_update_71423[9] = add_71421 == 32'h0000_0009 ? TestBlock__B_op41 : array_index_71420[9];
  assign array_update_71424[0] = add_71405 == 32'h0000_0000 ? array_update_71422 : array_update_71414[0];
  assign array_update_71424[1] = add_71405 == 32'h0000_0001 ? array_update_71422 : array_update_71414[1];
  assign array_update_71424[2] = add_71405 == 32'h0000_0002 ? array_update_71422 : array_update_71414[2];
  assign array_update_71424[3] = add_71405 == 32'h0000_0003 ? array_update_71422 : array_update_71414[3];
  assign array_update_71424[4] = add_71405 == 32'h0000_0004 ? array_update_71422 : array_update_71414[4];
  assign array_update_71424[5] = add_71405 == 32'h0000_0005 ? array_update_71422 : array_update_71414[5];
  assign array_update_71424[6] = add_71405 == 32'h0000_0006 ? array_update_71422 : array_update_71414[6];
  assign array_update_71424[7] = add_71405 == 32'h0000_0007 ? array_update_71422 : array_update_71414[7];
  assign array_update_71424[8] = add_71405 == 32'h0000_0008 ? array_update_71422 : array_update_71414[8];
  assign array_update_71424[9] = add_71405 == 32'h0000_0009 ? array_update_71422 : array_update_71414[9];
  assign array_update_71426[0] = add_71407 == 32'h0000_0000 ? array_update_71423 : array_update_71416[0];
  assign array_update_71426[1] = add_71407 == 32'h0000_0001 ? array_update_71423 : array_update_71416[1];
  assign array_update_71426[2] = add_71407 == 32'h0000_0002 ? array_update_71423 : array_update_71416[2];
  assign array_update_71426[3] = add_71407 == 32'h0000_0003 ? array_update_71423 : array_update_71416[3];
  assign array_update_71426[4] = add_71407 == 32'h0000_0004 ? array_update_71423 : array_update_71416[4];
  assign array_update_71426[5] = add_71407 == 32'h0000_0005 ? array_update_71423 : array_update_71416[5];
  assign array_update_71426[6] = add_71407 == 32'h0000_0006 ? array_update_71423 : array_update_71416[6];
  assign array_update_71426[7] = add_71407 == 32'h0000_0007 ? array_update_71423 : array_update_71416[7];
  assign array_update_71426[8] = add_71407 == 32'h0000_0008 ? array_update_71423 : array_update_71416[8];
  assign array_update_71426[9] = add_71407 == 32'h0000_0009 ? array_update_71423 : array_update_71416[9];
  assign array_index_71428 = array_update_71424[add_71405 > 32'h0000_0009 ? 4'h9 : add_71405[3:0]];
  assign add_71429 = add_71419 + 32'h0000_0001;
  assign array_index_71430 = array_update_71426[add_71407 > 32'h0000_0009 ? 4'h9 : add_71407[3:0]];
  assign add_71431 = add_71421 + 32'h0000_0001;
  assign array_update_71432[0] = add_71429 == 32'h0000_0000 ? TestBlock__A_op42 : array_index_71428[0];
  assign array_update_71432[1] = add_71429 == 32'h0000_0001 ? TestBlock__A_op42 : array_index_71428[1];
  assign array_update_71432[2] = add_71429 == 32'h0000_0002 ? TestBlock__A_op42 : array_index_71428[2];
  assign array_update_71432[3] = add_71429 == 32'h0000_0003 ? TestBlock__A_op42 : array_index_71428[3];
  assign array_update_71432[4] = add_71429 == 32'h0000_0004 ? TestBlock__A_op42 : array_index_71428[4];
  assign array_update_71432[5] = add_71429 == 32'h0000_0005 ? TestBlock__A_op42 : array_index_71428[5];
  assign array_update_71432[6] = add_71429 == 32'h0000_0006 ? TestBlock__A_op42 : array_index_71428[6];
  assign array_update_71432[7] = add_71429 == 32'h0000_0007 ? TestBlock__A_op42 : array_index_71428[7];
  assign array_update_71432[8] = add_71429 == 32'h0000_0008 ? TestBlock__A_op42 : array_index_71428[8];
  assign array_update_71432[9] = add_71429 == 32'h0000_0009 ? TestBlock__A_op42 : array_index_71428[9];
  assign array_update_71433[0] = add_71431 == 32'h0000_0000 ? TestBlock__B_op42 : array_index_71430[0];
  assign array_update_71433[1] = add_71431 == 32'h0000_0001 ? TestBlock__B_op42 : array_index_71430[1];
  assign array_update_71433[2] = add_71431 == 32'h0000_0002 ? TestBlock__B_op42 : array_index_71430[2];
  assign array_update_71433[3] = add_71431 == 32'h0000_0003 ? TestBlock__B_op42 : array_index_71430[3];
  assign array_update_71433[4] = add_71431 == 32'h0000_0004 ? TestBlock__B_op42 : array_index_71430[4];
  assign array_update_71433[5] = add_71431 == 32'h0000_0005 ? TestBlock__B_op42 : array_index_71430[5];
  assign array_update_71433[6] = add_71431 == 32'h0000_0006 ? TestBlock__B_op42 : array_index_71430[6];
  assign array_update_71433[7] = add_71431 == 32'h0000_0007 ? TestBlock__B_op42 : array_index_71430[7];
  assign array_update_71433[8] = add_71431 == 32'h0000_0008 ? TestBlock__B_op42 : array_index_71430[8];
  assign array_update_71433[9] = add_71431 == 32'h0000_0009 ? TestBlock__B_op42 : array_index_71430[9];
  assign array_update_71434[0] = add_71405 == 32'h0000_0000 ? array_update_71432 : array_update_71424[0];
  assign array_update_71434[1] = add_71405 == 32'h0000_0001 ? array_update_71432 : array_update_71424[1];
  assign array_update_71434[2] = add_71405 == 32'h0000_0002 ? array_update_71432 : array_update_71424[2];
  assign array_update_71434[3] = add_71405 == 32'h0000_0003 ? array_update_71432 : array_update_71424[3];
  assign array_update_71434[4] = add_71405 == 32'h0000_0004 ? array_update_71432 : array_update_71424[4];
  assign array_update_71434[5] = add_71405 == 32'h0000_0005 ? array_update_71432 : array_update_71424[5];
  assign array_update_71434[6] = add_71405 == 32'h0000_0006 ? array_update_71432 : array_update_71424[6];
  assign array_update_71434[7] = add_71405 == 32'h0000_0007 ? array_update_71432 : array_update_71424[7];
  assign array_update_71434[8] = add_71405 == 32'h0000_0008 ? array_update_71432 : array_update_71424[8];
  assign array_update_71434[9] = add_71405 == 32'h0000_0009 ? array_update_71432 : array_update_71424[9];
  assign array_update_71436[0] = add_71407 == 32'h0000_0000 ? array_update_71433 : array_update_71426[0];
  assign array_update_71436[1] = add_71407 == 32'h0000_0001 ? array_update_71433 : array_update_71426[1];
  assign array_update_71436[2] = add_71407 == 32'h0000_0002 ? array_update_71433 : array_update_71426[2];
  assign array_update_71436[3] = add_71407 == 32'h0000_0003 ? array_update_71433 : array_update_71426[3];
  assign array_update_71436[4] = add_71407 == 32'h0000_0004 ? array_update_71433 : array_update_71426[4];
  assign array_update_71436[5] = add_71407 == 32'h0000_0005 ? array_update_71433 : array_update_71426[5];
  assign array_update_71436[6] = add_71407 == 32'h0000_0006 ? array_update_71433 : array_update_71426[6];
  assign array_update_71436[7] = add_71407 == 32'h0000_0007 ? array_update_71433 : array_update_71426[7];
  assign array_update_71436[8] = add_71407 == 32'h0000_0008 ? array_update_71433 : array_update_71426[8];
  assign array_update_71436[9] = add_71407 == 32'h0000_0009 ? array_update_71433 : array_update_71426[9];
  assign array_index_71438 = array_update_71434[add_71405 > 32'h0000_0009 ? 4'h9 : add_71405[3:0]];
  assign add_71439 = add_71429 + 32'h0000_0001;
  assign array_index_71440 = array_update_71436[add_71407 > 32'h0000_0009 ? 4'h9 : add_71407[3:0]];
  assign add_71441 = add_71431 + 32'h0000_0001;
  assign array_update_71442[0] = add_71439 == 32'h0000_0000 ? TestBlock__A_op43 : array_index_71438[0];
  assign array_update_71442[1] = add_71439 == 32'h0000_0001 ? TestBlock__A_op43 : array_index_71438[1];
  assign array_update_71442[2] = add_71439 == 32'h0000_0002 ? TestBlock__A_op43 : array_index_71438[2];
  assign array_update_71442[3] = add_71439 == 32'h0000_0003 ? TestBlock__A_op43 : array_index_71438[3];
  assign array_update_71442[4] = add_71439 == 32'h0000_0004 ? TestBlock__A_op43 : array_index_71438[4];
  assign array_update_71442[5] = add_71439 == 32'h0000_0005 ? TestBlock__A_op43 : array_index_71438[5];
  assign array_update_71442[6] = add_71439 == 32'h0000_0006 ? TestBlock__A_op43 : array_index_71438[6];
  assign array_update_71442[7] = add_71439 == 32'h0000_0007 ? TestBlock__A_op43 : array_index_71438[7];
  assign array_update_71442[8] = add_71439 == 32'h0000_0008 ? TestBlock__A_op43 : array_index_71438[8];
  assign array_update_71442[9] = add_71439 == 32'h0000_0009 ? TestBlock__A_op43 : array_index_71438[9];
  assign array_update_71443[0] = add_71441 == 32'h0000_0000 ? TestBlock__B_op43 : array_index_71440[0];
  assign array_update_71443[1] = add_71441 == 32'h0000_0001 ? TestBlock__B_op43 : array_index_71440[1];
  assign array_update_71443[2] = add_71441 == 32'h0000_0002 ? TestBlock__B_op43 : array_index_71440[2];
  assign array_update_71443[3] = add_71441 == 32'h0000_0003 ? TestBlock__B_op43 : array_index_71440[3];
  assign array_update_71443[4] = add_71441 == 32'h0000_0004 ? TestBlock__B_op43 : array_index_71440[4];
  assign array_update_71443[5] = add_71441 == 32'h0000_0005 ? TestBlock__B_op43 : array_index_71440[5];
  assign array_update_71443[6] = add_71441 == 32'h0000_0006 ? TestBlock__B_op43 : array_index_71440[6];
  assign array_update_71443[7] = add_71441 == 32'h0000_0007 ? TestBlock__B_op43 : array_index_71440[7];
  assign array_update_71443[8] = add_71441 == 32'h0000_0008 ? TestBlock__B_op43 : array_index_71440[8];
  assign array_update_71443[9] = add_71441 == 32'h0000_0009 ? TestBlock__B_op43 : array_index_71440[9];
  assign array_update_71444[0] = add_71405 == 32'h0000_0000 ? array_update_71442 : array_update_71434[0];
  assign array_update_71444[1] = add_71405 == 32'h0000_0001 ? array_update_71442 : array_update_71434[1];
  assign array_update_71444[2] = add_71405 == 32'h0000_0002 ? array_update_71442 : array_update_71434[2];
  assign array_update_71444[3] = add_71405 == 32'h0000_0003 ? array_update_71442 : array_update_71434[3];
  assign array_update_71444[4] = add_71405 == 32'h0000_0004 ? array_update_71442 : array_update_71434[4];
  assign array_update_71444[5] = add_71405 == 32'h0000_0005 ? array_update_71442 : array_update_71434[5];
  assign array_update_71444[6] = add_71405 == 32'h0000_0006 ? array_update_71442 : array_update_71434[6];
  assign array_update_71444[7] = add_71405 == 32'h0000_0007 ? array_update_71442 : array_update_71434[7];
  assign array_update_71444[8] = add_71405 == 32'h0000_0008 ? array_update_71442 : array_update_71434[8];
  assign array_update_71444[9] = add_71405 == 32'h0000_0009 ? array_update_71442 : array_update_71434[9];
  assign array_update_71446[0] = add_71407 == 32'h0000_0000 ? array_update_71443 : array_update_71436[0];
  assign array_update_71446[1] = add_71407 == 32'h0000_0001 ? array_update_71443 : array_update_71436[1];
  assign array_update_71446[2] = add_71407 == 32'h0000_0002 ? array_update_71443 : array_update_71436[2];
  assign array_update_71446[3] = add_71407 == 32'h0000_0003 ? array_update_71443 : array_update_71436[3];
  assign array_update_71446[4] = add_71407 == 32'h0000_0004 ? array_update_71443 : array_update_71436[4];
  assign array_update_71446[5] = add_71407 == 32'h0000_0005 ? array_update_71443 : array_update_71436[5];
  assign array_update_71446[6] = add_71407 == 32'h0000_0006 ? array_update_71443 : array_update_71436[6];
  assign array_update_71446[7] = add_71407 == 32'h0000_0007 ? array_update_71443 : array_update_71436[7];
  assign array_update_71446[8] = add_71407 == 32'h0000_0008 ? array_update_71443 : array_update_71436[8];
  assign array_update_71446[9] = add_71407 == 32'h0000_0009 ? array_update_71443 : array_update_71436[9];
  assign array_index_71448 = array_update_71444[add_71405 > 32'h0000_0009 ? 4'h9 : add_71405[3:0]];
  assign add_71449 = add_71439 + 32'h0000_0001;
  assign array_index_71450 = array_update_71446[add_71407 > 32'h0000_0009 ? 4'h9 : add_71407[3:0]];
  assign add_71451 = add_71441 + 32'h0000_0001;
  assign array_update_71452[0] = add_71449 == 32'h0000_0000 ? TestBlock__A_op44 : array_index_71448[0];
  assign array_update_71452[1] = add_71449 == 32'h0000_0001 ? TestBlock__A_op44 : array_index_71448[1];
  assign array_update_71452[2] = add_71449 == 32'h0000_0002 ? TestBlock__A_op44 : array_index_71448[2];
  assign array_update_71452[3] = add_71449 == 32'h0000_0003 ? TestBlock__A_op44 : array_index_71448[3];
  assign array_update_71452[4] = add_71449 == 32'h0000_0004 ? TestBlock__A_op44 : array_index_71448[4];
  assign array_update_71452[5] = add_71449 == 32'h0000_0005 ? TestBlock__A_op44 : array_index_71448[5];
  assign array_update_71452[6] = add_71449 == 32'h0000_0006 ? TestBlock__A_op44 : array_index_71448[6];
  assign array_update_71452[7] = add_71449 == 32'h0000_0007 ? TestBlock__A_op44 : array_index_71448[7];
  assign array_update_71452[8] = add_71449 == 32'h0000_0008 ? TestBlock__A_op44 : array_index_71448[8];
  assign array_update_71452[9] = add_71449 == 32'h0000_0009 ? TestBlock__A_op44 : array_index_71448[9];
  assign array_update_71453[0] = add_71451 == 32'h0000_0000 ? TestBlock__B_op44 : array_index_71450[0];
  assign array_update_71453[1] = add_71451 == 32'h0000_0001 ? TestBlock__B_op44 : array_index_71450[1];
  assign array_update_71453[2] = add_71451 == 32'h0000_0002 ? TestBlock__B_op44 : array_index_71450[2];
  assign array_update_71453[3] = add_71451 == 32'h0000_0003 ? TestBlock__B_op44 : array_index_71450[3];
  assign array_update_71453[4] = add_71451 == 32'h0000_0004 ? TestBlock__B_op44 : array_index_71450[4];
  assign array_update_71453[5] = add_71451 == 32'h0000_0005 ? TestBlock__B_op44 : array_index_71450[5];
  assign array_update_71453[6] = add_71451 == 32'h0000_0006 ? TestBlock__B_op44 : array_index_71450[6];
  assign array_update_71453[7] = add_71451 == 32'h0000_0007 ? TestBlock__B_op44 : array_index_71450[7];
  assign array_update_71453[8] = add_71451 == 32'h0000_0008 ? TestBlock__B_op44 : array_index_71450[8];
  assign array_update_71453[9] = add_71451 == 32'h0000_0009 ? TestBlock__B_op44 : array_index_71450[9];
  assign array_update_71454[0] = add_71405 == 32'h0000_0000 ? array_update_71452 : array_update_71444[0];
  assign array_update_71454[1] = add_71405 == 32'h0000_0001 ? array_update_71452 : array_update_71444[1];
  assign array_update_71454[2] = add_71405 == 32'h0000_0002 ? array_update_71452 : array_update_71444[2];
  assign array_update_71454[3] = add_71405 == 32'h0000_0003 ? array_update_71452 : array_update_71444[3];
  assign array_update_71454[4] = add_71405 == 32'h0000_0004 ? array_update_71452 : array_update_71444[4];
  assign array_update_71454[5] = add_71405 == 32'h0000_0005 ? array_update_71452 : array_update_71444[5];
  assign array_update_71454[6] = add_71405 == 32'h0000_0006 ? array_update_71452 : array_update_71444[6];
  assign array_update_71454[7] = add_71405 == 32'h0000_0007 ? array_update_71452 : array_update_71444[7];
  assign array_update_71454[8] = add_71405 == 32'h0000_0008 ? array_update_71452 : array_update_71444[8];
  assign array_update_71454[9] = add_71405 == 32'h0000_0009 ? array_update_71452 : array_update_71444[9];
  assign array_update_71456[0] = add_71407 == 32'h0000_0000 ? array_update_71453 : array_update_71446[0];
  assign array_update_71456[1] = add_71407 == 32'h0000_0001 ? array_update_71453 : array_update_71446[1];
  assign array_update_71456[2] = add_71407 == 32'h0000_0002 ? array_update_71453 : array_update_71446[2];
  assign array_update_71456[3] = add_71407 == 32'h0000_0003 ? array_update_71453 : array_update_71446[3];
  assign array_update_71456[4] = add_71407 == 32'h0000_0004 ? array_update_71453 : array_update_71446[4];
  assign array_update_71456[5] = add_71407 == 32'h0000_0005 ? array_update_71453 : array_update_71446[5];
  assign array_update_71456[6] = add_71407 == 32'h0000_0006 ? array_update_71453 : array_update_71446[6];
  assign array_update_71456[7] = add_71407 == 32'h0000_0007 ? array_update_71453 : array_update_71446[7];
  assign array_update_71456[8] = add_71407 == 32'h0000_0008 ? array_update_71453 : array_update_71446[8];
  assign array_update_71456[9] = add_71407 == 32'h0000_0009 ? array_update_71453 : array_update_71446[9];
  assign array_index_71458 = array_update_71454[add_71405 > 32'h0000_0009 ? 4'h9 : add_71405[3:0]];
  assign add_71459 = add_71449 + 32'h0000_0001;
  assign array_index_71460 = array_update_71456[add_71407 > 32'h0000_0009 ? 4'h9 : add_71407[3:0]];
  assign add_71461 = add_71451 + 32'h0000_0001;
  assign array_update_71462[0] = add_71459 == 32'h0000_0000 ? TestBlock__A_op45 : array_index_71458[0];
  assign array_update_71462[1] = add_71459 == 32'h0000_0001 ? TestBlock__A_op45 : array_index_71458[1];
  assign array_update_71462[2] = add_71459 == 32'h0000_0002 ? TestBlock__A_op45 : array_index_71458[2];
  assign array_update_71462[3] = add_71459 == 32'h0000_0003 ? TestBlock__A_op45 : array_index_71458[3];
  assign array_update_71462[4] = add_71459 == 32'h0000_0004 ? TestBlock__A_op45 : array_index_71458[4];
  assign array_update_71462[5] = add_71459 == 32'h0000_0005 ? TestBlock__A_op45 : array_index_71458[5];
  assign array_update_71462[6] = add_71459 == 32'h0000_0006 ? TestBlock__A_op45 : array_index_71458[6];
  assign array_update_71462[7] = add_71459 == 32'h0000_0007 ? TestBlock__A_op45 : array_index_71458[7];
  assign array_update_71462[8] = add_71459 == 32'h0000_0008 ? TestBlock__A_op45 : array_index_71458[8];
  assign array_update_71462[9] = add_71459 == 32'h0000_0009 ? TestBlock__A_op45 : array_index_71458[9];
  assign array_update_71463[0] = add_71461 == 32'h0000_0000 ? TestBlock__B_op45 : array_index_71460[0];
  assign array_update_71463[1] = add_71461 == 32'h0000_0001 ? TestBlock__B_op45 : array_index_71460[1];
  assign array_update_71463[2] = add_71461 == 32'h0000_0002 ? TestBlock__B_op45 : array_index_71460[2];
  assign array_update_71463[3] = add_71461 == 32'h0000_0003 ? TestBlock__B_op45 : array_index_71460[3];
  assign array_update_71463[4] = add_71461 == 32'h0000_0004 ? TestBlock__B_op45 : array_index_71460[4];
  assign array_update_71463[5] = add_71461 == 32'h0000_0005 ? TestBlock__B_op45 : array_index_71460[5];
  assign array_update_71463[6] = add_71461 == 32'h0000_0006 ? TestBlock__B_op45 : array_index_71460[6];
  assign array_update_71463[7] = add_71461 == 32'h0000_0007 ? TestBlock__B_op45 : array_index_71460[7];
  assign array_update_71463[8] = add_71461 == 32'h0000_0008 ? TestBlock__B_op45 : array_index_71460[8];
  assign array_update_71463[9] = add_71461 == 32'h0000_0009 ? TestBlock__B_op45 : array_index_71460[9];
  assign array_update_71464[0] = add_71405 == 32'h0000_0000 ? array_update_71462 : array_update_71454[0];
  assign array_update_71464[1] = add_71405 == 32'h0000_0001 ? array_update_71462 : array_update_71454[1];
  assign array_update_71464[2] = add_71405 == 32'h0000_0002 ? array_update_71462 : array_update_71454[2];
  assign array_update_71464[3] = add_71405 == 32'h0000_0003 ? array_update_71462 : array_update_71454[3];
  assign array_update_71464[4] = add_71405 == 32'h0000_0004 ? array_update_71462 : array_update_71454[4];
  assign array_update_71464[5] = add_71405 == 32'h0000_0005 ? array_update_71462 : array_update_71454[5];
  assign array_update_71464[6] = add_71405 == 32'h0000_0006 ? array_update_71462 : array_update_71454[6];
  assign array_update_71464[7] = add_71405 == 32'h0000_0007 ? array_update_71462 : array_update_71454[7];
  assign array_update_71464[8] = add_71405 == 32'h0000_0008 ? array_update_71462 : array_update_71454[8];
  assign array_update_71464[9] = add_71405 == 32'h0000_0009 ? array_update_71462 : array_update_71454[9];
  assign array_update_71466[0] = add_71407 == 32'h0000_0000 ? array_update_71463 : array_update_71456[0];
  assign array_update_71466[1] = add_71407 == 32'h0000_0001 ? array_update_71463 : array_update_71456[1];
  assign array_update_71466[2] = add_71407 == 32'h0000_0002 ? array_update_71463 : array_update_71456[2];
  assign array_update_71466[3] = add_71407 == 32'h0000_0003 ? array_update_71463 : array_update_71456[3];
  assign array_update_71466[4] = add_71407 == 32'h0000_0004 ? array_update_71463 : array_update_71456[4];
  assign array_update_71466[5] = add_71407 == 32'h0000_0005 ? array_update_71463 : array_update_71456[5];
  assign array_update_71466[6] = add_71407 == 32'h0000_0006 ? array_update_71463 : array_update_71456[6];
  assign array_update_71466[7] = add_71407 == 32'h0000_0007 ? array_update_71463 : array_update_71456[7];
  assign array_update_71466[8] = add_71407 == 32'h0000_0008 ? array_update_71463 : array_update_71456[8];
  assign array_update_71466[9] = add_71407 == 32'h0000_0009 ? array_update_71463 : array_update_71456[9];
  assign array_index_71468 = array_update_71464[add_71405 > 32'h0000_0009 ? 4'h9 : add_71405[3:0]];
  assign add_71469 = add_71459 + 32'h0000_0001;
  assign array_index_71470 = array_update_71466[add_71407 > 32'h0000_0009 ? 4'h9 : add_71407[3:0]];
  assign add_71471 = add_71461 + 32'h0000_0001;
  assign array_update_71472[0] = add_71469 == 32'h0000_0000 ? TestBlock__A_op46 : array_index_71468[0];
  assign array_update_71472[1] = add_71469 == 32'h0000_0001 ? TestBlock__A_op46 : array_index_71468[1];
  assign array_update_71472[2] = add_71469 == 32'h0000_0002 ? TestBlock__A_op46 : array_index_71468[2];
  assign array_update_71472[3] = add_71469 == 32'h0000_0003 ? TestBlock__A_op46 : array_index_71468[3];
  assign array_update_71472[4] = add_71469 == 32'h0000_0004 ? TestBlock__A_op46 : array_index_71468[4];
  assign array_update_71472[5] = add_71469 == 32'h0000_0005 ? TestBlock__A_op46 : array_index_71468[5];
  assign array_update_71472[6] = add_71469 == 32'h0000_0006 ? TestBlock__A_op46 : array_index_71468[6];
  assign array_update_71472[7] = add_71469 == 32'h0000_0007 ? TestBlock__A_op46 : array_index_71468[7];
  assign array_update_71472[8] = add_71469 == 32'h0000_0008 ? TestBlock__A_op46 : array_index_71468[8];
  assign array_update_71472[9] = add_71469 == 32'h0000_0009 ? TestBlock__A_op46 : array_index_71468[9];
  assign array_update_71473[0] = add_71471 == 32'h0000_0000 ? TestBlock__B_op46 : array_index_71470[0];
  assign array_update_71473[1] = add_71471 == 32'h0000_0001 ? TestBlock__B_op46 : array_index_71470[1];
  assign array_update_71473[2] = add_71471 == 32'h0000_0002 ? TestBlock__B_op46 : array_index_71470[2];
  assign array_update_71473[3] = add_71471 == 32'h0000_0003 ? TestBlock__B_op46 : array_index_71470[3];
  assign array_update_71473[4] = add_71471 == 32'h0000_0004 ? TestBlock__B_op46 : array_index_71470[4];
  assign array_update_71473[5] = add_71471 == 32'h0000_0005 ? TestBlock__B_op46 : array_index_71470[5];
  assign array_update_71473[6] = add_71471 == 32'h0000_0006 ? TestBlock__B_op46 : array_index_71470[6];
  assign array_update_71473[7] = add_71471 == 32'h0000_0007 ? TestBlock__B_op46 : array_index_71470[7];
  assign array_update_71473[8] = add_71471 == 32'h0000_0008 ? TestBlock__B_op46 : array_index_71470[8];
  assign array_update_71473[9] = add_71471 == 32'h0000_0009 ? TestBlock__B_op46 : array_index_71470[9];
  assign array_update_71474[0] = add_71405 == 32'h0000_0000 ? array_update_71472 : array_update_71464[0];
  assign array_update_71474[1] = add_71405 == 32'h0000_0001 ? array_update_71472 : array_update_71464[1];
  assign array_update_71474[2] = add_71405 == 32'h0000_0002 ? array_update_71472 : array_update_71464[2];
  assign array_update_71474[3] = add_71405 == 32'h0000_0003 ? array_update_71472 : array_update_71464[3];
  assign array_update_71474[4] = add_71405 == 32'h0000_0004 ? array_update_71472 : array_update_71464[4];
  assign array_update_71474[5] = add_71405 == 32'h0000_0005 ? array_update_71472 : array_update_71464[5];
  assign array_update_71474[6] = add_71405 == 32'h0000_0006 ? array_update_71472 : array_update_71464[6];
  assign array_update_71474[7] = add_71405 == 32'h0000_0007 ? array_update_71472 : array_update_71464[7];
  assign array_update_71474[8] = add_71405 == 32'h0000_0008 ? array_update_71472 : array_update_71464[8];
  assign array_update_71474[9] = add_71405 == 32'h0000_0009 ? array_update_71472 : array_update_71464[9];
  assign array_update_71476[0] = add_71407 == 32'h0000_0000 ? array_update_71473 : array_update_71466[0];
  assign array_update_71476[1] = add_71407 == 32'h0000_0001 ? array_update_71473 : array_update_71466[1];
  assign array_update_71476[2] = add_71407 == 32'h0000_0002 ? array_update_71473 : array_update_71466[2];
  assign array_update_71476[3] = add_71407 == 32'h0000_0003 ? array_update_71473 : array_update_71466[3];
  assign array_update_71476[4] = add_71407 == 32'h0000_0004 ? array_update_71473 : array_update_71466[4];
  assign array_update_71476[5] = add_71407 == 32'h0000_0005 ? array_update_71473 : array_update_71466[5];
  assign array_update_71476[6] = add_71407 == 32'h0000_0006 ? array_update_71473 : array_update_71466[6];
  assign array_update_71476[7] = add_71407 == 32'h0000_0007 ? array_update_71473 : array_update_71466[7];
  assign array_update_71476[8] = add_71407 == 32'h0000_0008 ? array_update_71473 : array_update_71466[8];
  assign array_update_71476[9] = add_71407 == 32'h0000_0009 ? array_update_71473 : array_update_71466[9];
  assign array_index_71478 = array_update_71474[add_71405 > 32'h0000_0009 ? 4'h9 : add_71405[3:0]];
  assign add_71479 = add_71469 + 32'h0000_0001;
  assign array_index_71480 = array_update_71476[add_71407 > 32'h0000_0009 ? 4'h9 : add_71407[3:0]];
  assign add_71481 = add_71471 + 32'h0000_0001;
  assign array_update_71482[0] = add_71479 == 32'h0000_0000 ? TestBlock__A_op47 : array_index_71478[0];
  assign array_update_71482[1] = add_71479 == 32'h0000_0001 ? TestBlock__A_op47 : array_index_71478[1];
  assign array_update_71482[2] = add_71479 == 32'h0000_0002 ? TestBlock__A_op47 : array_index_71478[2];
  assign array_update_71482[3] = add_71479 == 32'h0000_0003 ? TestBlock__A_op47 : array_index_71478[3];
  assign array_update_71482[4] = add_71479 == 32'h0000_0004 ? TestBlock__A_op47 : array_index_71478[4];
  assign array_update_71482[5] = add_71479 == 32'h0000_0005 ? TestBlock__A_op47 : array_index_71478[5];
  assign array_update_71482[6] = add_71479 == 32'h0000_0006 ? TestBlock__A_op47 : array_index_71478[6];
  assign array_update_71482[7] = add_71479 == 32'h0000_0007 ? TestBlock__A_op47 : array_index_71478[7];
  assign array_update_71482[8] = add_71479 == 32'h0000_0008 ? TestBlock__A_op47 : array_index_71478[8];
  assign array_update_71482[9] = add_71479 == 32'h0000_0009 ? TestBlock__A_op47 : array_index_71478[9];
  assign array_update_71483[0] = add_71481 == 32'h0000_0000 ? TestBlock__B_op47 : array_index_71480[0];
  assign array_update_71483[1] = add_71481 == 32'h0000_0001 ? TestBlock__B_op47 : array_index_71480[1];
  assign array_update_71483[2] = add_71481 == 32'h0000_0002 ? TestBlock__B_op47 : array_index_71480[2];
  assign array_update_71483[3] = add_71481 == 32'h0000_0003 ? TestBlock__B_op47 : array_index_71480[3];
  assign array_update_71483[4] = add_71481 == 32'h0000_0004 ? TestBlock__B_op47 : array_index_71480[4];
  assign array_update_71483[5] = add_71481 == 32'h0000_0005 ? TestBlock__B_op47 : array_index_71480[5];
  assign array_update_71483[6] = add_71481 == 32'h0000_0006 ? TestBlock__B_op47 : array_index_71480[6];
  assign array_update_71483[7] = add_71481 == 32'h0000_0007 ? TestBlock__B_op47 : array_index_71480[7];
  assign array_update_71483[8] = add_71481 == 32'h0000_0008 ? TestBlock__B_op47 : array_index_71480[8];
  assign array_update_71483[9] = add_71481 == 32'h0000_0009 ? TestBlock__B_op47 : array_index_71480[9];
  assign array_update_71484[0] = add_71405 == 32'h0000_0000 ? array_update_71482 : array_update_71474[0];
  assign array_update_71484[1] = add_71405 == 32'h0000_0001 ? array_update_71482 : array_update_71474[1];
  assign array_update_71484[2] = add_71405 == 32'h0000_0002 ? array_update_71482 : array_update_71474[2];
  assign array_update_71484[3] = add_71405 == 32'h0000_0003 ? array_update_71482 : array_update_71474[3];
  assign array_update_71484[4] = add_71405 == 32'h0000_0004 ? array_update_71482 : array_update_71474[4];
  assign array_update_71484[5] = add_71405 == 32'h0000_0005 ? array_update_71482 : array_update_71474[5];
  assign array_update_71484[6] = add_71405 == 32'h0000_0006 ? array_update_71482 : array_update_71474[6];
  assign array_update_71484[7] = add_71405 == 32'h0000_0007 ? array_update_71482 : array_update_71474[7];
  assign array_update_71484[8] = add_71405 == 32'h0000_0008 ? array_update_71482 : array_update_71474[8];
  assign array_update_71484[9] = add_71405 == 32'h0000_0009 ? array_update_71482 : array_update_71474[9];
  assign array_update_71486[0] = add_71407 == 32'h0000_0000 ? array_update_71483 : array_update_71476[0];
  assign array_update_71486[1] = add_71407 == 32'h0000_0001 ? array_update_71483 : array_update_71476[1];
  assign array_update_71486[2] = add_71407 == 32'h0000_0002 ? array_update_71483 : array_update_71476[2];
  assign array_update_71486[3] = add_71407 == 32'h0000_0003 ? array_update_71483 : array_update_71476[3];
  assign array_update_71486[4] = add_71407 == 32'h0000_0004 ? array_update_71483 : array_update_71476[4];
  assign array_update_71486[5] = add_71407 == 32'h0000_0005 ? array_update_71483 : array_update_71476[5];
  assign array_update_71486[6] = add_71407 == 32'h0000_0006 ? array_update_71483 : array_update_71476[6];
  assign array_update_71486[7] = add_71407 == 32'h0000_0007 ? array_update_71483 : array_update_71476[7];
  assign array_update_71486[8] = add_71407 == 32'h0000_0008 ? array_update_71483 : array_update_71476[8];
  assign array_update_71486[9] = add_71407 == 32'h0000_0009 ? array_update_71483 : array_update_71476[9];
  assign array_index_71488 = array_update_71484[add_71405 > 32'h0000_0009 ? 4'h9 : add_71405[3:0]];
  assign add_71489 = add_71479 + 32'h0000_0001;
  assign array_index_71490 = array_update_71486[add_71407 > 32'h0000_0009 ? 4'h9 : add_71407[3:0]];
  assign add_71491 = add_71481 + 32'h0000_0001;
  assign array_update_71492[0] = add_71489 == 32'h0000_0000 ? TestBlock__A_op48 : array_index_71488[0];
  assign array_update_71492[1] = add_71489 == 32'h0000_0001 ? TestBlock__A_op48 : array_index_71488[1];
  assign array_update_71492[2] = add_71489 == 32'h0000_0002 ? TestBlock__A_op48 : array_index_71488[2];
  assign array_update_71492[3] = add_71489 == 32'h0000_0003 ? TestBlock__A_op48 : array_index_71488[3];
  assign array_update_71492[4] = add_71489 == 32'h0000_0004 ? TestBlock__A_op48 : array_index_71488[4];
  assign array_update_71492[5] = add_71489 == 32'h0000_0005 ? TestBlock__A_op48 : array_index_71488[5];
  assign array_update_71492[6] = add_71489 == 32'h0000_0006 ? TestBlock__A_op48 : array_index_71488[6];
  assign array_update_71492[7] = add_71489 == 32'h0000_0007 ? TestBlock__A_op48 : array_index_71488[7];
  assign array_update_71492[8] = add_71489 == 32'h0000_0008 ? TestBlock__A_op48 : array_index_71488[8];
  assign array_update_71492[9] = add_71489 == 32'h0000_0009 ? TestBlock__A_op48 : array_index_71488[9];
  assign array_update_71493[0] = add_71491 == 32'h0000_0000 ? TestBlock__B_op48 : array_index_71490[0];
  assign array_update_71493[1] = add_71491 == 32'h0000_0001 ? TestBlock__B_op48 : array_index_71490[1];
  assign array_update_71493[2] = add_71491 == 32'h0000_0002 ? TestBlock__B_op48 : array_index_71490[2];
  assign array_update_71493[3] = add_71491 == 32'h0000_0003 ? TestBlock__B_op48 : array_index_71490[3];
  assign array_update_71493[4] = add_71491 == 32'h0000_0004 ? TestBlock__B_op48 : array_index_71490[4];
  assign array_update_71493[5] = add_71491 == 32'h0000_0005 ? TestBlock__B_op48 : array_index_71490[5];
  assign array_update_71493[6] = add_71491 == 32'h0000_0006 ? TestBlock__B_op48 : array_index_71490[6];
  assign array_update_71493[7] = add_71491 == 32'h0000_0007 ? TestBlock__B_op48 : array_index_71490[7];
  assign array_update_71493[8] = add_71491 == 32'h0000_0008 ? TestBlock__B_op48 : array_index_71490[8];
  assign array_update_71493[9] = add_71491 == 32'h0000_0009 ? TestBlock__B_op48 : array_index_71490[9];
  assign array_update_71494[0] = add_71405 == 32'h0000_0000 ? array_update_71492 : array_update_71484[0];
  assign array_update_71494[1] = add_71405 == 32'h0000_0001 ? array_update_71492 : array_update_71484[1];
  assign array_update_71494[2] = add_71405 == 32'h0000_0002 ? array_update_71492 : array_update_71484[2];
  assign array_update_71494[3] = add_71405 == 32'h0000_0003 ? array_update_71492 : array_update_71484[3];
  assign array_update_71494[4] = add_71405 == 32'h0000_0004 ? array_update_71492 : array_update_71484[4];
  assign array_update_71494[5] = add_71405 == 32'h0000_0005 ? array_update_71492 : array_update_71484[5];
  assign array_update_71494[6] = add_71405 == 32'h0000_0006 ? array_update_71492 : array_update_71484[6];
  assign array_update_71494[7] = add_71405 == 32'h0000_0007 ? array_update_71492 : array_update_71484[7];
  assign array_update_71494[8] = add_71405 == 32'h0000_0008 ? array_update_71492 : array_update_71484[8];
  assign array_update_71494[9] = add_71405 == 32'h0000_0009 ? array_update_71492 : array_update_71484[9];
  assign array_update_71496[0] = add_71407 == 32'h0000_0000 ? array_update_71493 : array_update_71486[0];
  assign array_update_71496[1] = add_71407 == 32'h0000_0001 ? array_update_71493 : array_update_71486[1];
  assign array_update_71496[2] = add_71407 == 32'h0000_0002 ? array_update_71493 : array_update_71486[2];
  assign array_update_71496[3] = add_71407 == 32'h0000_0003 ? array_update_71493 : array_update_71486[3];
  assign array_update_71496[4] = add_71407 == 32'h0000_0004 ? array_update_71493 : array_update_71486[4];
  assign array_update_71496[5] = add_71407 == 32'h0000_0005 ? array_update_71493 : array_update_71486[5];
  assign array_update_71496[6] = add_71407 == 32'h0000_0006 ? array_update_71493 : array_update_71486[6];
  assign array_update_71496[7] = add_71407 == 32'h0000_0007 ? array_update_71493 : array_update_71486[7];
  assign array_update_71496[8] = add_71407 == 32'h0000_0008 ? array_update_71493 : array_update_71486[8];
  assign array_update_71496[9] = add_71407 == 32'h0000_0009 ? array_update_71493 : array_update_71486[9];
  assign array_index_71498 = array_update_71494[add_71405 > 32'h0000_0009 ? 4'h9 : add_71405[3:0]];
  assign add_71499 = add_71489 + 32'h0000_0001;
  assign array_index_71500 = array_update_71496[add_71407 > 32'h0000_0009 ? 4'h9 : add_71407[3:0]];
  assign add_71501 = add_71491 + 32'h0000_0001;
  assign array_update_71502[0] = add_71499 == 32'h0000_0000 ? TestBlock__A_op49 : array_index_71498[0];
  assign array_update_71502[1] = add_71499 == 32'h0000_0001 ? TestBlock__A_op49 : array_index_71498[1];
  assign array_update_71502[2] = add_71499 == 32'h0000_0002 ? TestBlock__A_op49 : array_index_71498[2];
  assign array_update_71502[3] = add_71499 == 32'h0000_0003 ? TestBlock__A_op49 : array_index_71498[3];
  assign array_update_71502[4] = add_71499 == 32'h0000_0004 ? TestBlock__A_op49 : array_index_71498[4];
  assign array_update_71502[5] = add_71499 == 32'h0000_0005 ? TestBlock__A_op49 : array_index_71498[5];
  assign array_update_71502[6] = add_71499 == 32'h0000_0006 ? TestBlock__A_op49 : array_index_71498[6];
  assign array_update_71502[7] = add_71499 == 32'h0000_0007 ? TestBlock__A_op49 : array_index_71498[7];
  assign array_update_71502[8] = add_71499 == 32'h0000_0008 ? TestBlock__A_op49 : array_index_71498[8];
  assign array_update_71502[9] = add_71499 == 32'h0000_0009 ? TestBlock__A_op49 : array_index_71498[9];
  assign array_update_71504[0] = add_71501 == 32'h0000_0000 ? TestBlock__B_op49 : array_index_71500[0];
  assign array_update_71504[1] = add_71501 == 32'h0000_0001 ? TestBlock__B_op49 : array_index_71500[1];
  assign array_update_71504[2] = add_71501 == 32'h0000_0002 ? TestBlock__B_op49 : array_index_71500[2];
  assign array_update_71504[3] = add_71501 == 32'h0000_0003 ? TestBlock__B_op49 : array_index_71500[3];
  assign array_update_71504[4] = add_71501 == 32'h0000_0004 ? TestBlock__B_op49 : array_index_71500[4];
  assign array_update_71504[5] = add_71501 == 32'h0000_0005 ? TestBlock__B_op49 : array_index_71500[5];
  assign array_update_71504[6] = add_71501 == 32'h0000_0006 ? TestBlock__B_op49 : array_index_71500[6];
  assign array_update_71504[7] = add_71501 == 32'h0000_0007 ? TestBlock__B_op49 : array_index_71500[7];
  assign array_update_71504[8] = add_71501 == 32'h0000_0008 ? TestBlock__B_op49 : array_index_71500[8];
  assign array_update_71504[9] = add_71501 == 32'h0000_0009 ? TestBlock__B_op49 : array_index_71500[9];
  assign array_update_71506[0] = add_71405 == 32'h0000_0000 ? array_update_71502 : array_update_71494[0];
  assign array_update_71506[1] = add_71405 == 32'h0000_0001 ? array_update_71502 : array_update_71494[1];
  assign array_update_71506[2] = add_71405 == 32'h0000_0002 ? array_update_71502 : array_update_71494[2];
  assign array_update_71506[3] = add_71405 == 32'h0000_0003 ? array_update_71502 : array_update_71494[3];
  assign array_update_71506[4] = add_71405 == 32'h0000_0004 ? array_update_71502 : array_update_71494[4];
  assign array_update_71506[5] = add_71405 == 32'h0000_0005 ? array_update_71502 : array_update_71494[5];
  assign array_update_71506[6] = add_71405 == 32'h0000_0006 ? array_update_71502 : array_update_71494[6];
  assign array_update_71506[7] = add_71405 == 32'h0000_0007 ? array_update_71502 : array_update_71494[7];
  assign array_update_71506[8] = add_71405 == 32'h0000_0008 ? array_update_71502 : array_update_71494[8];
  assign array_update_71506[9] = add_71405 == 32'h0000_0009 ? array_update_71502 : array_update_71494[9];
  assign add_71507 = add_71405 + 32'h0000_0001;
  assign array_update_71508[0] = add_71407 == 32'h0000_0000 ? array_update_71504 : array_update_71496[0];
  assign array_update_71508[1] = add_71407 == 32'h0000_0001 ? array_update_71504 : array_update_71496[1];
  assign array_update_71508[2] = add_71407 == 32'h0000_0002 ? array_update_71504 : array_update_71496[2];
  assign array_update_71508[3] = add_71407 == 32'h0000_0003 ? array_update_71504 : array_update_71496[3];
  assign array_update_71508[4] = add_71407 == 32'h0000_0004 ? array_update_71504 : array_update_71496[4];
  assign array_update_71508[5] = add_71407 == 32'h0000_0005 ? array_update_71504 : array_update_71496[5];
  assign array_update_71508[6] = add_71407 == 32'h0000_0006 ? array_update_71504 : array_update_71496[6];
  assign array_update_71508[7] = add_71407 == 32'h0000_0007 ? array_update_71504 : array_update_71496[7];
  assign array_update_71508[8] = add_71407 == 32'h0000_0008 ? array_update_71504 : array_update_71496[8];
  assign array_update_71508[9] = add_71407 == 32'h0000_0009 ? array_update_71504 : array_update_71496[9];
  assign add_71509 = add_71407 + 32'h0000_0001;
  assign array_index_71510 = array_update_71506[add_71507 > 32'h0000_0009 ? 4'h9 : add_71507[3:0]];
  assign literal_71511 = 32'h0000_0000;
  assign array_index_71512 = array_update_71508[add_71509 > 32'h0000_0009 ? 4'h9 : add_71509[3:0]];
  assign literal_71513 = 32'h0000_0000;
  assign array_update_71514[0] = literal_71511 == 32'h0000_0000 ? TestBlock__A_op50 : array_index_71510[0];
  assign array_update_71514[1] = literal_71511 == 32'h0000_0001 ? TestBlock__A_op50 : array_index_71510[1];
  assign array_update_71514[2] = literal_71511 == 32'h0000_0002 ? TestBlock__A_op50 : array_index_71510[2];
  assign array_update_71514[3] = literal_71511 == 32'h0000_0003 ? TestBlock__A_op50 : array_index_71510[3];
  assign array_update_71514[4] = literal_71511 == 32'h0000_0004 ? TestBlock__A_op50 : array_index_71510[4];
  assign array_update_71514[5] = literal_71511 == 32'h0000_0005 ? TestBlock__A_op50 : array_index_71510[5];
  assign array_update_71514[6] = literal_71511 == 32'h0000_0006 ? TestBlock__A_op50 : array_index_71510[6];
  assign array_update_71514[7] = literal_71511 == 32'h0000_0007 ? TestBlock__A_op50 : array_index_71510[7];
  assign array_update_71514[8] = literal_71511 == 32'h0000_0008 ? TestBlock__A_op50 : array_index_71510[8];
  assign array_update_71514[9] = literal_71511 == 32'h0000_0009 ? TestBlock__A_op50 : array_index_71510[9];
  assign array_update_71515[0] = literal_71513 == 32'h0000_0000 ? TestBlock__B_op50 : array_index_71512[0];
  assign array_update_71515[1] = literal_71513 == 32'h0000_0001 ? TestBlock__B_op50 : array_index_71512[1];
  assign array_update_71515[2] = literal_71513 == 32'h0000_0002 ? TestBlock__B_op50 : array_index_71512[2];
  assign array_update_71515[3] = literal_71513 == 32'h0000_0003 ? TestBlock__B_op50 : array_index_71512[3];
  assign array_update_71515[4] = literal_71513 == 32'h0000_0004 ? TestBlock__B_op50 : array_index_71512[4];
  assign array_update_71515[5] = literal_71513 == 32'h0000_0005 ? TestBlock__B_op50 : array_index_71512[5];
  assign array_update_71515[6] = literal_71513 == 32'h0000_0006 ? TestBlock__B_op50 : array_index_71512[6];
  assign array_update_71515[7] = literal_71513 == 32'h0000_0007 ? TestBlock__B_op50 : array_index_71512[7];
  assign array_update_71515[8] = literal_71513 == 32'h0000_0008 ? TestBlock__B_op50 : array_index_71512[8];
  assign array_update_71515[9] = literal_71513 == 32'h0000_0009 ? TestBlock__B_op50 : array_index_71512[9];
  assign array_update_71516[0] = add_71507 == 32'h0000_0000 ? array_update_71514 : array_update_71506[0];
  assign array_update_71516[1] = add_71507 == 32'h0000_0001 ? array_update_71514 : array_update_71506[1];
  assign array_update_71516[2] = add_71507 == 32'h0000_0002 ? array_update_71514 : array_update_71506[2];
  assign array_update_71516[3] = add_71507 == 32'h0000_0003 ? array_update_71514 : array_update_71506[3];
  assign array_update_71516[4] = add_71507 == 32'h0000_0004 ? array_update_71514 : array_update_71506[4];
  assign array_update_71516[5] = add_71507 == 32'h0000_0005 ? array_update_71514 : array_update_71506[5];
  assign array_update_71516[6] = add_71507 == 32'h0000_0006 ? array_update_71514 : array_update_71506[6];
  assign array_update_71516[7] = add_71507 == 32'h0000_0007 ? array_update_71514 : array_update_71506[7];
  assign array_update_71516[8] = add_71507 == 32'h0000_0008 ? array_update_71514 : array_update_71506[8];
  assign array_update_71516[9] = add_71507 == 32'h0000_0009 ? array_update_71514 : array_update_71506[9];
  assign array_update_71518[0] = add_71509 == 32'h0000_0000 ? array_update_71515 : array_update_71508[0];
  assign array_update_71518[1] = add_71509 == 32'h0000_0001 ? array_update_71515 : array_update_71508[1];
  assign array_update_71518[2] = add_71509 == 32'h0000_0002 ? array_update_71515 : array_update_71508[2];
  assign array_update_71518[3] = add_71509 == 32'h0000_0003 ? array_update_71515 : array_update_71508[3];
  assign array_update_71518[4] = add_71509 == 32'h0000_0004 ? array_update_71515 : array_update_71508[4];
  assign array_update_71518[5] = add_71509 == 32'h0000_0005 ? array_update_71515 : array_update_71508[5];
  assign array_update_71518[6] = add_71509 == 32'h0000_0006 ? array_update_71515 : array_update_71508[6];
  assign array_update_71518[7] = add_71509 == 32'h0000_0007 ? array_update_71515 : array_update_71508[7];
  assign array_update_71518[8] = add_71509 == 32'h0000_0008 ? array_update_71515 : array_update_71508[8];
  assign array_update_71518[9] = add_71509 == 32'h0000_0009 ? array_update_71515 : array_update_71508[9];
  assign array_index_71520 = array_update_71516[add_71507 > 32'h0000_0009 ? 4'h9 : add_71507[3:0]];
  assign add_71521 = literal_71511 + 32'h0000_0001;
  assign array_index_71522 = array_update_71518[add_71509 > 32'h0000_0009 ? 4'h9 : add_71509[3:0]];
  assign add_71523 = literal_71513 + 32'h0000_0001;
  assign array_update_71524[0] = add_71521 == 32'h0000_0000 ? TestBlock__A_op51 : array_index_71520[0];
  assign array_update_71524[1] = add_71521 == 32'h0000_0001 ? TestBlock__A_op51 : array_index_71520[1];
  assign array_update_71524[2] = add_71521 == 32'h0000_0002 ? TestBlock__A_op51 : array_index_71520[2];
  assign array_update_71524[3] = add_71521 == 32'h0000_0003 ? TestBlock__A_op51 : array_index_71520[3];
  assign array_update_71524[4] = add_71521 == 32'h0000_0004 ? TestBlock__A_op51 : array_index_71520[4];
  assign array_update_71524[5] = add_71521 == 32'h0000_0005 ? TestBlock__A_op51 : array_index_71520[5];
  assign array_update_71524[6] = add_71521 == 32'h0000_0006 ? TestBlock__A_op51 : array_index_71520[6];
  assign array_update_71524[7] = add_71521 == 32'h0000_0007 ? TestBlock__A_op51 : array_index_71520[7];
  assign array_update_71524[8] = add_71521 == 32'h0000_0008 ? TestBlock__A_op51 : array_index_71520[8];
  assign array_update_71524[9] = add_71521 == 32'h0000_0009 ? TestBlock__A_op51 : array_index_71520[9];
  assign array_update_71525[0] = add_71523 == 32'h0000_0000 ? TestBlock__B_op51 : array_index_71522[0];
  assign array_update_71525[1] = add_71523 == 32'h0000_0001 ? TestBlock__B_op51 : array_index_71522[1];
  assign array_update_71525[2] = add_71523 == 32'h0000_0002 ? TestBlock__B_op51 : array_index_71522[2];
  assign array_update_71525[3] = add_71523 == 32'h0000_0003 ? TestBlock__B_op51 : array_index_71522[3];
  assign array_update_71525[4] = add_71523 == 32'h0000_0004 ? TestBlock__B_op51 : array_index_71522[4];
  assign array_update_71525[5] = add_71523 == 32'h0000_0005 ? TestBlock__B_op51 : array_index_71522[5];
  assign array_update_71525[6] = add_71523 == 32'h0000_0006 ? TestBlock__B_op51 : array_index_71522[6];
  assign array_update_71525[7] = add_71523 == 32'h0000_0007 ? TestBlock__B_op51 : array_index_71522[7];
  assign array_update_71525[8] = add_71523 == 32'h0000_0008 ? TestBlock__B_op51 : array_index_71522[8];
  assign array_update_71525[9] = add_71523 == 32'h0000_0009 ? TestBlock__B_op51 : array_index_71522[9];
  assign array_update_71526[0] = add_71507 == 32'h0000_0000 ? array_update_71524 : array_update_71516[0];
  assign array_update_71526[1] = add_71507 == 32'h0000_0001 ? array_update_71524 : array_update_71516[1];
  assign array_update_71526[2] = add_71507 == 32'h0000_0002 ? array_update_71524 : array_update_71516[2];
  assign array_update_71526[3] = add_71507 == 32'h0000_0003 ? array_update_71524 : array_update_71516[3];
  assign array_update_71526[4] = add_71507 == 32'h0000_0004 ? array_update_71524 : array_update_71516[4];
  assign array_update_71526[5] = add_71507 == 32'h0000_0005 ? array_update_71524 : array_update_71516[5];
  assign array_update_71526[6] = add_71507 == 32'h0000_0006 ? array_update_71524 : array_update_71516[6];
  assign array_update_71526[7] = add_71507 == 32'h0000_0007 ? array_update_71524 : array_update_71516[7];
  assign array_update_71526[8] = add_71507 == 32'h0000_0008 ? array_update_71524 : array_update_71516[8];
  assign array_update_71526[9] = add_71507 == 32'h0000_0009 ? array_update_71524 : array_update_71516[9];
  assign array_update_71528[0] = add_71509 == 32'h0000_0000 ? array_update_71525 : array_update_71518[0];
  assign array_update_71528[1] = add_71509 == 32'h0000_0001 ? array_update_71525 : array_update_71518[1];
  assign array_update_71528[2] = add_71509 == 32'h0000_0002 ? array_update_71525 : array_update_71518[2];
  assign array_update_71528[3] = add_71509 == 32'h0000_0003 ? array_update_71525 : array_update_71518[3];
  assign array_update_71528[4] = add_71509 == 32'h0000_0004 ? array_update_71525 : array_update_71518[4];
  assign array_update_71528[5] = add_71509 == 32'h0000_0005 ? array_update_71525 : array_update_71518[5];
  assign array_update_71528[6] = add_71509 == 32'h0000_0006 ? array_update_71525 : array_update_71518[6];
  assign array_update_71528[7] = add_71509 == 32'h0000_0007 ? array_update_71525 : array_update_71518[7];
  assign array_update_71528[8] = add_71509 == 32'h0000_0008 ? array_update_71525 : array_update_71518[8];
  assign array_update_71528[9] = add_71509 == 32'h0000_0009 ? array_update_71525 : array_update_71518[9];
  assign array_index_71530 = array_update_71526[add_71507 > 32'h0000_0009 ? 4'h9 : add_71507[3:0]];
  assign add_71531 = add_71521 + 32'h0000_0001;
  assign array_index_71532 = array_update_71528[add_71509 > 32'h0000_0009 ? 4'h9 : add_71509[3:0]];
  assign add_71533 = add_71523 + 32'h0000_0001;
  assign array_update_71534[0] = add_71531 == 32'h0000_0000 ? TestBlock__A_op52 : array_index_71530[0];
  assign array_update_71534[1] = add_71531 == 32'h0000_0001 ? TestBlock__A_op52 : array_index_71530[1];
  assign array_update_71534[2] = add_71531 == 32'h0000_0002 ? TestBlock__A_op52 : array_index_71530[2];
  assign array_update_71534[3] = add_71531 == 32'h0000_0003 ? TestBlock__A_op52 : array_index_71530[3];
  assign array_update_71534[4] = add_71531 == 32'h0000_0004 ? TestBlock__A_op52 : array_index_71530[4];
  assign array_update_71534[5] = add_71531 == 32'h0000_0005 ? TestBlock__A_op52 : array_index_71530[5];
  assign array_update_71534[6] = add_71531 == 32'h0000_0006 ? TestBlock__A_op52 : array_index_71530[6];
  assign array_update_71534[7] = add_71531 == 32'h0000_0007 ? TestBlock__A_op52 : array_index_71530[7];
  assign array_update_71534[8] = add_71531 == 32'h0000_0008 ? TestBlock__A_op52 : array_index_71530[8];
  assign array_update_71534[9] = add_71531 == 32'h0000_0009 ? TestBlock__A_op52 : array_index_71530[9];
  assign array_update_71535[0] = add_71533 == 32'h0000_0000 ? TestBlock__B_op52 : array_index_71532[0];
  assign array_update_71535[1] = add_71533 == 32'h0000_0001 ? TestBlock__B_op52 : array_index_71532[1];
  assign array_update_71535[2] = add_71533 == 32'h0000_0002 ? TestBlock__B_op52 : array_index_71532[2];
  assign array_update_71535[3] = add_71533 == 32'h0000_0003 ? TestBlock__B_op52 : array_index_71532[3];
  assign array_update_71535[4] = add_71533 == 32'h0000_0004 ? TestBlock__B_op52 : array_index_71532[4];
  assign array_update_71535[5] = add_71533 == 32'h0000_0005 ? TestBlock__B_op52 : array_index_71532[5];
  assign array_update_71535[6] = add_71533 == 32'h0000_0006 ? TestBlock__B_op52 : array_index_71532[6];
  assign array_update_71535[7] = add_71533 == 32'h0000_0007 ? TestBlock__B_op52 : array_index_71532[7];
  assign array_update_71535[8] = add_71533 == 32'h0000_0008 ? TestBlock__B_op52 : array_index_71532[8];
  assign array_update_71535[9] = add_71533 == 32'h0000_0009 ? TestBlock__B_op52 : array_index_71532[9];
  assign array_update_71536[0] = add_71507 == 32'h0000_0000 ? array_update_71534 : array_update_71526[0];
  assign array_update_71536[1] = add_71507 == 32'h0000_0001 ? array_update_71534 : array_update_71526[1];
  assign array_update_71536[2] = add_71507 == 32'h0000_0002 ? array_update_71534 : array_update_71526[2];
  assign array_update_71536[3] = add_71507 == 32'h0000_0003 ? array_update_71534 : array_update_71526[3];
  assign array_update_71536[4] = add_71507 == 32'h0000_0004 ? array_update_71534 : array_update_71526[4];
  assign array_update_71536[5] = add_71507 == 32'h0000_0005 ? array_update_71534 : array_update_71526[5];
  assign array_update_71536[6] = add_71507 == 32'h0000_0006 ? array_update_71534 : array_update_71526[6];
  assign array_update_71536[7] = add_71507 == 32'h0000_0007 ? array_update_71534 : array_update_71526[7];
  assign array_update_71536[8] = add_71507 == 32'h0000_0008 ? array_update_71534 : array_update_71526[8];
  assign array_update_71536[9] = add_71507 == 32'h0000_0009 ? array_update_71534 : array_update_71526[9];
  assign array_update_71538[0] = add_71509 == 32'h0000_0000 ? array_update_71535 : array_update_71528[0];
  assign array_update_71538[1] = add_71509 == 32'h0000_0001 ? array_update_71535 : array_update_71528[1];
  assign array_update_71538[2] = add_71509 == 32'h0000_0002 ? array_update_71535 : array_update_71528[2];
  assign array_update_71538[3] = add_71509 == 32'h0000_0003 ? array_update_71535 : array_update_71528[3];
  assign array_update_71538[4] = add_71509 == 32'h0000_0004 ? array_update_71535 : array_update_71528[4];
  assign array_update_71538[5] = add_71509 == 32'h0000_0005 ? array_update_71535 : array_update_71528[5];
  assign array_update_71538[6] = add_71509 == 32'h0000_0006 ? array_update_71535 : array_update_71528[6];
  assign array_update_71538[7] = add_71509 == 32'h0000_0007 ? array_update_71535 : array_update_71528[7];
  assign array_update_71538[8] = add_71509 == 32'h0000_0008 ? array_update_71535 : array_update_71528[8];
  assign array_update_71538[9] = add_71509 == 32'h0000_0009 ? array_update_71535 : array_update_71528[9];
  assign array_index_71540 = array_update_71536[add_71507 > 32'h0000_0009 ? 4'h9 : add_71507[3:0]];
  assign add_71541 = add_71531 + 32'h0000_0001;
  assign array_index_71542 = array_update_71538[add_71509 > 32'h0000_0009 ? 4'h9 : add_71509[3:0]];
  assign add_71543 = add_71533 + 32'h0000_0001;
  assign array_update_71544[0] = add_71541 == 32'h0000_0000 ? TestBlock__A_op53 : array_index_71540[0];
  assign array_update_71544[1] = add_71541 == 32'h0000_0001 ? TestBlock__A_op53 : array_index_71540[1];
  assign array_update_71544[2] = add_71541 == 32'h0000_0002 ? TestBlock__A_op53 : array_index_71540[2];
  assign array_update_71544[3] = add_71541 == 32'h0000_0003 ? TestBlock__A_op53 : array_index_71540[3];
  assign array_update_71544[4] = add_71541 == 32'h0000_0004 ? TestBlock__A_op53 : array_index_71540[4];
  assign array_update_71544[5] = add_71541 == 32'h0000_0005 ? TestBlock__A_op53 : array_index_71540[5];
  assign array_update_71544[6] = add_71541 == 32'h0000_0006 ? TestBlock__A_op53 : array_index_71540[6];
  assign array_update_71544[7] = add_71541 == 32'h0000_0007 ? TestBlock__A_op53 : array_index_71540[7];
  assign array_update_71544[8] = add_71541 == 32'h0000_0008 ? TestBlock__A_op53 : array_index_71540[8];
  assign array_update_71544[9] = add_71541 == 32'h0000_0009 ? TestBlock__A_op53 : array_index_71540[9];
  assign array_update_71545[0] = add_71543 == 32'h0000_0000 ? TestBlock__B_op53 : array_index_71542[0];
  assign array_update_71545[1] = add_71543 == 32'h0000_0001 ? TestBlock__B_op53 : array_index_71542[1];
  assign array_update_71545[2] = add_71543 == 32'h0000_0002 ? TestBlock__B_op53 : array_index_71542[2];
  assign array_update_71545[3] = add_71543 == 32'h0000_0003 ? TestBlock__B_op53 : array_index_71542[3];
  assign array_update_71545[4] = add_71543 == 32'h0000_0004 ? TestBlock__B_op53 : array_index_71542[4];
  assign array_update_71545[5] = add_71543 == 32'h0000_0005 ? TestBlock__B_op53 : array_index_71542[5];
  assign array_update_71545[6] = add_71543 == 32'h0000_0006 ? TestBlock__B_op53 : array_index_71542[6];
  assign array_update_71545[7] = add_71543 == 32'h0000_0007 ? TestBlock__B_op53 : array_index_71542[7];
  assign array_update_71545[8] = add_71543 == 32'h0000_0008 ? TestBlock__B_op53 : array_index_71542[8];
  assign array_update_71545[9] = add_71543 == 32'h0000_0009 ? TestBlock__B_op53 : array_index_71542[9];
  assign array_update_71546[0] = add_71507 == 32'h0000_0000 ? array_update_71544 : array_update_71536[0];
  assign array_update_71546[1] = add_71507 == 32'h0000_0001 ? array_update_71544 : array_update_71536[1];
  assign array_update_71546[2] = add_71507 == 32'h0000_0002 ? array_update_71544 : array_update_71536[2];
  assign array_update_71546[3] = add_71507 == 32'h0000_0003 ? array_update_71544 : array_update_71536[3];
  assign array_update_71546[4] = add_71507 == 32'h0000_0004 ? array_update_71544 : array_update_71536[4];
  assign array_update_71546[5] = add_71507 == 32'h0000_0005 ? array_update_71544 : array_update_71536[5];
  assign array_update_71546[6] = add_71507 == 32'h0000_0006 ? array_update_71544 : array_update_71536[6];
  assign array_update_71546[7] = add_71507 == 32'h0000_0007 ? array_update_71544 : array_update_71536[7];
  assign array_update_71546[8] = add_71507 == 32'h0000_0008 ? array_update_71544 : array_update_71536[8];
  assign array_update_71546[9] = add_71507 == 32'h0000_0009 ? array_update_71544 : array_update_71536[9];
  assign array_update_71548[0] = add_71509 == 32'h0000_0000 ? array_update_71545 : array_update_71538[0];
  assign array_update_71548[1] = add_71509 == 32'h0000_0001 ? array_update_71545 : array_update_71538[1];
  assign array_update_71548[2] = add_71509 == 32'h0000_0002 ? array_update_71545 : array_update_71538[2];
  assign array_update_71548[3] = add_71509 == 32'h0000_0003 ? array_update_71545 : array_update_71538[3];
  assign array_update_71548[4] = add_71509 == 32'h0000_0004 ? array_update_71545 : array_update_71538[4];
  assign array_update_71548[5] = add_71509 == 32'h0000_0005 ? array_update_71545 : array_update_71538[5];
  assign array_update_71548[6] = add_71509 == 32'h0000_0006 ? array_update_71545 : array_update_71538[6];
  assign array_update_71548[7] = add_71509 == 32'h0000_0007 ? array_update_71545 : array_update_71538[7];
  assign array_update_71548[8] = add_71509 == 32'h0000_0008 ? array_update_71545 : array_update_71538[8];
  assign array_update_71548[9] = add_71509 == 32'h0000_0009 ? array_update_71545 : array_update_71538[9];
  assign array_index_71550 = array_update_71546[add_71507 > 32'h0000_0009 ? 4'h9 : add_71507[3:0]];
  assign add_71551 = add_71541 + 32'h0000_0001;
  assign array_index_71552 = array_update_71548[add_71509 > 32'h0000_0009 ? 4'h9 : add_71509[3:0]];
  assign add_71553 = add_71543 + 32'h0000_0001;
  assign array_update_71554[0] = add_71551 == 32'h0000_0000 ? TestBlock__A_op54 : array_index_71550[0];
  assign array_update_71554[1] = add_71551 == 32'h0000_0001 ? TestBlock__A_op54 : array_index_71550[1];
  assign array_update_71554[2] = add_71551 == 32'h0000_0002 ? TestBlock__A_op54 : array_index_71550[2];
  assign array_update_71554[3] = add_71551 == 32'h0000_0003 ? TestBlock__A_op54 : array_index_71550[3];
  assign array_update_71554[4] = add_71551 == 32'h0000_0004 ? TestBlock__A_op54 : array_index_71550[4];
  assign array_update_71554[5] = add_71551 == 32'h0000_0005 ? TestBlock__A_op54 : array_index_71550[5];
  assign array_update_71554[6] = add_71551 == 32'h0000_0006 ? TestBlock__A_op54 : array_index_71550[6];
  assign array_update_71554[7] = add_71551 == 32'h0000_0007 ? TestBlock__A_op54 : array_index_71550[7];
  assign array_update_71554[8] = add_71551 == 32'h0000_0008 ? TestBlock__A_op54 : array_index_71550[8];
  assign array_update_71554[9] = add_71551 == 32'h0000_0009 ? TestBlock__A_op54 : array_index_71550[9];
  assign array_update_71555[0] = add_71553 == 32'h0000_0000 ? TestBlock__B_op54 : array_index_71552[0];
  assign array_update_71555[1] = add_71553 == 32'h0000_0001 ? TestBlock__B_op54 : array_index_71552[1];
  assign array_update_71555[2] = add_71553 == 32'h0000_0002 ? TestBlock__B_op54 : array_index_71552[2];
  assign array_update_71555[3] = add_71553 == 32'h0000_0003 ? TestBlock__B_op54 : array_index_71552[3];
  assign array_update_71555[4] = add_71553 == 32'h0000_0004 ? TestBlock__B_op54 : array_index_71552[4];
  assign array_update_71555[5] = add_71553 == 32'h0000_0005 ? TestBlock__B_op54 : array_index_71552[5];
  assign array_update_71555[6] = add_71553 == 32'h0000_0006 ? TestBlock__B_op54 : array_index_71552[6];
  assign array_update_71555[7] = add_71553 == 32'h0000_0007 ? TestBlock__B_op54 : array_index_71552[7];
  assign array_update_71555[8] = add_71553 == 32'h0000_0008 ? TestBlock__B_op54 : array_index_71552[8];
  assign array_update_71555[9] = add_71553 == 32'h0000_0009 ? TestBlock__B_op54 : array_index_71552[9];
  assign array_update_71556[0] = add_71507 == 32'h0000_0000 ? array_update_71554 : array_update_71546[0];
  assign array_update_71556[1] = add_71507 == 32'h0000_0001 ? array_update_71554 : array_update_71546[1];
  assign array_update_71556[2] = add_71507 == 32'h0000_0002 ? array_update_71554 : array_update_71546[2];
  assign array_update_71556[3] = add_71507 == 32'h0000_0003 ? array_update_71554 : array_update_71546[3];
  assign array_update_71556[4] = add_71507 == 32'h0000_0004 ? array_update_71554 : array_update_71546[4];
  assign array_update_71556[5] = add_71507 == 32'h0000_0005 ? array_update_71554 : array_update_71546[5];
  assign array_update_71556[6] = add_71507 == 32'h0000_0006 ? array_update_71554 : array_update_71546[6];
  assign array_update_71556[7] = add_71507 == 32'h0000_0007 ? array_update_71554 : array_update_71546[7];
  assign array_update_71556[8] = add_71507 == 32'h0000_0008 ? array_update_71554 : array_update_71546[8];
  assign array_update_71556[9] = add_71507 == 32'h0000_0009 ? array_update_71554 : array_update_71546[9];
  assign array_update_71558[0] = add_71509 == 32'h0000_0000 ? array_update_71555 : array_update_71548[0];
  assign array_update_71558[1] = add_71509 == 32'h0000_0001 ? array_update_71555 : array_update_71548[1];
  assign array_update_71558[2] = add_71509 == 32'h0000_0002 ? array_update_71555 : array_update_71548[2];
  assign array_update_71558[3] = add_71509 == 32'h0000_0003 ? array_update_71555 : array_update_71548[3];
  assign array_update_71558[4] = add_71509 == 32'h0000_0004 ? array_update_71555 : array_update_71548[4];
  assign array_update_71558[5] = add_71509 == 32'h0000_0005 ? array_update_71555 : array_update_71548[5];
  assign array_update_71558[6] = add_71509 == 32'h0000_0006 ? array_update_71555 : array_update_71548[6];
  assign array_update_71558[7] = add_71509 == 32'h0000_0007 ? array_update_71555 : array_update_71548[7];
  assign array_update_71558[8] = add_71509 == 32'h0000_0008 ? array_update_71555 : array_update_71548[8];
  assign array_update_71558[9] = add_71509 == 32'h0000_0009 ? array_update_71555 : array_update_71548[9];
  assign array_index_71560 = array_update_71556[add_71507 > 32'h0000_0009 ? 4'h9 : add_71507[3:0]];
  assign add_71561 = add_71551 + 32'h0000_0001;
  assign array_index_71562 = array_update_71558[add_71509 > 32'h0000_0009 ? 4'h9 : add_71509[3:0]];
  assign add_71563 = add_71553 + 32'h0000_0001;
  assign array_update_71564[0] = add_71561 == 32'h0000_0000 ? TestBlock__A_op55 : array_index_71560[0];
  assign array_update_71564[1] = add_71561 == 32'h0000_0001 ? TestBlock__A_op55 : array_index_71560[1];
  assign array_update_71564[2] = add_71561 == 32'h0000_0002 ? TestBlock__A_op55 : array_index_71560[2];
  assign array_update_71564[3] = add_71561 == 32'h0000_0003 ? TestBlock__A_op55 : array_index_71560[3];
  assign array_update_71564[4] = add_71561 == 32'h0000_0004 ? TestBlock__A_op55 : array_index_71560[4];
  assign array_update_71564[5] = add_71561 == 32'h0000_0005 ? TestBlock__A_op55 : array_index_71560[5];
  assign array_update_71564[6] = add_71561 == 32'h0000_0006 ? TestBlock__A_op55 : array_index_71560[6];
  assign array_update_71564[7] = add_71561 == 32'h0000_0007 ? TestBlock__A_op55 : array_index_71560[7];
  assign array_update_71564[8] = add_71561 == 32'h0000_0008 ? TestBlock__A_op55 : array_index_71560[8];
  assign array_update_71564[9] = add_71561 == 32'h0000_0009 ? TestBlock__A_op55 : array_index_71560[9];
  assign array_update_71565[0] = add_71563 == 32'h0000_0000 ? TestBlock__B_op55 : array_index_71562[0];
  assign array_update_71565[1] = add_71563 == 32'h0000_0001 ? TestBlock__B_op55 : array_index_71562[1];
  assign array_update_71565[2] = add_71563 == 32'h0000_0002 ? TestBlock__B_op55 : array_index_71562[2];
  assign array_update_71565[3] = add_71563 == 32'h0000_0003 ? TestBlock__B_op55 : array_index_71562[3];
  assign array_update_71565[4] = add_71563 == 32'h0000_0004 ? TestBlock__B_op55 : array_index_71562[4];
  assign array_update_71565[5] = add_71563 == 32'h0000_0005 ? TestBlock__B_op55 : array_index_71562[5];
  assign array_update_71565[6] = add_71563 == 32'h0000_0006 ? TestBlock__B_op55 : array_index_71562[6];
  assign array_update_71565[7] = add_71563 == 32'h0000_0007 ? TestBlock__B_op55 : array_index_71562[7];
  assign array_update_71565[8] = add_71563 == 32'h0000_0008 ? TestBlock__B_op55 : array_index_71562[8];
  assign array_update_71565[9] = add_71563 == 32'h0000_0009 ? TestBlock__B_op55 : array_index_71562[9];
  assign array_update_71566[0] = add_71507 == 32'h0000_0000 ? array_update_71564 : array_update_71556[0];
  assign array_update_71566[1] = add_71507 == 32'h0000_0001 ? array_update_71564 : array_update_71556[1];
  assign array_update_71566[2] = add_71507 == 32'h0000_0002 ? array_update_71564 : array_update_71556[2];
  assign array_update_71566[3] = add_71507 == 32'h0000_0003 ? array_update_71564 : array_update_71556[3];
  assign array_update_71566[4] = add_71507 == 32'h0000_0004 ? array_update_71564 : array_update_71556[4];
  assign array_update_71566[5] = add_71507 == 32'h0000_0005 ? array_update_71564 : array_update_71556[5];
  assign array_update_71566[6] = add_71507 == 32'h0000_0006 ? array_update_71564 : array_update_71556[6];
  assign array_update_71566[7] = add_71507 == 32'h0000_0007 ? array_update_71564 : array_update_71556[7];
  assign array_update_71566[8] = add_71507 == 32'h0000_0008 ? array_update_71564 : array_update_71556[8];
  assign array_update_71566[9] = add_71507 == 32'h0000_0009 ? array_update_71564 : array_update_71556[9];
  assign array_update_71568[0] = add_71509 == 32'h0000_0000 ? array_update_71565 : array_update_71558[0];
  assign array_update_71568[1] = add_71509 == 32'h0000_0001 ? array_update_71565 : array_update_71558[1];
  assign array_update_71568[2] = add_71509 == 32'h0000_0002 ? array_update_71565 : array_update_71558[2];
  assign array_update_71568[3] = add_71509 == 32'h0000_0003 ? array_update_71565 : array_update_71558[3];
  assign array_update_71568[4] = add_71509 == 32'h0000_0004 ? array_update_71565 : array_update_71558[4];
  assign array_update_71568[5] = add_71509 == 32'h0000_0005 ? array_update_71565 : array_update_71558[5];
  assign array_update_71568[6] = add_71509 == 32'h0000_0006 ? array_update_71565 : array_update_71558[6];
  assign array_update_71568[7] = add_71509 == 32'h0000_0007 ? array_update_71565 : array_update_71558[7];
  assign array_update_71568[8] = add_71509 == 32'h0000_0008 ? array_update_71565 : array_update_71558[8];
  assign array_update_71568[9] = add_71509 == 32'h0000_0009 ? array_update_71565 : array_update_71558[9];
  assign array_index_71570 = array_update_71566[add_71507 > 32'h0000_0009 ? 4'h9 : add_71507[3:0]];
  assign add_71571 = add_71561 + 32'h0000_0001;
  assign array_index_71572 = array_update_71568[add_71509 > 32'h0000_0009 ? 4'h9 : add_71509[3:0]];
  assign add_71573 = add_71563 + 32'h0000_0001;
  assign array_update_71574[0] = add_71571 == 32'h0000_0000 ? TestBlock__A_op56 : array_index_71570[0];
  assign array_update_71574[1] = add_71571 == 32'h0000_0001 ? TestBlock__A_op56 : array_index_71570[1];
  assign array_update_71574[2] = add_71571 == 32'h0000_0002 ? TestBlock__A_op56 : array_index_71570[2];
  assign array_update_71574[3] = add_71571 == 32'h0000_0003 ? TestBlock__A_op56 : array_index_71570[3];
  assign array_update_71574[4] = add_71571 == 32'h0000_0004 ? TestBlock__A_op56 : array_index_71570[4];
  assign array_update_71574[5] = add_71571 == 32'h0000_0005 ? TestBlock__A_op56 : array_index_71570[5];
  assign array_update_71574[6] = add_71571 == 32'h0000_0006 ? TestBlock__A_op56 : array_index_71570[6];
  assign array_update_71574[7] = add_71571 == 32'h0000_0007 ? TestBlock__A_op56 : array_index_71570[7];
  assign array_update_71574[8] = add_71571 == 32'h0000_0008 ? TestBlock__A_op56 : array_index_71570[8];
  assign array_update_71574[9] = add_71571 == 32'h0000_0009 ? TestBlock__A_op56 : array_index_71570[9];
  assign array_update_71575[0] = add_71573 == 32'h0000_0000 ? TestBlock__B_op56 : array_index_71572[0];
  assign array_update_71575[1] = add_71573 == 32'h0000_0001 ? TestBlock__B_op56 : array_index_71572[1];
  assign array_update_71575[2] = add_71573 == 32'h0000_0002 ? TestBlock__B_op56 : array_index_71572[2];
  assign array_update_71575[3] = add_71573 == 32'h0000_0003 ? TestBlock__B_op56 : array_index_71572[3];
  assign array_update_71575[4] = add_71573 == 32'h0000_0004 ? TestBlock__B_op56 : array_index_71572[4];
  assign array_update_71575[5] = add_71573 == 32'h0000_0005 ? TestBlock__B_op56 : array_index_71572[5];
  assign array_update_71575[6] = add_71573 == 32'h0000_0006 ? TestBlock__B_op56 : array_index_71572[6];
  assign array_update_71575[7] = add_71573 == 32'h0000_0007 ? TestBlock__B_op56 : array_index_71572[7];
  assign array_update_71575[8] = add_71573 == 32'h0000_0008 ? TestBlock__B_op56 : array_index_71572[8];
  assign array_update_71575[9] = add_71573 == 32'h0000_0009 ? TestBlock__B_op56 : array_index_71572[9];
  assign array_update_71576[0] = add_71507 == 32'h0000_0000 ? array_update_71574 : array_update_71566[0];
  assign array_update_71576[1] = add_71507 == 32'h0000_0001 ? array_update_71574 : array_update_71566[1];
  assign array_update_71576[2] = add_71507 == 32'h0000_0002 ? array_update_71574 : array_update_71566[2];
  assign array_update_71576[3] = add_71507 == 32'h0000_0003 ? array_update_71574 : array_update_71566[3];
  assign array_update_71576[4] = add_71507 == 32'h0000_0004 ? array_update_71574 : array_update_71566[4];
  assign array_update_71576[5] = add_71507 == 32'h0000_0005 ? array_update_71574 : array_update_71566[5];
  assign array_update_71576[6] = add_71507 == 32'h0000_0006 ? array_update_71574 : array_update_71566[6];
  assign array_update_71576[7] = add_71507 == 32'h0000_0007 ? array_update_71574 : array_update_71566[7];
  assign array_update_71576[8] = add_71507 == 32'h0000_0008 ? array_update_71574 : array_update_71566[8];
  assign array_update_71576[9] = add_71507 == 32'h0000_0009 ? array_update_71574 : array_update_71566[9];
  assign array_update_71578[0] = add_71509 == 32'h0000_0000 ? array_update_71575 : array_update_71568[0];
  assign array_update_71578[1] = add_71509 == 32'h0000_0001 ? array_update_71575 : array_update_71568[1];
  assign array_update_71578[2] = add_71509 == 32'h0000_0002 ? array_update_71575 : array_update_71568[2];
  assign array_update_71578[3] = add_71509 == 32'h0000_0003 ? array_update_71575 : array_update_71568[3];
  assign array_update_71578[4] = add_71509 == 32'h0000_0004 ? array_update_71575 : array_update_71568[4];
  assign array_update_71578[5] = add_71509 == 32'h0000_0005 ? array_update_71575 : array_update_71568[5];
  assign array_update_71578[6] = add_71509 == 32'h0000_0006 ? array_update_71575 : array_update_71568[6];
  assign array_update_71578[7] = add_71509 == 32'h0000_0007 ? array_update_71575 : array_update_71568[7];
  assign array_update_71578[8] = add_71509 == 32'h0000_0008 ? array_update_71575 : array_update_71568[8];
  assign array_update_71578[9] = add_71509 == 32'h0000_0009 ? array_update_71575 : array_update_71568[9];
  assign array_index_71580 = array_update_71576[add_71507 > 32'h0000_0009 ? 4'h9 : add_71507[3:0]];
  assign add_71581 = add_71571 + 32'h0000_0001;
  assign array_index_71582 = array_update_71578[add_71509 > 32'h0000_0009 ? 4'h9 : add_71509[3:0]];
  assign add_71583 = add_71573 + 32'h0000_0001;
  assign array_update_71584[0] = add_71581 == 32'h0000_0000 ? TestBlock__A_op57 : array_index_71580[0];
  assign array_update_71584[1] = add_71581 == 32'h0000_0001 ? TestBlock__A_op57 : array_index_71580[1];
  assign array_update_71584[2] = add_71581 == 32'h0000_0002 ? TestBlock__A_op57 : array_index_71580[2];
  assign array_update_71584[3] = add_71581 == 32'h0000_0003 ? TestBlock__A_op57 : array_index_71580[3];
  assign array_update_71584[4] = add_71581 == 32'h0000_0004 ? TestBlock__A_op57 : array_index_71580[4];
  assign array_update_71584[5] = add_71581 == 32'h0000_0005 ? TestBlock__A_op57 : array_index_71580[5];
  assign array_update_71584[6] = add_71581 == 32'h0000_0006 ? TestBlock__A_op57 : array_index_71580[6];
  assign array_update_71584[7] = add_71581 == 32'h0000_0007 ? TestBlock__A_op57 : array_index_71580[7];
  assign array_update_71584[8] = add_71581 == 32'h0000_0008 ? TestBlock__A_op57 : array_index_71580[8];
  assign array_update_71584[9] = add_71581 == 32'h0000_0009 ? TestBlock__A_op57 : array_index_71580[9];
  assign array_update_71585[0] = add_71583 == 32'h0000_0000 ? TestBlock__B_op57 : array_index_71582[0];
  assign array_update_71585[1] = add_71583 == 32'h0000_0001 ? TestBlock__B_op57 : array_index_71582[1];
  assign array_update_71585[2] = add_71583 == 32'h0000_0002 ? TestBlock__B_op57 : array_index_71582[2];
  assign array_update_71585[3] = add_71583 == 32'h0000_0003 ? TestBlock__B_op57 : array_index_71582[3];
  assign array_update_71585[4] = add_71583 == 32'h0000_0004 ? TestBlock__B_op57 : array_index_71582[4];
  assign array_update_71585[5] = add_71583 == 32'h0000_0005 ? TestBlock__B_op57 : array_index_71582[5];
  assign array_update_71585[6] = add_71583 == 32'h0000_0006 ? TestBlock__B_op57 : array_index_71582[6];
  assign array_update_71585[7] = add_71583 == 32'h0000_0007 ? TestBlock__B_op57 : array_index_71582[7];
  assign array_update_71585[8] = add_71583 == 32'h0000_0008 ? TestBlock__B_op57 : array_index_71582[8];
  assign array_update_71585[9] = add_71583 == 32'h0000_0009 ? TestBlock__B_op57 : array_index_71582[9];
  assign array_update_71586[0] = add_71507 == 32'h0000_0000 ? array_update_71584 : array_update_71576[0];
  assign array_update_71586[1] = add_71507 == 32'h0000_0001 ? array_update_71584 : array_update_71576[1];
  assign array_update_71586[2] = add_71507 == 32'h0000_0002 ? array_update_71584 : array_update_71576[2];
  assign array_update_71586[3] = add_71507 == 32'h0000_0003 ? array_update_71584 : array_update_71576[3];
  assign array_update_71586[4] = add_71507 == 32'h0000_0004 ? array_update_71584 : array_update_71576[4];
  assign array_update_71586[5] = add_71507 == 32'h0000_0005 ? array_update_71584 : array_update_71576[5];
  assign array_update_71586[6] = add_71507 == 32'h0000_0006 ? array_update_71584 : array_update_71576[6];
  assign array_update_71586[7] = add_71507 == 32'h0000_0007 ? array_update_71584 : array_update_71576[7];
  assign array_update_71586[8] = add_71507 == 32'h0000_0008 ? array_update_71584 : array_update_71576[8];
  assign array_update_71586[9] = add_71507 == 32'h0000_0009 ? array_update_71584 : array_update_71576[9];
  assign array_update_71588[0] = add_71509 == 32'h0000_0000 ? array_update_71585 : array_update_71578[0];
  assign array_update_71588[1] = add_71509 == 32'h0000_0001 ? array_update_71585 : array_update_71578[1];
  assign array_update_71588[2] = add_71509 == 32'h0000_0002 ? array_update_71585 : array_update_71578[2];
  assign array_update_71588[3] = add_71509 == 32'h0000_0003 ? array_update_71585 : array_update_71578[3];
  assign array_update_71588[4] = add_71509 == 32'h0000_0004 ? array_update_71585 : array_update_71578[4];
  assign array_update_71588[5] = add_71509 == 32'h0000_0005 ? array_update_71585 : array_update_71578[5];
  assign array_update_71588[6] = add_71509 == 32'h0000_0006 ? array_update_71585 : array_update_71578[6];
  assign array_update_71588[7] = add_71509 == 32'h0000_0007 ? array_update_71585 : array_update_71578[7];
  assign array_update_71588[8] = add_71509 == 32'h0000_0008 ? array_update_71585 : array_update_71578[8];
  assign array_update_71588[9] = add_71509 == 32'h0000_0009 ? array_update_71585 : array_update_71578[9];
  assign array_index_71590 = array_update_71586[add_71507 > 32'h0000_0009 ? 4'h9 : add_71507[3:0]];
  assign add_71591 = add_71581 + 32'h0000_0001;
  assign array_index_71592 = array_update_71588[add_71509 > 32'h0000_0009 ? 4'h9 : add_71509[3:0]];
  assign add_71593 = add_71583 + 32'h0000_0001;
  assign array_update_71594[0] = add_71591 == 32'h0000_0000 ? TestBlock__A_op58 : array_index_71590[0];
  assign array_update_71594[1] = add_71591 == 32'h0000_0001 ? TestBlock__A_op58 : array_index_71590[1];
  assign array_update_71594[2] = add_71591 == 32'h0000_0002 ? TestBlock__A_op58 : array_index_71590[2];
  assign array_update_71594[3] = add_71591 == 32'h0000_0003 ? TestBlock__A_op58 : array_index_71590[3];
  assign array_update_71594[4] = add_71591 == 32'h0000_0004 ? TestBlock__A_op58 : array_index_71590[4];
  assign array_update_71594[5] = add_71591 == 32'h0000_0005 ? TestBlock__A_op58 : array_index_71590[5];
  assign array_update_71594[6] = add_71591 == 32'h0000_0006 ? TestBlock__A_op58 : array_index_71590[6];
  assign array_update_71594[7] = add_71591 == 32'h0000_0007 ? TestBlock__A_op58 : array_index_71590[7];
  assign array_update_71594[8] = add_71591 == 32'h0000_0008 ? TestBlock__A_op58 : array_index_71590[8];
  assign array_update_71594[9] = add_71591 == 32'h0000_0009 ? TestBlock__A_op58 : array_index_71590[9];
  assign array_update_71595[0] = add_71593 == 32'h0000_0000 ? TestBlock__B_op58 : array_index_71592[0];
  assign array_update_71595[1] = add_71593 == 32'h0000_0001 ? TestBlock__B_op58 : array_index_71592[1];
  assign array_update_71595[2] = add_71593 == 32'h0000_0002 ? TestBlock__B_op58 : array_index_71592[2];
  assign array_update_71595[3] = add_71593 == 32'h0000_0003 ? TestBlock__B_op58 : array_index_71592[3];
  assign array_update_71595[4] = add_71593 == 32'h0000_0004 ? TestBlock__B_op58 : array_index_71592[4];
  assign array_update_71595[5] = add_71593 == 32'h0000_0005 ? TestBlock__B_op58 : array_index_71592[5];
  assign array_update_71595[6] = add_71593 == 32'h0000_0006 ? TestBlock__B_op58 : array_index_71592[6];
  assign array_update_71595[7] = add_71593 == 32'h0000_0007 ? TestBlock__B_op58 : array_index_71592[7];
  assign array_update_71595[8] = add_71593 == 32'h0000_0008 ? TestBlock__B_op58 : array_index_71592[8];
  assign array_update_71595[9] = add_71593 == 32'h0000_0009 ? TestBlock__B_op58 : array_index_71592[9];
  assign array_update_71596[0] = add_71507 == 32'h0000_0000 ? array_update_71594 : array_update_71586[0];
  assign array_update_71596[1] = add_71507 == 32'h0000_0001 ? array_update_71594 : array_update_71586[1];
  assign array_update_71596[2] = add_71507 == 32'h0000_0002 ? array_update_71594 : array_update_71586[2];
  assign array_update_71596[3] = add_71507 == 32'h0000_0003 ? array_update_71594 : array_update_71586[3];
  assign array_update_71596[4] = add_71507 == 32'h0000_0004 ? array_update_71594 : array_update_71586[4];
  assign array_update_71596[5] = add_71507 == 32'h0000_0005 ? array_update_71594 : array_update_71586[5];
  assign array_update_71596[6] = add_71507 == 32'h0000_0006 ? array_update_71594 : array_update_71586[6];
  assign array_update_71596[7] = add_71507 == 32'h0000_0007 ? array_update_71594 : array_update_71586[7];
  assign array_update_71596[8] = add_71507 == 32'h0000_0008 ? array_update_71594 : array_update_71586[8];
  assign array_update_71596[9] = add_71507 == 32'h0000_0009 ? array_update_71594 : array_update_71586[9];
  assign array_update_71598[0] = add_71509 == 32'h0000_0000 ? array_update_71595 : array_update_71588[0];
  assign array_update_71598[1] = add_71509 == 32'h0000_0001 ? array_update_71595 : array_update_71588[1];
  assign array_update_71598[2] = add_71509 == 32'h0000_0002 ? array_update_71595 : array_update_71588[2];
  assign array_update_71598[3] = add_71509 == 32'h0000_0003 ? array_update_71595 : array_update_71588[3];
  assign array_update_71598[4] = add_71509 == 32'h0000_0004 ? array_update_71595 : array_update_71588[4];
  assign array_update_71598[5] = add_71509 == 32'h0000_0005 ? array_update_71595 : array_update_71588[5];
  assign array_update_71598[6] = add_71509 == 32'h0000_0006 ? array_update_71595 : array_update_71588[6];
  assign array_update_71598[7] = add_71509 == 32'h0000_0007 ? array_update_71595 : array_update_71588[7];
  assign array_update_71598[8] = add_71509 == 32'h0000_0008 ? array_update_71595 : array_update_71588[8];
  assign array_update_71598[9] = add_71509 == 32'h0000_0009 ? array_update_71595 : array_update_71588[9];
  assign array_index_71600 = array_update_71596[add_71507 > 32'h0000_0009 ? 4'h9 : add_71507[3:0]];
  assign add_71601 = add_71591 + 32'h0000_0001;
  assign array_index_71602 = array_update_71598[add_71509 > 32'h0000_0009 ? 4'h9 : add_71509[3:0]];
  assign add_71603 = add_71593 + 32'h0000_0001;
  assign array_update_71604[0] = add_71601 == 32'h0000_0000 ? TestBlock__A_op59 : array_index_71600[0];
  assign array_update_71604[1] = add_71601 == 32'h0000_0001 ? TestBlock__A_op59 : array_index_71600[1];
  assign array_update_71604[2] = add_71601 == 32'h0000_0002 ? TestBlock__A_op59 : array_index_71600[2];
  assign array_update_71604[3] = add_71601 == 32'h0000_0003 ? TestBlock__A_op59 : array_index_71600[3];
  assign array_update_71604[4] = add_71601 == 32'h0000_0004 ? TestBlock__A_op59 : array_index_71600[4];
  assign array_update_71604[5] = add_71601 == 32'h0000_0005 ? TestBlock__A_op59 : array_index_71600[5];
  assign array_update_71604[6] = add_71601 == 32'h0000_0006 ? TestBlock__A_op59 : array_index_71600[6];
  assign array_update_71604[7] = add_71601 == 32'h0000_0007 ? TestBlock__A_op59 : array_index_71600[7];
  assign array_update_71604[8] = add_71601 == 32'h0000_0008 ? TestBlock__A_op59 : array_index_71600[8];
  assign array_update_71604[9] = add_71601 == 32'h0000_0009 ? TestBlock__A_op59 : array_index_71600[9];
  assign array_update_71606[0] = add_71603 == 32'h0000_0000 ? TestBlock__B_op59 : array_index_71602[0];
  assign array_update_71606[1] = add_71603 == 32'h0000_0001 ? TestBlock__B_op59 : array_index_71602[1];
  assign array_update_71606[2] = add_71603 == 32'h0000_0002 ? TestBlock__B_op59 : array_index_71602[2];
  assign array_update_71606[3] = add_71603 == 32'h0000_0003 ? TestBlock__B_op59 : array_index_71602[3];
  assign array_update_71606[4] = add_71603 == 32'h0000_0004 ? TestBlock__B_op59 : array_index_71602[4];
  assign array_update_71606[5] = add_71603 == 32'h0000_0005 ? TestBlock__B_op59 : array_index_71602[5];
  assign array_update_71606[6] = add_71603 == 32'h0000_0006 ? TestBlock__B_op59 : array_index_71602[6];
  assign array_update_71606[7] = add_71603 == 32'h0000_0007 ? TestBlock__B_op59 : array_index_71602[7];
  assign array_update_71606[8] = add_71603 == 32'h0000_0008 ? TestBlock__B_op59 : array_index_71602[8];
  assign array_update_71606[9] = add_71603 == 32'h0000_0009 ? TestBlock__B_op59 : array_index_71602[9];
  assign array_update_71608[0] = add_71507 == 32'h0000_0000 ? array_update_71604 : array_update_71596[0];
  assign array_update_71608[1] = add_71507 == 32'h0000_0001 ? array_update_71604 : array_update_71596[1];
  assign array_update_71608[2] = add_71507 == 32'h0000_0002 ? array_update_71604 : array_update_71596[2];
  assign array_update_71608[3] = add_71507 == 32'h0000_0003 ? array_update_71604 : array_update_71596[3];
  assign array_update_71608[4] = add_71507 == 32'h0000_0004 ? array_update_71604 : array_update_71596[4];
  assign array_update_71608[5] = add_71507 == 32'h0000_0005 ? array_update_71604 : array_update_71596[5];
  assign array_update_71608[6] = add_71507 == 32'h0000_0006 ? array_update_71604 : array_update_71596[6];
  assign array_update_71608[7] = add_71507 == 32'h0000_0007 ? array_update_71604 : array_update_71596[7];
  assign array_update_71608[8] = add_71507 == 32'h0000_0008 ? array_update_71604 : array_update_71596[8];
  assign array_update_71608[9] = add_71507 == 32'h0000_0009 ? array_update_71604 : array_update_71596[9];
  assign add_71609 = add_71507 + 32'h0000_0001;
  assign array_update_71610[0] = add_71509 == 32'h0000_0000 ? array_update_71606 : array_update_71598[0];
  assign array_update_71610[1] = add_71509 == 32'h0000_0001 ? array_update_71606 : array_update_71598[1];
  assign array_update_71610[2] = add_71509 == 32'h0000_0002 ? array_update_71606 : array_update_71598[2];
  assign array_update_71610[3] = add_71509 == 32'h0000_0003 ? array_update_71606 : array_update_71598[3];
  assign array_update_71610[4] = add_71509 == 32'h0000_0004 ? array_update_71606 : array_update_71598[4];
  assign array_update_71610[5] = add_71509 == 32'h0000_0005 ? array_update_71606 : array_update_71598[5];
  assign array_update_71610[6] = add_71509 == 32'h0000_0006 ? array_update_71606 : array_update_71598[6];
  assign array_update_71610[7] = add_71509 == 32'h0000_0007 ? array_update_71606 : array_update_71598[7];
  assign array_update_71610[8] = add_71509 == 32'h0000_0008 ? array_update_71606 : array_update_71598[8];
  assign array_update_71610[9] = add_71509 == 32'h0000_0009 ? array_update_71606 : array_update_71598[9];
  assign add_71611 = add_71509 + 32'h0000_0001;
  assign array_index_71612 = array_update_71608[add_71609 > 32'h0000_0009 ? 4'h9 : add_71609[3:0]];
  assign literal_71613 = 32'h0000_0000;
  assign array_index_71614 = array_update_71610[add_71611 > 32'h0000_0009 ? 4'h9 : add_71611[3:0]];
  assign literal_71615 = 32'h0000_0000;
  assign array_update_71616[0] = literal_71613 == 32'h0000_0000 ? TestBlock__A_op60 : array_index_71612[0];
  assign array_update_71616[1] = literal_71613 == 32'h0000_0001 ? TestBlock__A_op60 : array_index_71612[1];
  assign array_update_71616[2] = literal_71613 == 32'h0000_0002 ? TestBlock__A_op60 : array_index_71612[2];
  assign array_update_71616[3] = literal_71613 == 32'h0000_0003 ? TestBlock__A_op60 : array_index_71612[3];
  assign array_update_71616[4] = literal_71613 == 32'h0000_0004 ? TestBlock__A_op60 : array_index_71612[4];
  assign array_update_71616[5] = literal_71613 == 32'h0000_0005 ? TestBlock__A_op60 : array_index_71612[5];
  assign array_update_71616[6] = literal_71613 == 32'h0000_0006 ? TestBlock__A_op60 : array_index_71612[6];
  assign array_update_71616[7] = literal_71613 == 32'h0000_0007 ? TestBlock__A_op60 : array_index_71612[7];
  assign array_update_71616[8] = literal_71613 == 32'h0000_0008 ? TestBlock__A_op60 : array_index_71612[8];
  assign array_update_71616[9] = literal_71613 == 32'h0000_0009 ? TestBlock__A_op60 : array_index_71612[9];
  assign array_update_71617[0] = literal_71615 == 32'h0000_0000 ? TestBlock__B_op60 : array_index_71614[0];
  assign array_update_71617[1] = literal_71615 == 32'h0000_0001 ? TestBlock__B_op60 : array_index_71614[1];
  assign array_update_71617[2] = literal_71615 == 32'h0000_0002 ? TestBlock__B_op60 : array_index_71614[2];
  assign array_update_71617[3] = literal_71615 == 32'h0000_0003 ? TestBlock__B_op60 : array_index_71614[3];
  assign array_update_71617[4] = literal_71615 == 32'h0000_0004 ? TestBlock__B_op60 : array_index_71614[4];
  assign array_update_71617[5] = literal_71615 == 32'h0000_0005 ? TestBlock__B_op60 : array_index_71614[5];
  assign array_update_71617[6] = literal_71615 == 32'h0000_0006 ? TestBlock__B_op60 : array_index_71614[6];
  assign array_update_71617[7] = literal_71615 == 32'h0000_0007 ? TestBlock__B_op60 : array_index_71614[7];
  assign array_update_71617[8] = literal_71615 == 32'h0000_0008 ? TestBlock__B_op60 : array_index_71614[8];
  assign array_update_71617[9] = literal_71615 == 32'h0000_0009 ? TestBlock__B_op60 : array_index_71614[9];
  assign array_update_71618[0] = add_71609 == 32'h0000_0000 ? array_update_71616 : array_update_71608[0];
  assign array_update_71618[1] = add_71609 == 32'h0000_0001 ? array_update_71616 : array_update_71608[1];
  assign array_update_71618[2] = add_71609 == 32'h0000_0002 ? array_update_71616 : array_update_71608[2];
  assign array_update_71618[3] = add_71609 == 32'h0000_0003 ? array_update_71616 : array_update_71608[3];
  assign array_update_71618[4] = add_71609 == 32'h0000_0004 ? array_update_71616 : array_update_71608[4];
  assign array_update_71618[5] = add_71609 == 32'h0000_0005 ? array_update_71616 : array_update_71608[5];
  assign array_update_71618[6] = add_71609 == 32'h0000_0006 ? array_update_71616 : array_update_71608[6];
  assign array_update_71618[7] = add_71609 == 32'h0000_0007 ? array_update_71616 : array_update_71608[7];
  assign array_update_71618[8] = add_71609 == 32'h0000_0008 ? array_update_71616 : array_update_71608[8];
  assign array_update_71618[9] = add_71609 == 32'h0000_0009 ? array_update_71616 : array_update_71608[9];
  assign array_update_71620[0] = add_71611 == 32'h0000_0000 ? array_update_71617 : array_update_71610[0];
  assign array_update_71620[1] = add_71611 == 32'h0000_0001 ? array_update_71617 : array_update_71610[1];
  assign array_update_71620[2] = add_71611 == 32'h0000_0002 ? array_update_71617 : array_update_71610[2];
  assign array_update_71620[3] = add_71611 == 32'h0000_0003 ? array_update_71617 : array_update_71610[3];
  assign array_update_71620[4] = add_71611 == 32'h0000_0004 ? array_update_71617 : array_update_71610[4];
  assign array_update_71620[5] = add_71611 == 32'h0000_0005 ? array_update_71617 : array_update_71610[5];
  assign array_update_71620[6] = add_71611 == 32'h0000_0006 ? array_update_71617 : array_update_71610[6];
  assign array_update_71620[7] = add_71611 == 32'h0000_0007 ? array_update_71617 : array_update_71610[7];
  assign array_update_71620[8] = add_71611 == 32'h0000_0008 ? array_update_71617 : array_update_71610[8];
  assign array_update_71620[9] = add_71611 == 32'h0000_0009 ? array_update_71617 : array_update_71610[9];
  assign array_index_71622 = array_update_71618[add_71609 > 32'h0000_0009 ? 4'h9 : add_71609[3:0]];
  assign add_71623 = literal_71613 + 32'h0000_0001;
  assign array_index_71624 = array_update_71620[add_71611 > 32'h0000_0009 ? 4'h9 : add_71611[3:0]];
  assign add_71625 = literal_71615 + 32'h0000_0001;
  assign array_update_71626[0] = add_71623 == 32'h0000_0000 ? TestBlock__A_op61 : array_index_71622[0];
  assign array_update_71626[1] = add_71623 == 32'h0000_0001 ? TestBlock__A_op61 : array_index_71622[1];
  assign array_update_71626[2] = add_71623 == 32'h0000_0002 ? TestBlock__A_op61 : array_index_71622[2];
  assign array_update_71626[3] = add_71623 == 32'h0000_0003 ? TestBlock__A_op61 : array_index_71622[3];
  assign array_update_71626[4] = add_71623 == 32'h0000_0004 ? TestBlock__A_op61 : array_index_71622[4];
  assign array_update_71626[5] = add_71623 == 32'h0000_0005 ? TestBlock__A_op61 : array_index_71622[5];
  assign array_update_71626[6] = add_71623 == 32'h0000_0006 ? TestBlock__A_op61 : array_index_71622[6];
  assign array_update_71626[7] = add_71623 == 32'h0000_0007 ? TestBlock__A_op61 : array_index_71622[7];
  assign array_update_71626[8] = add_71623 == 32'h0000_0008 ? TestBlock__A_op61 : array_index_71622[8];
  assign array_update_71626[9] = add_71623 == 32'h0000_0009 ? TestBlock__A_op61 : array_index_71622[9];
  assign array_update_71627[0] = add_71625 == 32'h0000_0000 ? TestBlock__B_op61 : array_index_71624[0];
  assign array_update_71627[1] = add_71625 == 32'h0000_0001 ? TestBlock__B_op61 : array_index_71624[1];
  assign array_update_71627[2] = add_71625 == 32'h0000_0002 ? TestBlock__B_op61 : array_index_71624[2];
  assign array_update_71627[3] = add_71625 == 32'h0000_0003 ? TestBlock__B_op61 : array_index_71624[3];
  assign array_update_71627[4] = add_71625 == 32'h0000_0004 ? TestBlock__B_op61 : array_index_71624[4];
  assign array_update_71627[5] = add_71625 == 32'h0000_0005 ? TestBlock__B_op61 : array_index_71624[5];
  assign array_update_71627[6] = add_71625 == 32'h0000_0006 ? TestBlock__B_op61 : array_index_71624[6];
  assign array_update_71627[7] = add_71625 == 32'h0000_0007 ? TestBlock__B_op61 : array_index_71624[7];
  assign array_update_71627[8] = add_71625 == 32'h0000_0008 ? TestBlock__B_op61 : array_index_71624[8];
  assign array_update_71627[9] = add_71625 == 32'h0000_0009 ? TestBlock__B_op61 : array_index_71624[9];
  assign array_update_71628[0] = add_71609 == 32'h0000_0000 ? array_update_71626 : array_update_71618[0];
  assign array_update_71628[1] = add_71609 == 32'h0000_0001 ? array_update_71626 : array_update_71618[1];
  assign array_update_71628[2] = add_71609 == 32'h0000_0002 ? array_update_71626 : array_update_71618[2];
  assign array_update_71628[3] = add_71609 == 32'h0000_0003 ? array_update_71626 : array_update_71618[3];
  assign array_update_71628[4] = add_71609 == 32'h0000_0004 ? array_update_71626 : array_update_71618[4];
  assign array_update_71628[5] = add_71609 == 32'h0000_0005 ? array_update_71626 : array_update_71618[5];
  assign array_update_71628[6] = add_71609 == 32'h0000_0006 ? array_update_71626 : array_update_71618[6];
  assign array_update_71628[7] = add_71609 == 32'h0000_0007 ? array_update_71626 : array_update_71618[7];
  assign array_update_71628[8] = add_71609 == 32'h0000_0008 ? array_update_71626 : array_update_71618[8];
  assign array_update_71628[9] = add_71609 == 32'h0000_0009 ? array_update_71626 : array_update_71618[9];
  assign array_update_71630[0] = add_71611 == 32'h0000_0000 ? array_update_71627 : array_update_71620[0];
  assign array_update_71630[1] = add_71611 == 32'h0000_0001 ? array_update_71627 : array_update_71620[1];
  assign array_update_71630[2] = add_71611 == 32'h0000_0002 ? array_update_71627 : array_update_71620[2];
  assign array_update_71630[3] = add_71611 == 32'h0000_0003 ? array_update_71627 : array_update_71620[3];
  assign array_update_71630[4] = add_71611 == 32'h0000_0004 ? array_update_71627 : array_update_71620[4];
  assign array_update_71630[5] = add_71611 == 32'h0000_0005 ? array_update_71627 : array_update_71620[5];
  assign array_update_71630[6] = add_71611 == 32'h0000_0006 ? array_update_71627 : array_update_71620[6];
  assign array_update_71630[7] = add_71611 == 32'h0000_0007 ? array_update_71627 : array_update_71620[7];
  assign array_update_71630[8] = add_71611 == 32'h0000_0008 ? array_update_71627 : array_update_71620[8];
  assign array_update_71630[9] = add_71611 == 32'h0000_0009 ? array_update_71627 : array_update_71620[9];
  assign array_index_71632 = array_update_71628[add_71609 > 32'h0000_0009 ? 4'h9 : add_71609[3:0]];
  assign add_71633 = add_71623 + 32'h0000_0001;
  assign array_index_71634 = array_update_71630[add_71611 > 32'h0000_0009 ? 4'h9 : add_71611[3:0]];
  assign add_71635 = add_71625 + 32'h0000_0001;
  assign array_update_71636[0] = add_71633 == 32'h0000_0000 ? TestBlock__A_op62 : array_index_71632[0];
  assign array_update_71636[1] = add_71633 == 32'h0000_0001 ? TestBlock__A_op62 : array_index_71632[1];
  assign array_update_71636[2] = add_71633 == 32'h0000_0002 ? TestBlock__A_op62 : array_index_71632[2];
  assign array_update_71636[3] = add_71633 == 32'h0000_0003 ? TestBlock__A_op62 : array_index_71632[3];
  assign array_update_71636[4] = add_71633 == 32'h0000_0004 ? TestBlock__A_op62 : array_index_71632[4];
  assign array_update_71636[5] = add_71633 == 32'h0000_0005 ? TestBlock__A_op62 : array_index_71632[5];
  assign array_update_71636[6] = add_71633 == 32'h0000_0006 ? TestBlock__A_op62 : array_index_71632[6];
  assign array_update_71636[7] = add_71633 == 32'h0000_0007 ? TestBlock__A_op62 : array_index_71632[7];
  assign array_update_71636[8] = add_71633 == 32'h0000_0008 ? TestBlock__A_op62 : array_index_71632[8];
  assign array_update_71636[9] = add_71633 == 32'h0000_0009 ? TestBlock__A_op62 : array_index_71632[9];
  assign array_update_71637[0] = add_71635 == 32'h0000_0000 ? TestBlock__B_op62 : array_index_71634[0];
  assign array_update_71637[1] = add_71635 == 32'h0000_0001 ? TestBlock__B_op62 : array_index_71634[1];
  assign array_update_71637[2] = add_71635 == 32'h0000_0002 ? TestBlock__B_op62 : array_index_71634[2];
  assign array_update_71637[3] = add_71635 == 32'h0000_0003 ? TestBlock__B_op62 : array_index_71634[3];
  assign array_update_71637[4] = add_71635 == 32'h0000_0004 ? TestBlock__B_op62 : array_index_71634[4];
  assign array_update_71637[5] = add_71635 == 32'h0000_0005 ? TestBlock__B_op62 : array_index_71634[5];
  assign array_update_71637[6] = add_71635 == 32'h0000_0006 ? TestBlock__B_op62 : array_index_71634[6];
  assign array_update_71637[7] = add_71635 == 32'h0000_0007 ? TestBlock__B_op62 : array_index_71634[7];
  assign array_update_71637[8] = add_71635 == 32'h0000_0008 ? TestBlock__B_op62 : array_index_71634[8];
  assign array_update_71637[9] = add_71635 == 32'h0000_0009 ? TestBlock__B_op62 : array_index_71634[9];
  assign array_update_71638[0] = add_71609 == 32'h0000_0000 ? array_update_71636 : array_update_71628[0];
  assign array_update_71638[1] = add_71609 == 32'h0000_0001 ? array_update_71636 : array_update_71628[1];
  assign array_update_71638[2] = add_71609 == 32'h0000_0002 ? array_update_71636 : array_update_71628[2];
  assign array_update_71638[3] = add_71609 == 32'h0000_0003 ? array_update_71636 : array_update_71628[3];
  assign array_update_71638[4] = add_71609 == 32'h0000_0004 ? array_update_71636 : array_update_71628[4];
  assign array_update_71638[5] = add_71609 == 32'h0000_0005 ? array_update_71636 : array_update_71628[5];
  assign array_update_71638[6] = add_71609 == 32'h0000_0006 ? array_update_71636 : array_update_71628[6];
  assign array_update_71638[7] = add_71609 == 32'h0000_0007 ? array_update_71636 : array_update_71628[7];
  assign array_update_71638[8] = add_71609 == 32'h0000_0008 ? array_update_71636 : array_update_71628[8];
  assign array_update_71638[9] = add_71609 == 32'h0000_0009 ? array_update_71636 : array_update_71628[9];
  assign array_update_71640[0] = add_71611 == 32'h0000_0000 ? array_update_71637 : array_update_71630[0];
  assign array_update_71640[1] = add_71611 == 32'h0000_0001 ? array_update_71637 : array_update_71630[1];
  assign array_update_71640[2] = add_71611 == 32'h0000_0002 ? array_update_71637 : array_update_71630[2];
  assign array_update_71640[3] = add_71611 == 32'h0000_0003 ? array_update_71637 : array_update_71630[3];
  assign array_update_71640[4] = add_71611 == 32'h0000_0004 ? array_update_71637 : array_update_71630[4];
  assign array_update_71640[5] = add_71611 == 32'h0000_0005 ? array_update_71637 : array_update_71630[5];
  assign array_update_71640[6] = add_71611 == 32'h0000_0006 ? array_update_71637 : array_update_71630[6];
  assign array_update_71640[7] = add_71611 == 32'h0000_0007 ? array_update_71637 : array_update_71630[7];
  assign array_update_71640[8] = add_71611 == 32'h0000_0008 ? array_update_71637 : array_update_71630[8];
  assign array_update_71640[9] = add_71611 == 32'h0000_0009 ? array_update_71637 : array_update_71630[9];
  assign array_index_71642 = array_update_71638[add_71609 > 32'h0000_0009 ? 4'h9 : add_71609[3:0]];
  assign add_71643 = add_71633 + 32'h0000_0001;
  assign array_index_71644 = array_update_71640[add_71611 > 32'h0000_0009 ? 4'h9 : add_71611[3:0]];
  assign add_71645 = add_71635 + 32'h0000_0001;
  assign array_update_71646[0] = add_71643 == 32'h0000_0000 ? TestBlock__A_op63 : array_index_71642[0];
  assign array_update_71646[1] = add_71643 == 32'h0000_0001 ? TestBlock__A_op63 : array_index_71642[1];
  assign array_update_71646[2] = add_71643 == 32'h0000_0002 ? TestBlock__A_op63 : array_index_71642[2];
  assign array_update_71646[3] = add_71643 == 32'h0000_0003 ? TestBlock__A_op63 : array_index_71642[3];
  assign array_update_71646[4] = add_71643 == 32'h0000_0004 ? TestBlock__A_op63 : array_index_71642[4];
  assign array_update_71646[5] = add_71643 == 32'h0000_0005 ? TestBlock__A_op63 : array_index_71642[5];
  assign array_update_71646[6] = add_71643 == 32'h0000_0006 ? TestBlock__A_op63 : array_index_71642[6];
  assign array_update_71646[7] = add_71643 == 32'h0000_0007 ? TestBlock__A_op63 : array_index_71642[7];
  assign array_update_71646[8] = add_71643 == 32'h0000_0008 ? TestBlock__A_op63 : array_index_71642[8];
  assign array_update_71646[9] = add_71643 == 32'h0000_0009 ? TestBlock__A_op63 : array_index_71642[9];
  assign array_update_71647[0] = add_71645 == 32'h0000_0000 ? TestBlock__B_op63 : array_index_71644[0];
  assign array_update_71647[1] = add_71645 == 32'h0000_0001 ? TestBlock__B_op63 : array_index_71644[1];
  assign array_update_71647[2] = add_71645 == 32'h0000_0002 ? TestBlock__B_op63 : array_index_71644[2];
  assign array_update_71647[3] = add_71645 == 32'h0000_0003 ? TestBlock__B_op63 : array_index_71644[3];
  assign array_update_71647[4] = add_71645 == 32'h0000_0004 ? TestBlock__B_op63 : array_index_71644[4];
  assign array_update_71647[5] = add_71645 == 32'h0000_0005 ? TestBlock__B_op63 : array_index_71644[5];
  assign array_update_71647[6] = add_71645 == 32'h0000_0006 ? TestBlock__B_op63 : array_index_71644[6];
  assign array_update_71647[7] = add_71645 == 32'h0000_0007 ? TestBlock__B_op63 : array_index_71644[7];
  assign array_update_71647[8] = add_71645 == 32'h0000_0008 ? TestBlock__B_op63 : array_index_71644[8];
  assign array_update_71647[9] = add_71645 == 32'h0000_0009 ? TestBlock__B_op63 : array_index_71644[9];
  assign array_update_71648[0] = add_71609 == 32'h0000_0000 ? array_update_71646 : array_update_71638[0];
  assign array_update_71648[1] = add_71609 == 32'h0000_0001 ? array_update_71646 : array_update_71638[1];
  assign array_update_71648[2] = add_71609 == 32'h0000_0002 ? array_update_71646 : array_update_71638[2];
  assign array_update_71648[3] = add_71609 == 32'h0000_0003 ? array_update_71646 : array_update_71638[3];
  assign array_update_71648[4] = add_71609 == 32'h0000_0004 ? array_update_71646 : array_update_71638[4];
  assign array_update_71648[5] = add_71609 == 32'h0000_0005 ? array_update_71646 : array_update_71638[5];
  assign array_update_71648[6] = add_71609 == 32'h0000_0006 ? array_update_71646 : array_update_71638[6];
  assign array_update_71648[7] = add_71609 == 32'h0000_0007 ? array_update_71646 : array_update_71638[7];
  assign array_update_71648[8] = add_71609 == 32'h0000_0008 ? array_update_71646 : array_update_71638[8];
  assign array_update_71648[9] = add_71609 == 32'h0000_0009 ? array_update_71646 : array_update_71638[9];
  assign array_update_71650[0] = add_71611 == 32'h0000_0000 ? array_update_71647 : array_update_71640[0];
  assign array_update_71650[1] = add_71611 == 32'h0000_0001 ? array_update_71647 : array_update_71640[1];
  assign array_update_71650[2] = add_71611 == 32'h0000_0002 ? array_update_71647 : array_update_71640[2];
  assign array_update_71650[3] = add_71611 == 32'h0000_0003 ? array_update_71647 : array_update_71640[3];
  assign array_update_71650[4] = add_71611 == 32'h0000_0004 ? array_update_71647 : array_update_71640[4];
  assign array_update_71650[5] = add_71611 == 32'h0000_0005 ? array_update_71647 : array_update_71640[5];
  assign array_update_71650[6] = add_71611 == 32'h0000_0006 ? array_update_71647 : array_update_71640[6];
  assign array_update_71650[7] = add_71611 == 32'h0000_0007 ? array_update_71647 : array_update_71640[7];
  assign array_update_71650[8] = add_71611 == 32'h0000_0008 ? array_update_71647 : array_update_71640[8];
  assign array_update_71650[9] = add_71611 == 32'h0000_0009 ? array_update_71647 : array_update_71640[9];
  assign array_index_71652 = array_update_71648[add_71609 > 32'h0000_0009 ? 4'h9 : add_71609[3:0]];
  assign add_71653 = add_71643 + 32'h0000_0001;
  assign array_index_71654 = array_update_71650[add_71611 > 32'h0000_0009 ? 4'h9 : add_71611[3:0]];
  assign add_71655 = add_71645 + 32'h0000_0001;
  assign array_update_71656[0] = add_71653 == 32'h0000_0000 ? TestBlock__A_op64 : array_index_71652[0];
  assign array_update_71656[1] = add_71653 == 32'h0000_0001 ? TestBlock__A_op64 : array_index_71652[1];
  assign array_update_71656[2] = add_71653 == 32'h0000_0002 ? TestBlock__A_op64 : array_index_71652[2];
  assign array_update_71656[3] = add_71653 == 32'h0000_0003 ? TestBlock__A_op64 : array_index_71652[3];
  assign array_update_71656[4] = add_71653 == 32'h0000_0004 ? TestBlock__A_op64 : array_index_71652[4];
  assign array_update_71656[5] = add_71653 == 32'h0000_0005 ? TestBlock__A_op64 : array_index_71652[5];
  assign array_update_71656[6] = add_71653 == 32'h0000_0006 ? TestBlock__A_op64 : array_index_71652[6];
  assign array_update_71656[7] = add_71653 == 32'h0000_0007 ? TestBlock__A_op64 : array_index_71652[7];
  assign array_update_71656[8] = add_71653 == 32'h0000_0008 ? TestBlock__A_op64 : array_index_71652[8];
  assign array_update_71656[9] = add_71653 == 32'h0000_0009 ? TestBlock__A_op64 : array_index_71652[9];
  assign array_update_71657[0] = add_71655 == 32'h0000_0000 ? TestBlock__B_op64 : array_index_71654[0];
  assign array_update_71657[1] = add_71655 == 32'h0000_0001 ? TestBlock__B_op64 : array_index_71654[1];
  assign array_update_71657[2] = add_71655 == 32'h0000_0002 ? TestBlock__B_op64 : array_index_71654[2];
  assign array_update_71657[3] = add_71655 == 32'h0000_0003 ? TestBlock__B_op64 : array_index_71654[3];
  assign array_update_71657[4] = add_71655 == 32'h0000_0004 ? TestBlock__B_op64 : array_index_71654[4];
  assign array_update_71657[5] = add_71655 == 32'h0000_0005 ? TestBlock__B_op64 : array_index_71654[5];
  assign array_update_71657[6] = add_71655 == 32'h0000_0006 ? TestBlock__B_op64 : array_index_71654[6];
  assign array_update_71657[7] = add_71655 == 32'h0000_0007 ? TestBlock__B_op64 : array_index_71654[7];
  assign array_update_71657[8] = add_71655 == 32'h0000_0008 ? TestBlock__B_op64 : array_index_71654[8];
  assign array_update_71657[9] = add_71655 == 32'h0000_0009 ? TestBlock__B_op64 : array_index_71654[9];
  assign array_update_71658[0] = add_71609 == 32'h0000_0000 ? array_update_71656 : array_update_71648[0];
  assign array_update_71658[1] = add_71609 == 32'h0000_0001 ? array_update_71656 : array_update_71648[1];
  assign array_update_71658[2] = add_71609 == 32'h0000_0002 ? array_update_71656 : array_update_71648[2];
  assign array_update_71658[3] = add_71609 == 32'h0000_0003 ? array_update_71656 : array_update_71648[3];
  assign array_update_71658[4] = add_71609 == 32'h0000_0004 ? array_update_71656 : array_update_71648[4];
  assign array_update_71658[5] = add_71609 == 32'h0000_0005 ? array_update_71656 : array_update_71648[5];
  assign array_update_71658[6] = add_71609 == 32'h0000_0006 ? array_update_71656 : array_update_71648[6];
  assign array_update_71658[7] = add_71609 == 32'h0000_0007 ? array_update_71656 : array_update_71648[7];
  assign array_update_71658[8] = add_71609 == 32'h0000_0008 ? array_update_71656 : array_update_71648[8];
  assign array_update_71658[9] = add_71609 == 32'h0000_0009 ? array_update_71656 : array_update_71648[9];
  assign array_update_71660[0] = add_71611 == 32'h0000_0000 ? array_update_71657 : array_update_71650[0];
  assign array_update_71660[1] = add_71611 == 32'h0000_0001 ? array_update_71657 : array_update_71650[1];
  assign array_update_71660[2] = add_71611 == 32'h0000_0002 ? array_update_71657 : array_update_71650[2];
  assign array_update_71660[3] = add_71611 == 32'h0000_0003 ? array_update_71657 : array_update_71650[3];
  assign array_update_71660[4] = add_71611 == 32'h0000_0004 ? array_update_71657 : array_update_71650[4];
  assign array_update_71660[5] = add_71611 == 32'h0000_0005 ? array_update_71657 : array_update_71650[5];
  assign array_update_71660[6] = add_71611 == 32'h0000_0006 ? array_update_71657 : array_update_71650[6];
  assign array_update_71660[7] = add_71611 == 32'h0000_0007 ? array_update_71657 : array_update_71650[7];
  assign array_update_71660[8] = add_71611 == 32'h0000_0008 ? array_update_71657 : array_update_71650[8];
  assign array_update_71660[9] = add_71611 == 32'h0000_0009 ? array_update_71657 : array_update_71650[9];
  assign array_index_71662 = array_update_71658[add_71609 > 32'h0000_0009 ? 4'h9 : add_71609[3:0]];
  assign add_71663 = add_71653 + 32'h0000_0001;
  assign array_index_71664 = array_update_71660[add_71611 > 32'h0000_0009 ? 4'h9 : add_71611[3:0]];
  assign add_71665 = add_71655 + 32'h0000_0001;
  assign array_update_71666[0] = add_71663 == 32'h0000_0000 ? TestBlock__A_op65 : array_index_71662[0];
  assign array_update_71666[1] = add_71663 == 32'h0000_0001 ? TestBlock__A_op65 : array_index_71662[1];
  assign array_update_71666[2] = add_71663 == 32'h0000_0002 ? TestBlock__A_op65 : array_index_71662[2];
  assign array_update_71666[3] = add_71663 == 32'h0000_0003 ? TestBlock__A_op65 : array_index_71662[3];
  assign array_update_71666[4] = add_71663 == 32'h0000_0004 ? TestBlock__A_op65 : array_index_71662[4];
  assign array_update_71666[5] = add_71663 == 32'h0000_0005 ? TestBlock__A_op65 : array_index_71662[5];
  assign array_update_71666[6] = add_71663 == 32'h0000_0006 ? TestBlock__A_op65 : array_index_71662[6];
  assign array_update_71666[7] = add_71663 == 32'h0000_0007 ? TestBlock__A_op65 : array_index_71662[7];
  assign array_update_71666[8] = add_71663 == 32'h0000_0008 ? TestBlock__A_op65 : array_index_71662[8];
  assign array_update_71666[9] = add_71663 == 32'h0000_0009 ? TestBlock__A_op65 : array_index_71662[9];
  assign array_update_71667[0] = add_71665 == 32'h0000_0000 ? TestBlock__B_op65 : array_index_71664[0];
  assign array_update_71667[1] = add_71665 == 32'h0000_0001 ? TestBlock__B_op65 : array_index_71664[1];
  assign array_update_71667[2] = add_71665 == 32'h0000_0002 ? TestBlock__B_op65 : array_index_71664[2];
  assign array_update_71667[3] = add_71665 == 32'h0000_0003 ? TestBlock__B_op65 : array_index_71664[3];
  assign array_update_71667[4] = add_71665 == 32'h0000_0004 ? TestBlock__B_op65 : array_index_71664[4];
  assign array_update_71667[5] = add_71665 == 32'h0000_0005 ? TestBlock__B_op65 : array_index_71664[5];
  assign array_update_71667[6] = add_71665 == 32'h0000_0006 ? TestBlock__B_op65 : array_index_71664[6];
  assign array_update_71667[7] = add_71665 == 32'h0000_0007 ? TestBlock__B_op65 : array_index_71664[7];
  assign array_update_71667[8] = add_71665 == 32'h0000_0008 ? TestBlock__B_op65 : array_index_71664[8];
  assign array_update_71667[9] = add_71665 == 32'h0000_0009 ? TestBlock__B_op65 : array_index_71664[9];
  assign array_update_71668[0] = add_71609 == 32'h0000_0000 ? array_update_71666 : array_update_71658[0];
  assign array_update_71668[1] = add_71609 == 32'h0000_0001 ? array_update_71666 : array_update_71658[1];
  assign array_update_71668[2] = add_71609 == 32'h0000_0002 ? array_update_71666 : array_update_71658[2];
  assign array_update_71668[3] = add_71609 == 32'h0000_0003 ? array_update_71666 : array_update_71658[3];
  assign array_update_71668[4] = add_71609 == 32'h0000_0004 ? array_update_71666 : array_update_71658[4];
  assign array_update_71668[5] = add_71609 == 32'h0000_0005 ? array_update_71666 : array_update_71658[5];
  assign array_update_71668[6] = add_71609 == 32'h0000_0006 ? array_update_71666 : array_update_71658[6];
  assign array_update_71668[7] = add_71609 == 32'h0000_0007 ? array_update_71666 : array_update_71658[7];
  assign array_update_71668[8] = add_71609 == 32'h0000_0008 ? array_update_71666 : array_update_71658[8];
  assign array_update_71668[9] = add_71609 == 32'h0000_0009 ? array_update_71666 : array_update_71658[9];
  assign array_update_71670[0] = add_71611 == 32'h0000_0000 ? array_update_71667 : array_update_71660[0];
  assign array_update_71670[1] = add_71611 == 32'h0000_0001 ? array_update_71667 : array_update_71660[1];
  assign array_update_71670[2] = add_71611 == 32'h0000_0002 ? array_update_71667 : array_update_71660[2];
  assign array_update_71670[3] = add_71611 == 32'h0000_0003 ? array_update_71667 : array_update_71660[3];
  assign array_update_71670[4] = add_71611 == 32'h0000_0004 ? array_update_71667 : array_update_71660[4];
  assign array_update_71670[5] = add_71611 == 32'h0000_0005 ? array_update_71667 : array_update_71660[5];
  assign array_update_71670[6] = add_71611 == 32'h0000_0006 ? array_update_71667 : array_update_71660[6];
  assign array_update_71670[7] = add_71611 == 32'h0000_0007 ? array_update_71667 : array_update_71660[7];
  assign array_update_71670[8] = add_71611 == 32'h0000_0008 ? array_update_71667 : array_update_71660[8];
  assign array_update_71670[9] = add_71611 == 32'h0000_0009 ? array_update_71667 : array_update_71660[9];
  assign array_index_71672 = array_update_71668[add_71609 > 32'h0000_0009 ? 4'h9 : add_71609[3:0]];
  assign add_71673 = add_71663 + 32'h0000_0001;
  assign array_index_71674 = array_update_71670[add_71611 > 32'h0000_0009 ? 4'h9 : add_71611[3:0]];
  assign add_71675 = add_71665 + 32'h0000_0001;
  assign array_update_71676[0] = add_71673 == 32'h0000_0000 ? TestBlock__A_op66 : array_index_71672[0];
  assign array_update_71676[1] = add_71673 == 32'h0000_0001 ? TestBlock__A_op66 : array_index_71672[1];
  assign array_update_71676[2] = add_71673 == 32'h0000_0002 ? TestBlock__A_op66 : array_index_71672[2];
  assign array_update_71676[3] = add_71673 == 32'h0000_0003 ? TestBlock__A_op66 : array_index_71672[3];
  assign array_update_71676[4] = add_71673 == 32'h0000_0004 ? TestBlock__A_op66 : array_index_71672[4];
  assign array_update_71676[5] = add_71673 == 32'h0000_0005 ? TestBlock__A_op66 : array_index_71672[5];
  assign array_update_71676[6] = add_71673 == 32'h0000_0006 ? TestBlock__A_op66 : array_index_71672[6];
  assign array_update_71676[7] = add_71673 == 32'h0000_0007 ? TestBlock__A_op66 : array_index_71672[7];
  assign array_update_71676[8] = add_71673 == 32'h0000_0008 ? TestBlock__A_op66 : array_index_71672[8];
  assign array_update_71676[9] = add_71673 == 32'h0000_0009 ? TestBlock__A_op66 : array_index_71672[9];
  assign array_update_71677[0] = add_71675 == 32'h0000_0000 ? TestBlock__B_op66 : array_index_71674[0];
  assign array_update_71677[1] = add_71675 == 32'h0000_0001 ? TestBlock__B_op66 : array_index_71674[1];
  assign array_update_71677[2] = add_71675 == 32'h0000_0002 ? TestBlock__B_op66 : array_index_71674[2];
  assign array_update_71677[3] = add_71675 == 32'h0000_0003 ? TestBlock__B_op66 : array_index_71674[3];
  assign array_update_71677[4] = add_71675 == 32'h0000_0004 ? TestBlock__B_op66 : array_index_71674[4];
  assign array_update_71677[5] = add_71675 == 32'h0000_0005 ? TestBlock__B_op66 : array_index_71674[5];
  assign array_update_71677[6] = add_71675 == 32'h0000_0006 ? TestBlock__B_op66 : array_index_71674[6];
  assign array_update_71677[7] = add_71675 == 32'h0000_0007 ? TestBlock__B_op66 : array_index_71674[7];
  assign array_update_71677[8] = add_71675 == 32'h0000_0008 ? TestBlock__B_op66 : array_index_71674[8];
  assign array_update_71677[9] = add_71675 == 32'h0000_0009 ? TestBlock__B_op66 : array_index_71674[9];
  assign array_update_71678[0] = add_71609 == 32'h0000_0000 ? array_update_71676 : array_update_71668[0];
  assign array_update_71678[1] = add_71609 == 32'h0000_0001 ? array_update_71676 : array_update_71668[1];
  assign array_update_71678[2] = add_71609 == 32'h0000_0002 ? array_update_71676 : array_update_71668[2];
  assign array_update_71678[3] = add_71609 == 32'h0000_0003 ? array_update_71676 : array_update_71668[3];
  assign array_update_71678[4] = add_71609 == 32'h0000_0004 ? array_update_71676 : array_update_71668[4];
  assign array_update_71678[5] = add_71609 == 32'h0000_0005 ? array_update_71676 : array_update_71668[5];
  assign array_update_71678[6] = add_71609 == 32'h0000_0006 ? array_update_71676 : array_update_71668[6];
  assign array_update_71678[7] = add_71609 == 32'h0000_0007 ? array_update_71676 : array_update_71668[7];
  assign array_update_71678[8] = add_71609 == 32'h0000_0008 ? array_update_71676 : array_update_71668[8];
  assign array_update_71678[9] = add_71609 == 32'h0000_0009 ? array_update_71676 : array_update_71668[9];
  assign array_update_71680[0] = add_71611 == 32'h0000_0000 ? array_update_71677 : array_update_71670[0];
  assign array_update_71680[1] = add_71611 == 32'h0000_0001 ? array_update_71677 : array_update_71670[1];
  assign array_update_71680[2] = add_71611 == 32'h0000_0002 ? array_update_71677 : array_update_71670[2];
  assign array_update_71680[3] = add_71611 == 32'h0000_0003 ? array_update_71677 : array_update_71670[3];
  assign array_update_71680[4] = add_71611 == 32'h0000_0004 ? array_update_71677 : array_update_71670[4];
  assign array_update_71680[5] = add_71611 == 32'h0000_0005 ? array_update_71677 : array_update_71670[5];
  assign array_update_71680[6] = add_71611 == 32'h0000_0006 ? array_update_71677 : array_update_71670[6];
  assign array_update_71680[7] = add_71611 == 32'h0000_0007 ? array_update_71677 : array_update_71670[7];
  assign array_update_71680[8] = add_71611 == 32'h0000_0008 ? array_update_71677 : array_update_71670[8];
  assign array_update_71680[9] = add_71611 == 32'h0000_0009 ? array_update_71677 : array_update_71670[9];
  assign array_index_71682 = array_update_71678[add_71609 > 32'h0000_0009 ? 4'h9 : add_71609[3:0]];
  assign add_71683 = add_71673 + 32'h0000_0001;
  assign array_index_71684 = array_update_71680[add_71611 > 32'h0000_0009 ? 4'h9 : add_71611[3:0]];
  assign add_71685 = add_71675 + 32'h0000_0001;
  assign array_update_71686[0] = add_71683 == 32'h0000_0000 ? TestBlock__A_op67 : array_index_71682[0];
  assign array_update_71686[1] = add_71683 == 32'h0000_0001 ? TestBlock__A_op67 : array_index_71682[1];
  assign array_update_71686[2] = add_71683 == 32'h0000_0002 ? TestBlock__A_op67 : array_index_71682[2];
  assign array_update_71686[3] = add_71683 == 32'h0000_0003 ? TestBlock__A_op67 : array_index_71682[3];
  assign array_update_71686[4] = add_71683 == 32'h0000_0004 ? TestBlock__A_op67 : array_index_71682[4];
  assign array_update_71686[5] = add_71683 == 32'h0000_0005 ? TestBlock__A_op67 : array_index_71682[5];
  assign array_update_71686[6] = add_71683 == 32'h0000_0006 ? TestBlock__A_op67 : array_index_71682[6];
  assign array_update_71686[7] = add_71683 == 32'h0000_0007 ? TestBlock__A_op67 : array_index_71682[7];
  assign array_update_71686[8] = add_71683 == 32'h0000_0008 ? TestBlock__A_op67 : array_index_71682[8];
  assign array_update_71686[9] = add_71683 == 32'h0000_0009 ? TestBlock__A_op67 : array_index_71682[9];
  assign array_update_71687[0] = add_71685 == 32'h0000_0000 ? TestBlock__B_op67 : array_index_71684[0];
  assign array_update_71687[1] = add_71685 == 32'h0000_0001 ? TestBlock__B_op67 : array_index_71684[1];
  assign array_update_71687[2] = add_71685 == 32'h0000_0002 ? TestBlock__B_op67 : array_index_71684[2];
  assign array_update_71687[3] = add_71685 == 32'h0000_0003 ? TestBlock__B_op67 : array_index_71684[3];
  assign array_update_71687[4] = add_71685 == 32'h0000_0004 ? TestBlock__B_op67 : array_index_71684[4];
  assign array_update_71687[5] = add_71685 == 32'h0000_0005 ? TestBlock__B_op67 : array_index_71684[5];
  assign array_update_71687[6] = add_71685 == 32'h0000_0006 ? TestBlock__B_op67 : array_index_71684[6];
  assign array_update_71687[7] = add_71685 == 32'h0000_0007 ? TestBlock__B_op67 : array_index_71684[7];
  assign array_update_71687[8] = add_71685 == 32'h0000_0008 ? TestBlock__B_op67 : array_index_71684[8];
  assign array_update_71687[9] = add_71685 == 32'h0000_0009 ? TestBlock__B_op67 : array_index_71684[9];
  assign array_update_71688[0] = add_71609 == 32'h0000_0000 ? array_update_71686 : array_update_71678[0];
  assign array_update_71688[1] = add_71609 == 32'h0000_0001 ? array_update_71686 : array_update_71678[1];
  assign array_update_71688[2] = add_71609 == 32'h0000_0002 ? array_update_71686 : array_update_71678[2];
  assign array_update_71688[3] = add_71609 == 32'h0000_0003 ? array_update_71686 : array_update_71678[3];
  assign array_update_71688[4] = add_71609 == 32'h0000_0004 ? array_update_71686 : array_update_71678[4];
  assign array_update_71688[5] = add_71609 == 32'h0000_0005 ? array_update_71686 : array_update_71678[5];
  assign array_update_71688[6] = add_71609 == 32'h0000_0006 ? array_update_71686 : array_update_71678[6];
  assign array_update_71688[7] = add_71609 == 32'h0000_0007 ? array_update_71686 : array_update_71678[7];
  assign array_update_71688[8] = add_71609 == 32'h0000_0008 ? array_update_71686 : array_update_71678[8];
  assign array_update_71688[9] = add_71609 == 32'h0000_0009 ? array_update_71686 : array_update_71678[9];
  assign array_update_71690[0] = add_71611 == 32'h0000_0000 ? array_update_71687 : array_update_71680[0];
  assign array_update_71690[1] = add_71611 == 32'h0000_0001 ? array_update_71687 : array_update_71680[1];
  assign array_update_71690[2] = add_71611 == 32'h0000_0002 ? array_update_71687 : array_update_71680[2];
  assign array_update_71690[3] = add_71611 == 32'h0000_0003 ? array_update_71687 : array_update_71680[3];
  assign array_update_71690[4] = add_71611 == 32'h0000_0004 ? array_update_71687 : array_update_71680[4];
  assign array_update_71690[5] = add_71611 == 32'h0000_0005 ? array_update_71687 : array_update_71680[5];
  assign array_update_71690[6] = add_71611 == 32'h0000_0006 ? array_update_71687 : array_update_71680[6];
  assign array_update_71690[7] = add_71611 == 32'h0000_0007 ? array_update_71687 : array_update_71680[7];
  assign array_update_71690[8] = add_71611 == 32'h0000_0008 ? array_update_71687 : array_update_71680[8];
  assign array_update_71690[9] = add_71611 == 32'h0000_0009 ? array_update_71687 : array_update_71680[9];
  assign array_index_71692 = array_update_71688[add_71609 > 32'h0000_0009 ? 4'h9 : add_71609[3:0]];
  assign add_71693 = add_71683 + 32'h0000_0001;
  assign array_index_71694 = array_update_71690[add_71611 > 32'h0000_0009 ? 4'h9 : add_71611[3:0]];
  assign add_71695 = add_71685 + 32'h0000_0001;
  assign array_update_71696[0] = add_71693 == 32'h0000_0000 ? TestBlock__A_op68 : array_index_71692[0];
  assign array_update_71696[1] = add_71693 == 32'h0000_0001 ? TestBlock__A_op68 : array_index_71692[1];
  assign array_update_71696[2] = add_71693 == 32'h0000_0002 ? TestBlock__A_op68 : array_index_71692[2];
  assign array_update_71696[3] = add_71693 == 32'h0000_0003 ? TestBlock__A_op68 : array_index_71692[3];
  assign array_update_71696[4] = add_71693 == 32'h0000_0004 ? TestBlock__A_op68 : array_index_71692[4];
  assign array_update_71696[5] = add_71693 == 32'h0000_0005 ? TestBlock__A_op68 : array_index_71692[5];
  assign array_update_71696[6] = add_71693 == 32'h0000_0006 ? TestBlock__A_op68 : array_index_71692[6];
  assign array_update_71696[7] = add_71693 == 32'h0000_0007 ? TestBlock__A_op68 : array_index_71692[7];
  assign array_update_71696[8] = add_71693 == 32'h0000_0008 ? TestBlock__A_op68 : array_index_71692[8];
  assign array_update_71696[9] = add_71693 == 32'h0000_0009 ? TestBlock__A_op68 : array_index_71692[9];
  assign array_update_71697[0] = add_71695 == 32'h0000_0000 ? TestBlock__B_op68 : array_index_71694[0];
  assign array_update_71697[1] = add_71695 == 32'h0000_0001 ? TestBlock__B_op68 : array_index_71694[1];
  assign array_update_71697[2] = add_71695 == 32'h0000_0002 ? TestBlock__B_op68 : array_index_71694[2];
  assign array_update_71697[3] = add_71695 == 32'h0000_0003 ? TestBlock__B_op68 : array_index_71694[3];
  assign array_update_71697[4] = add_71695 == 32'h0000_0004 ? TestBlock__B_op68 : array_index_71694[4];
  assign array_update_71697[5] = add_71695 == 32'h0000_0005 ? TestBlock__B_op68 : array_index_71694[5];
  assign array_update_71697[6] = add_71695 == 32'h0000_0006 ? TestBlock__B_op68 : array_index_71694[6];
  assign array_update_71697[7] = add_71695 == 32'h0000_0007 ? TestBlock__B_op68 : array_index_71694[7];
  assign array_update_71697[8] = add_71695 == 32'h0000_0008 ? TestBlock__B_op68 : array_index_71694[8];
  assign array_update_71697[9] = add_71695 == 32'h0000_0009 ? TestBlock__B_op68 : array_index_71694[9];
  assign array_update_71698[0] = add_71609 == 32'h0000_0000 ? array_update_71696 : array_update_71688[0];
  assign array_update_71698[1] = add_71609 == 32'h0000_0001 ? array_update_71696 : array_update_71688[1];
  assign array_update_71698[2] = add_71609 == 32'h0000_0002 ? array_update_71696 : array_update_71688[2];
  assign array_update_71698[3] = add_71609 == 32'h0000_0003 ? array_update_71696 : array_update_71688[3];
  assign array_update_71698[4] = add_71609 == 32'h0000_0004 ? array_update_71696 : array_update_71688[4];
  assign array_update_71698[5] = add_71609 == 32'h0000_0005 ? array_update_71696 : array_update_71688[5];
  assign array_update_71698[6] = add_71609 == 32'h0000_0006 ? array_update_71696 : array_update_71688[6];
  assign array_update_71698[7] = add_71609 == 32'h0000_0007 ? array_update_71696 : array_update_71688[7];
  assign array_update_71698[8] = add_71609 == 32'h0000_0008 ? array_update_71696 : array_update_71688[8];
  assign array_update_71698[9] = add_71609 == 32'h0000_0009 ? array_update_71696 : array_update_71688[9];
  assign array_update_71700[0] = add_71611 == 32'h0000_0000 ? array_update_71697 : array_update_71690[0];
  assign array_update_71700[1] = add_71611 == 32'h0000_0001 ? array_update_71697 : array_update_71690[1];
  assign array_update_71700[2] = add_71611 == 32'h0000_0002 ? array_update_71697 : array_update_71690[2];
  assign array_update_71700[3] = add_71611 == 32'h0000_0003 ? array_update_71697 : array_update_71690[3];
  assign array_update_71700[4] = add_71611 == 32'h0000_0004 ? array_update_71697 : array_update_71690[4];
  assign array_update_71700[5] = add_71611 == 32'h0000_0005 ? array_update_71697 : array_update_71690[5];
  assign array_update_71700[6] = add_71611 == 32'h0000_0006 ? array_update_71697 : array_update_71690[6];
  assign array_update_71700[7] = add_71611 == 32'h0000_0007 ? array_update_71697 : array_update_71690[7];
  assign array_update_71700[8] = add_71611 == 32'h0000_0008 ? array_update_71697 : array_update_71690[8];
  assign array_update_71700[9] = add_71611 == 32'h0000_0009 ? array_update_71697 : array_update_71690[9];
  assign array_index_71702 = array_update_71698[add_71609 > 32'h0000_0009 ? 4'h9 : add_71609[3:0]];
  assign add_71703 = add_71693 + 32'h0000_0001;
  assign array_index_71704 = array_update_71700[add_71611 > 32'h0000_0009 ? 4'h9 : add_71611[3:0]];
  assign add_71705 = add_71695 + 32'h0000_0001;
  assign array_update_71706[0] = add_71703 == 32'h0000_0000 ? TestBlock__A_op69 : array_index_71702[0];
  assign array_update_71706[1] = add_71703 == 32'h0000_0001 ? TestBlock__A_op69 : array_index_71702[1];
  assign array_update_71706[2] = add_71703 == 32'h0000_0002 ? TestBlock__A_op69 : array_index_71702[2];
  assign array_update_71706[3] = add_71703 == 32'h0000_0003 ? TestBlock__A_op69 : array_index_71702[3];
  assign array_update_71706[4] = add_71703 == 32'h0000_0004 ? TestBlock__A_op69 : array_index_71702[4];
  assign array_update_71706[5] = add_71703 == 32'h0000_0005 ? TestBlock__A_op69 : array_index_71702[5];
  assign array_update_71706[6] = add_71703 == 32'h0000_0006 ? TestBlock__A_op69 : array_index_71702[6];
  assign array_update_71706[7] = add_71703 == 32'h0000_0007 ? TestBlock__A_op69 : array_index_71702[7];
  assign array_update_71706[8] = add_71703 == 32'h0000_0008 ? TestBlock__A_op69 : array_index_71702[8];
  assign array_update_71706[9] = add_71703 == 32'h0000_0009 ? TestBlock__A_op69 : array_index_71702[9];
  assign array_update_71708[0] = add_71705 == 32'h0000_0000 ? TestBlock__B_op69 : array_index_71704[0];
  assign array_update_71708[1] = add_71705 == 32'h0000_0001 ? TestBlock__B_op69 : array_index_71704[1];
  assign array_update_71708[2] = add_71705 == 32'h0000_0002 ? TestBlock__B_op69 : array_index_71704[2];
  assign array_update_71708[3] = add_71705 == 32'h0000_0003 ? TestBlock__B_op69 : array_index_71704[3];
  assign array_update_71708[4] = add_71705 == 32'h0000_0004 ? TestBlock__B_op69 : array_index_71704[4];
  assign array_update_71708[5] = add_71705 == 32'h0000_0005 ? TestBlock__B_op69 : array_index_71704[5];
  assign array_update_71708[6] = add_71705 == 32'h0000_0006 ? TestBlock__B_op69 : array_index_71704[6];
  assign array_update_71708[7] = add_71705 == 32'h0000_0007 ? TestBlock__B_op69 : array_index_71704[7];
  assign array_update_71708[8] = add_71705 == 32'h0000_0008 ? TestBlock__B_op69 : array_index_71704[8];
  assign array_update_71708[9] = add_71705 == 32'h0000_0009 ? TestBlock__B_op69 : array_index_71704[9];
  assign array_update_71710[0] = add_71609 == 32'h0000_0000 ? array_update_71706 : array_update_71698[0];
  assign array_update_71710[1] = add_71609 == 32'h0000_0001 ? array_update_71706 : array_update_71698[1];
  assign array_update_71710[2] = add_71609 == 32'h0000_0002 ? array_update_71706 : array_update_71698[2];
  assign array_update_71710[3] = add_71609 == 32'h0000_0003 ? array_update_71706 : array_update_71698[3];
  assign array_update_71710[4] = add_71609 == 32'h0000_0004 ? array_update_71706 : array_update_71698[4];
  assign array_update_71710[5] = add_71609 == 32'h0000_0005 ? array_update_71706 : array_update_71698[5];
  assign array_update_71710[6] = add_71609 == 32'h0000_0006 ? array_update_71706 : array_update_71698[6];
  assign array_update_71710[7] = add_71609 == 32'h0000_0007 ? array_update_71706 : array_update_71698[7];
  assign array_update_71710[8] = add_71609 == 32'h0000_0008 ? array_update_71706 : array_update_71698[8];
  assign array_update_71710[9] = add_71609 == 32'h0000_0009 ? array_update_71706 : array_update_71698[9];
  assign add_71711 = add_71609 + 32'h0000_0001;
  assign array_update_71712[0] = add_71611 == 32'h0000_0000 ? array_update_71708 : array_update_71700[0];
  assign array_update_71712[1] = add_71611 == 32'h0000_0001 ? array_update_71708 : array_update_71700[1];
  assign array_update_71712[2] = add_71611 == 32'h0000_0002 ? array_update_71708 : array_update_71700[2];
  assign array_update_71712[3] = add_71611 == 32'h0000_0003 ? array_update_71708 : array_update_71700[3];
  assign array_update_71712[4] = add_71611 == 32'h0000_0004 ? array_update_71708 : array_update_71700[4];
  assign array_update_71712[5] = add_71611 == 32'h0000_0005 ? array_update_71708 : array_update_71700[5];
  assign array_update_71712[6] = add_71611 == 32'h0000_0006 ? array_update_71708 : array_update_71700[6];
  assign array_update_71712[7] = add_71611 == 32'h0000_0007 ? array_update_71708 : array_update_71700[7];
  assign array_update_71712[8] = add_71611 == 32'h0000_0008 ? array_update_71708 : array_update_71700[8];
  assign array_update_71712[9] = add_71611 == 32'h0000_0009 ? array_update_71708 : array_update_71700[9];
  assign add_71713 = add_71611 + 32'h0000_0001;
  assign array_index_71714 = array_update_71710[add_71711 > 32'h0000_0009 ? 4'h9 : add_71711[3:0]];
  assign literal_71715 = 32'h0000_0000;
  assign array_index_71716 = array_update_71712[add_71713 > 32'h0000_0009 ? 4'h9 : add_71713[3:0]];
  assign literal_71717 = 32'h0000_0000;
  assign array_update_71718[0] = literal_71715 == 32'h0000_0000 ? TestBlock__A_op70 : array_index_71714[0];
  assign array_update_71718[1] = literal_71715 == 32'h0000_0001 ? TestBlock__A_op70 : array_index_71714[1];
  assign array_update_71718[2] = literal_71715 == 32'h0000_0002 ? TestBlock__A_op70 : array_index_71714[2];
  assign array_update_71718[3] = literal_71715 == 32'h0000_0003 ? TestBlock__A_op70 : array_index_71714[3];
  assign array_update_71718[4] = literal_71715 == 32'h0000_0004 ? TestBlock__A_op70 : array_index_71714[4];
  assign array_update_71718[5] = literal_71715 == 32'h0000_0005 ? TestBlock__A_op70 : array_index_71714[5];
  assign array_update_71718[6] = literal_71715 == 32'h0000_0006 ? TestBlock__A_op70 : array_index_71714[6];
  assign array_update_71718[7] = literal_71715 == 32'h0000_0007 ? TestBlock__A_op70 : array_index_71714[7];
  assign array_update_71718[8] = literal_71715 == 32'h0000_0008 ? TestBlock__A_op70 : array_index_71714[8];
  assign array_update_71718[9] = literal_71715 == 32'h0000_0009 ? TestBlock__A_op70 : array_index_71714[9];
  assign array_update_71719[0] = literal_71717 == 32'h0000_0000 ? TestBlock__B_op70 : array_index_71716[0];
  assign array_update_71719[1] = literal_71717 == 32'h0000_0001 ? TestBlock__B_op70 : array_index_71716[1];
  assign array_update_71719[2] = literal_71717 == 32'h0000_0002 ? TestBlock__B_op70 : array_index_71716[2];
  assign array_update_71719[3] = literal_71717 == 32'h0000_0003 ? TestBlock__B_op70 : array_index_71716[3];
  assign array_update_71719[4] = literal_71717 == 32'h0000_0004 ? TestBlock__B_op70 : array_index_71716[4];
  assign array_update_71719[5] = literal_71717 == 32'h0000_0005 ? TestBlock__B_op70 : array_index_71716[5];
  assign array_update_71719[6] = literal_71717 == 32'h0000_0006 ? TestBlock__B_op70 : array_index_71716[6];
  assign array_update_71719[7] = literal_71717 == 32'h0000_0007 ? TestBlock__B_op70 : array_index_71716[7];
  assign array_update_71719[8] = literal_71717 == 32'h0000_0008 ? TestBlock__B_op70 : array_index_71716[8];
  assign array_update_71719[9] = literal_71717 == 32'h0000_0009 ? TestBlock__B_op70 : array_index_71716[9];
  assign array_update_71720[0] = add_71711 == 32'h0000_0000 ? array_update_71718 : array_update_71710[0];
  assign array_update_71720[1] = add_71711 == 32'h0000_0001 ? array_update_71718 : array_update_71710[1];
  assign array_update_71720[2] = add_71711 == 32'h0000_0002 ? array_update_71718 : array_update_71710[2];
  assign array_update_71720[3] = add_71711 == 32'h0000_0003 ? array_update_71718 : array_update_71710[3];
  assign array_update_71720[4] = add_71711 == 32'h0000_0004 ? array_update_71718 : array_update_71710[4];
  assign array_update_71720[5] = add_71711 == 32'h0000_0005 ? array_update_71718 : array_update_71710[5];
  assign array_update_71720[6] = add_71711 == 32'h0000_0006 ? array_update_71718 : array_update_71710[6];
  assign array_update_71720[7] = add_71711 == 32'h0000_0007 ? array_update_71718 : array_update_71710[7];
  assign array_update_71720[8] = add_71711 == 32'h0000_0008 ? array_update_71718 : array_update_71710[8];
  assign array_update_71720[9] = add_71711 == 32'h0000_0009 ? array_update_71718 : array_update_71710[9];
  assign array_update_71722[0] = add_71713 == 32'h0000_0000 ? array_update_71719 : array_update_71712[0];
  assign array_update_71722[1] = add_71713 == 32'h0000_0001 ? array_update_71719 : array_update_71712[1];
  assign array_update_71722[2] = add_71713 == 32'h0000_0002 ? array_update_71719 : array_update_71712[2];
  assign array_update_71722[3] = add_71713 == 32'h0000_0003 ? array_update_71719 : array_update_71712[3];
  assign array_update_71722[4] = add_71713 == 32'h0000_0004 ? array_update_71719 : array_update_71712[4];
  assign array_update_71722[5] = add_71713 == 32'h0000_0005 ? array_update_71719 : array_update_71712[5];
  assign array_update_71722[6] = add_71713 == 32'h0000_0006 ? array_update_71719 : array_update_71712[6];
  assign array_update_71722[7] = add_71713 == 32'h0000_0007 ? array_update_71719 : array_update_71712[7];
  assign array_update_71722[8] = add_71713 == 32'h0000_0008 ? array_update_71719 : array_update_71712[8];
  assign array_update_71722[9] = add_71713 == 32'h0000_0009 ? array_update_71719 : array_update_71712[9];
  assign array_index_71724 = array_update_71720[add_71711 > 32'h0000_0009 ? 4'h9 : add_71711[3:0]];
  assign add_71725 = literal_71715 + 32'h0000_0001;
  assign array_index_71726 = array_update_71722[add_71713 > 32'h0000_0009 ? 4'h9 : add_71713[3:0]];
  assign add_71727 = literal_71717 + 32'h0000_0001;
  assign array_update_71728[0] = add_71725 == 32'h0000_0000 ? TestBlock__A_op71 : array_index_71724[0];
  assign array_update_71728[1] = add_71725 == 32'h0000_0001 ? TestBlock__A_op71 : array_index_71724[1];
  assign array_update_71728[2] = add_71725 == 32'h0000_0002 ? TestBlock__A_op71 : array_index_71724[2];
  assign array_update_71728[3] = add_71725 == 32'h0000_0003 ? TestBlock__A_op71 : array_index_71724[3];
  assign array_update_71728[4] = add_71725 == 32'h0000_0004 ? TestBlock__A_op71 : array_index_71724[4];
  assign array_update_71728[5] = add_71725 == 32'h0000_0005 ? TestBlock__A_op71 : array_index_71724[5];
  assign array_update_71728[6] = add_71725 == 32'h0000_0006 ? TestBlock__A_op71 : array_index_71724[6];
  assign array_update_71728[7] = add_71725 == 32'h0000_0007 ? TestBlock__A_op71 : array_index_71724[7];
  assign array_update_71728[8] = add_71725 == 32'h0000_0008 ? TestBlock__A_op71 : array_index_71724[8];
  assign array_update_71728[9] = add_71725 == 32'h0000_0009 ? TestBlock__A_op71 : array_index_71724[9];
  assign array_update_71729[0] = add_71727 == 32'h0000_0000 ? TestBlock__B_op71 : array_index_71726[0];
  assign array_update_71729[1] = add_71727 == 32'h0000_0001 ? TestBlock__B_op71 : array_index_71726[1];
  assign array_update_71729[2] = add_71727 == 32'h0000_0002 ? TestBlock__B_op71 : array_index_71726[2];
  assign array_update_71729[3] = add_71727 == 32'h0000_0003 ? TestBlock__B_op71 : array_index_71726[3];
  assign array_update_71729[4] = add_71727 == 32'h0000_0004 ? TestBlock__B_op71 : array_index_71726[4];
  assign array_update_71729[5] = add_71727 == 32'h0000_0005 ? TestBlock__B_op71 : array_index_71726[5];
  assign array_update_71729[6] = add_71727 == 32'h0000_0006 ? TestBlock__B_op71 : array_index_71726[6];
  assign array_update_71729[7] = add_71727 == 32'h0000_0007 ? TestBlock__B_op71 : array_index_71726[7];
  assign array_update_71729[8] = add_71727 == 32'h0000_0008 ? TestBlock__B_op71 : array_index_71726[8];
  assign array_update_71729[9] = add_71727 == 32'h0000_0009 ? TestBlock__B_op71 : array_index_71726[9];
  assign array_update_71730[0] = add_71711 == 32'h0000_0000 ? array_update_71728 : array_update_71720[0];
  assign array_update_71730[1] = add_71711 == 32'h0000_0001 ? array_update_71728 : array_update_71720[1];
  assign array_update_71730[2] = add_71711 == 32'h0000_0002 ? array_update_71728 : array_update_71720[2];
  assign array_update_71730[3] = add_71711 == 32'h0000_0003 ? array_update_71728 : array_update_71720[3];
  assign array_update_71730[4] = add_71711 == 32'h0000_0004 ? array_update_71728 : array_update_71720[4];
  assign array_update_71730[5] = add_71711 == 32'h0000_0005 ? array_update_71728 : array_update_71720[5];
  assign array_update_71730[6] = add_71711 == 32'h0000_0006 ? array_update_71728 : array_update_71720[6];
  assign array_update_71730[7] = add_71711 == 32'h0000_0007 ? array_update_71728 : array_update_71720[7];
  assign array_update_71730[8] = add_71711 == 32'h0000_0008 ? array_update_71728 : array_update_71720[8];
  assign array_update_71730[9] = add_71711 == 32'h0000_0009 ? array_update_71728 : array_update_71720[9];
  assign array_update_71732[0] = add_71713 == 32'h0000_0000 ? array_update_71729 : array_update_71722[0];
  assign array_update_71732[1] = add_71713 == 32'h0000_0001 ? array_update_71729 : array_update_71722[1];
  assign array_update_71732[2] = add_71713 == 32'h0000_0002 ? array_update_71729 : array_update_71722[2];
  assign array_update_71732[3] = add_71713 == 32'h0000_0003 ? array_update_71729 : array_update_71722[3];
  assign array_update_71732[4] = add_71713 == 32'h0000_0004 ? array_update_71729 : array_update_71722[4];
  assign array_update_71732[5] = add_71713 == 32'h0000_0005 ? array_update_71729 : array_update_71722[5];
  assign array_update_71732[6] = add_71713 == 32'h0000_0006 ? array_update_71729 : array_update_71722[6];
  assign array_update_71732[7] = add_71713 == 32'h0000_0007 ? array_update_71729 : array_update_71722[7];
  assign array_update_71732[8] = add_71713 == 32'h0000_0008 ? array_update_71729 : array_update_71722[8];
  assign array_update_71732[9] = add_71713 == 32'h0000_0009 ? array_update_71729 : array_update_71722[9];
  assign array_index_71734 = array_update_71730[add_71711 > 32'h0000_0009 ? 4'h9 : add_71711[3:0]];
  assign add_71735 = add_71725 + 32'h0000_0001;
  assign array_index_71736 = array_update_71732[add_71713 > 32'h0000_0009 ? 4'h9 : add_71713[3:0]];
  assign add_71737 = add_71727 + 32'h0000_0001;
  assign array_update_71738[0] = add_71735 == 32'h0000_0000 ? TestBlock__A_op72 : array_index_71734[0];
  assign array_update_71738[1] = add_71735 == 32'h0000_0001 ? TestBlock__A_op72 : array_index_71734[1];
  assign array_update_71738[2] = add_71735 == 32'h0000_0002 ? TestBlock__A_op72 : array_index_71734[2];
  assign array_update_71738[3] = add_71735 == 32'h0000_0003 ? TestBlock__A_op72 : array_index_71734[3];
  assign array_update_71738[4] = add_71735 == 32'h0000_0004 ? TestBlock__A_op72 : array_index_71734[4];
  assign array_update_71738[5] = add_71735 == 32'h0000_0005 ? TestBlock__A_op72 : array_index_71734[5];
  assign array_update_71738[6] = add_71735 == 32'h0000_0006 ? TestBlock__A_op72 : array_index_71734[6];
  assign array_update_71738[7] = add_71735 == 32'h0000_0007 ? TestBlock__A_op72 : array_index_71734[7];
  assign array_update_71738[8] = add_71735 == 32'h0000_0008 ? TestBlock__A_op72 : array_index_71734[8];
  assign array_update_71738[9] = add_71735 == 32'h0000_0009 ? TestBlock__A_op72 : array_index_71734[9];
  assign array_update_71739[0] = add_71737 == 32'h0000_0000 ? TestBlock__B_op72 : array_index_71736[0];
  assign array_update_71739[1] = add_71737 == 32'h0000_0001 ? TestBlock__B_op72 : array_index_71736[1];
  assign array_update_71739[2] = add_71737 == 32'h0000_0002 ? TestBlock__B_op72 : array_index_71736[2];
  assign array_update_71739[3] = add_71737 == 32'h0000_0003 ? TestBlock__B_op72 : array_index_71736[3];
  assign array_update_71739[4] = add_71737 == 32'h0000_0004 ? TestBlock__B_op72 : array_index_71736[4];
  assign array_update_71739[5] = add_71737 == 32'h0000_0005 ? TestBlock__B_op72 : array_index_71736[5];
  assign array_update_71739[6] = add_71737 == 32'h0000_0006 ? TestBlock__B_op72 : array_index_71736[6];
  assign array_update_71739[7] = add_71737 == 32'h0000_0007 ? TestBlock__B_op72 : array_index_71736[7];
  assign array_update_71739[8] = add_71737 == 32'h0000_0008 ? TestBlock__B_op72 : array_index_71736[8];
  assign array_update_71739[9] = add_71737 == 32'h0000_0009 ? TestBlock__B_op72 : array_index_71736[9];
  assign array_update_71740[0] = add_71711 == 32'h0000_0000 ? array_update_71738 : array_update_71730[0];
  assign array_update_71740[1] = add_71711 == 32'h0000_0001 ? array_update_71738 : array_update_71730[1];
  assign array_update_71740[2] = add_71711 == 32'h0000_0002 ? array_update_71738 : array_update_71730[2];
  assign array_update_71740[3] = add_71711 == 32'h0000_0003 ? array_update_71738 : array_update_71730[3];
  assign array_update_71740[4] = add_71711 == 32'h0000_0004 ? array_update_71738 : array_update_71730[4];
  assign array_update_71740[5] = add_71711 == 32'h0000_0005 ? array_update_71738 : array_update_71730[5];
  assign array_update_71740[6] = add_71711 == 32'h0000_0006 ? array_update_71738 : array_update_71730[6];
  assign array_update_71740[7] = add_71711 == 32'h0000_0007 ? array_update_71738 : array_update_71730[7];
  assign array_update_71740[8] = add_71711 == 32'h0000_0008 ? array_update_71738 : array_update_71730[8];
  assign array_update_71740[9] = add_71711 == 32'h0000_0009 ? array_update_71738 : array_update_71730[9];
  assign array_update_71742[0] = add_71713 == 32'h0000_0000 ? array_update_71739 : array_update_71732[0];
  assign array_update_71742[1] = add_71713 == 32'h0000_0001 ? array_update_71739 : array_update_71732[1];
  assign array_update_71742[2] = add_71713 == 32'h0000_0002 ? array_update_71739 : array_update_71732[2];
  assign array_update_71742[3] = add_71713 == 32'h0000_0003 ? array_update_71739 : array_update_71732[3];
  assign array_update_71742[4] = add_71713 == 32'h0000_0004 ? array_update_71739 : array_update_71732[4];
  assign array_update_71742[5] = add_71713 == 32'h0000_0005 ? array_update_71739 : array_update_71732[5];
  assign array_update_71742[6] = add_71713 == 32'h0000_0006 ? array_update_71739 : array_update_71732[6];
  assign array_update_71742[7] = add_71713 == 32'h0000_0007 ? array_update_71739 : array_update_71732[7];
  assign array_update_71742[8] = add_71713 == 32'h0000_0008 ? array_update_71739 : array_update_71732[8];
  assign array_update_71742[9] = add_71713 == 32'h0000_0009 ? array_update_71739 : array_update_71732[9];
  assign array_index_71744 = array_update_71740[add_71711 > 32'h0000_0009 ? 4'h9 : add_71711[3:0]];
  assign add_71745 = add_71735 + 32'h0000_0001;
  assign array_index_71746 = array_update_71742[add_71713 > 32'h0000_0009 ? 4'h9 : add_71713[3:0]];
  assign add_71747 = add_71737 + 32'h0000_0001;
  assign array_update_71748[0] = add_71745 == 32'h0000_0000 ? TestBlock__A_op73 : array_index_71744[0];
  assign array_update_71748[1] = add_71745 == 32'h0000_0001 ? TestBlock__A_op73 : array_index_71744[1];
  assign array_update_71748[2] = add_71745 == 32'h0000_0002 ? TestBlock__A_op73 : array_index_71744[2];
  assign array_update_71748[3] = add_71745 == 32'h0000_0003 ? TestBlock__A_op73 : array_index_71744[3];
  assign array_update_71748[4] = add_71745 == 32'h0000_0004 ? TestBlock__A_op73 : array_index_71744[4];
  assign array_update_71748[5] = add_71745 == 32'h0000_0005 ? TestBlock__A_op73 : array_index_71744[5];
  assign array_update_71748[6] = add_71745 == 32'h0000_0006 ? TestBlock__A_op73 : array_index_71744[6];
  assign array_update_71748[7] = add_71745 == 32'h0000_0007 ? TestBlock__A_op73 : array_index_71744[7];
  assign array_update_71748[8] = add_71745 == 32'h0000_0008 ? TestBlock__A_op73 : array_index_71744[8];
  assign array_update_71748[9] = add_71745 == 32'h0000_0009 ? TestBlock__A_op73 : array_index_71744[9];
  assign array_update_71749[0] = add_71747 == 32'h0000_0000 ? TestBlock__B_op73 : array_index_71746[0];
  assign array_update_71749[1] = add_71747 == 32'h0000_0001 ? TestBlock__B_op73 : array_index_71746[1];
  assign array_update_71749[2] = add_71747 == 32'h0000_0002 ? TestBlock__B_op73 : array_index_71746[2];
  assign array_update_71749[3] = add_71747 == 32'h0000_0003 ? TestBlock__B_op73 : array_index_71746[3];
  assign array_update_71749[4] = add_71747 == 32'h0000_0004 ? TestBlock__B_op73 : array_index_71746[4];
  assign array_update_71749[5] = add_71747 == 32'h0000_0005 ? TestBlock__B_op73 : array_index_71746[5];
  assign array_update_71749[6] = add_71747 == 32'h0000_0006 ? TestBlock__B_op73 : array_index_71746[6];
  assign array_update_71749[7] = add_71747 == 32'h0000_0007 ? TestBlock__B_op73 : array_index_71746[7];
  assign array_update_71749[8] = add_71747 == 32'h0000_0008 ? TestBlock__B_op73 : array_index_71746[8];
  assign array_update_71749[9] = add_71747 == 32'h0000_0009 ? TestBlock__B_op73 : array_index_71746[9];
  assign array_update_71750[0] = add_71711 == 32'h0000_0000 ? array_update_71748 : array_update_71740[0];
  assign array_update_71750[1] = add_71711 == 32'h0000_0001 ? array_update_71748 : array_update_71740[1];
  assign array_update_71750[2] = add_71711 == 32'h0000_0002 ? array_update_71748 : array_update_71740[2];
  assign array_update_71750[3] = add_71711 == 32'h0000_0003 ? array_update_71748 : array_update_71740[3];
  assign array_update_71750[4] = add_71711 == 32'h0000_0004 ? array_update_71748 : array_update_71740[4];
  assign array_update_71750[5] = add_71711 == 32'h0000_0005 ? array_update_71748 : array_update_71740[5];
  assign array_update_71750[6] = add_71711 == 32'h0000_0006 ? array_update_71748 : array_update_71740[6];
  assign array_update_71750[7] = add_71711 == 32'h0000_0007 ? array_update_71748 : array_update_71740[7];
  assign array_update_71750[8] = add_71711 == 32'h0000_0008 ? array_update_71748 : array_update_71740[8];
  assign array_update_71750[9] = add_71711 == 32'h0000_0009 ? array_update_71748 : array_update_71740[9];
  assign array_update_71752[0] = add_71713 == 32'h0000_0000 ? array_update_71749 : array_update_71742[0];
  assign array_update_71752[1] = add_71713 == 32'h0000_0001 ? array_update_71749 : array_update_71742[1];
  assign array_update_71752[2] = add_71713 == 32'h0000_0002 ? array_update_71749 : array_update_71742[2];
  assign array_update_71752[3] = add_71713 == 32'h0000_0003 ? array_update_71749 : array_update_71742[3];
  assign array_update_71752[4] = add_71713 == 32'h0000_0004 ? array_update_71749 : array_update_71742[4];
  assign array_update_71752[5] = add_71713 == 32'h0000_0005 ? array_update_71749 : array_update_71742[5];
  assign array_update_71752[6] = add_71713 == 32'h0000_0006 ? array_update_71749 : array_update_71742[6];
  assign array_update_71752[7] = add_71713 == 32'h0000_0007 ? array_update_71749 : array_update_71742[7];
  assign array_update_71752[8] = add_71713 == 32'h0000_0008 ? array_update_71749 : array_update_71742[8];
  assign array_update_71752[9] = add_71713 == 32'h0000_0009 ? array_update_71749 : array_update_71742[9];
  assign array_index_71754 = array_update_71750[add_71711 > 32'h0000_0009 ? 4'h9 : add_71711[3:0]];
  assign add_71755 = add_71745 + 32'h0000_0001;
  assign array_index_71756 = array_update_71752[add_71713 > 32'h0000_0009 ? 4'h9 : add_71713[3:0]];
  assign add_71757 = add_71747 + 32'h0000_0001;
  assign array_update_71758[0] = add_71755 == 32'h0000_0000 ? TestBlock__A_op74 : array_index_71754[0];
  assign array_update_71758[1] = add_71755 == 32'h0000_0001 ? TestBlock__A_op74 : array_index_71754[1];
  assign array_update_71758[2] = add_71755 == 32'h0000_0002 ? TestBlock__A_op74 : array_index_71754[2];
  assign array_update_71758[3] = add_71755 == 32'h0000_0003 ? TestBlock__A_op74 : array_index_71754[3];
  assign array_update_71758[4] = add_71755 == 32'h0000_0004 ? TestBlock__A_op74 : array_index_71754[4];
  assign array_update_71758[5] = add_71755 == 32'h0000_0005 ? TestBlock__A_op74 : array_index_71754[5];
  assign array_update_71758[6] = add_71755 == 32'h0000_0006 ? TestBlock__A_op74 : array_index_71754[6];
  assign array_update_71758[7] = add_71755 == 32'h0000_0007 ? TestBlock__A_op74 : array_index_71754[7];
  assign array_update_71758[8] = add_71755 == 32'h0000_0008 ? TestBlock__A_op74 : array_index_71754[8];
  assign array_update_71758[9] = add_71755 == 32'h0000_0009 ? TestBlock__A_op74 : array_index_71754[9];
  assign array_update_71759[0] = add_71757 == 32'h0000_0000 ? TestBlock__B_op74 : array_index_71756[0];
  assign array_update_71759[1] = add_71757 == 32'h0000_0001 ? TestBlock__B_op74 : array_index_71756[1];
  assign array_update_71759[2] = add_71757 == 32'h0000_0002 ? TestBlock__B_op74 : array_index_71756[2];
  assign array_update_71759[3] = add_71757 == 32'h0000_0003 ? TestBlock__B_op74 : array_index_71756[3];
  assign array_update_71759[4] = add_71757 == 32'h0000_0004 ? TestBlock__B_op74 : array_index_71756[4];
  assign array_update_71759[5] = add_71757 == 32'h0000_0005 ? TestBlock__B_op74 : array_index_71756[5];
  assign array_update_71759[6] = add_71757 == 32'h0000_0006 ? TestBlock__B_op74 : array_index_71756[6];
  assign array_update_71759[7] = add_71757 == 32'h0000_0007 ? TestBlock__B_op74 : array_index_71756[7];
  assign array_update_71759[8] = add_71757 == 32'h0000_0008 ? TestBlock__B_op74 : array_index_71756[8];
  assign array_update_71759[9] = add_71757 == 32'h0000_0009 ? TestBlock__B_op74 : array_index_71756[9];
  assign array_update_71760[0] = add_71711 == 32'h0000_0000 ? array_update_71758 : array_update_71750[0];
  assign array_update_71760[1] = add_71711 == 32'h0000_0001 ? array_update_71758 : array_update_71750[1];
  assign array_update_71760[2] = add_71711 == 32'h0000_0002 ? array_update_71758 : array_update_71750[2];
  assign array_update_71760[3] = add_71711 == 32'h0000_0003 ? array_update_71758 : array_update_71750[3];
  assign array_update_71760[4] = add_71711 == 32'h0000_0004 ? array_update_71758 : array_update_71750[4];
  assign array_update_71760[5] = add_71711 == 32'h0000_0005 ? array_update_71758 : array_update_71750[5];
  assign array_update_71760[6] = add_71711 == 32'h0000_0006 ? array_update_71758 : array_update_71750[6];
  assign array_update_71760[7] = add_71711 == 32'h0000_0007 ? array_update_71758 : array_update_71750[7];
  assign array_update_71760[8] = add_71711 == 32'h0000_0008 ? array_update_71758 : array_update_71750[8];
  assign array_update_71760[9] = add_71711 == 32'h0000_0009 ? array_update_71758 : array_update_71750[9];
  assign array_update_71762[0] = add_71713 == 32'h0000_0000 ? array_update_71759 : array_update_71752[0];
  assign array_update_71762[1] = add_71713 == 32'h0000_0001 ? array_update_71759 : array_update_71752[1];
  assign array_update_71762[2] = add_71713 == 32'h0000_0002 ? array_update_71759 : array_update_71752[2];
  assign array_update_71762[3] = add_71713 == 32'h0000_0003 ? array_update_71759 : array_update_71752[3];
  assign array_update_71762[4] = add_71713 == 32'h0000_0004 ? array_update_71759 : array_update_71752[4];
  assign array_update_71762[5] = add_71713 == 32'h0000_0005 ? array_update_71759 : array_update_71752[5];
  assign array_update_71762[6] = add_71713 == 32'h0000_0006 ? array_update_71759 : array_update_71752[6];
  assign array_update_71762[7] = add_71713 == 32'h0000_0007 ? array_update_71759 : array_update_71752[7];
  assign array_update_71762[8] = add_71713 == 32'h0000_0008 ? array_update_71759 : array_update_71752[8];
  assign array_update_71762[9] = add_71713 == 32'h0000_0009 ? array_update_71759 : array_update_71752[9];
  assign array_index_71764 = array_update_71760[add_71711 > 32'h0000_0009 ? 4'h9 : add_71711[3:0]];
  assign add_71765 = add_71755 + 32'h0000_0001;
  assign array_index_71766 = array_update_71762[add_71713 > 32'h0000_0009 ? 4'h9 : add_71713[3:0]];
  assign add_71767 = add_71757 + 32'h0000_0001;
  assign array_update_71768[0] = add_71765 == 32'h0000_0000 ? TestBlock__A_op75 : array_index_71764[0];
  assign array_update_71768[1] = add_71765 == 32'h0000_0001 ? TestBlock__A_op75 : array_index_71764[1];
  assign array_update_71768[2] = add_71765 == 32'h0000_0002 ? TestBlock__A_op75 : array_index_71764[2];
  assign array_update_71768[3] = add_71765 == 32'h0000_0003 ? TestBlock__A_op75 : array_index_71764[3];
  assign array_update_71768[4] = add_71765 == 32'h0000_0004 ? TestBlock__A_op75 : array_index_71764[4];
  assign array_update_71768[5] = add_71765 == 32'h0000_0005 ? TestBlock__A_op75 : array_index_71764[5];
  assign array_update_71768[6] = add_71765 == 32'h0000_0006 ? TestBlock__A_op75 : array_index_71764[6];
  assign array_update_71768[7] = add_71765 == 32'h0000_0007 ? TestBlock__A_op75 : array_index_71764[7];
  assign array_update_71768[8] = add_71765 == 32'h0000_0008 ? TestBlock__A_op75 : array_index_71764[8];
  assign array_update_71768[9] = add_71765 == 32'h0000_0009 ? TestBlock__A_op75 : array_index_71764[9];
  assign array_update_71769[0] = add_71767 == 32'h0000_0000 ? TestBlock__B_op75 : array_index_71766[0];
  assign array_update_71769[1] = add_71767 == 32'h0000_0001 ? TestBlock__B_op75 : array_index_71766[1];
  assign array_update_71769[2] = add_71767 == 32'h0000_0002 ? TestBlock__B_op75 : array_index_71766[2];
  assign array_update_71769[3] = add_71767 == 32'h0000_0003 ? TestBlock__B_op75 : array_index_71766[3];
  assign array_update_71769[4] = add_71767 == 32'h0000_0004 ? TestBlock__B_op75 : array_index_71766[4];
  assign array_update_71769[5] = add_71767 == 32'h0000_0005 ? TestBlock__B_op75 : array_index_71766[5];
  assign array_update_71769[6] = add_71767 == 32'h0000_0006 ? TestBlock__B_op75 : array_index_71766[6];
  assign array_update_71769[7] = add_71767 == 32'h0000_0007 ? TestBlock__B_op75 : array_index_71766[7];
  assign array_update_71769[8] = add_71767 == 32'h0000_0008 ? TestBlock__B_op75 : array_index_71766[8];
  assign array_update_71769[9] = add_71767 == 32'h0000_0009 ? TestBlock__B_op75 : array_index_71766[9];
  assign array_update_71770[0] = add_71711 == 32'h0000_0000 ? array_update_71768 : array_update_71760[0];
  assign array_update_71770[1] = add_71711 == 32'h0000_0001 ? array_update_71768 : array_update_71760[1];
  assign array_update_71770[2] = add_71711 == 32'h0000_0002 ? array_update_71768 : array_update_71760[2];
  assign array_update_71770[3] = add_71711 == 32'h0000_0003 ? array_update_71768 : array_update_71760[3];
  assign array_update_71770[4] = add_71711 == 32'h0000_0004 ? array_update_71768 : array_update_71760[4];
  assign array_update_71770[5] = add_71711 == 32'h0000_0005 ? array_update_71768 : array_update_71760[5];
  assign array_update_71770[6] = add_71711 == 32'h0000_0006 ? array_update_71768 : array_update_71760[6];
  assign array_update_71770[7] = add_71711 == 32'h0000_0007 ? array_update_71768 : array_update_71760[7];
  assign array_update_71770[8] = add_71711 == 32'h0000_0008 ? array_update_71768 : array_update_71760[8];
  assign array_update_71770[9] = add_71711 == 32'h0000_0009 ? array_update_71768 : array_update_71760[9];
  assign array_update_71772[0] = add_71713 == 32'h0000_0000 ? array_update_71769 : array_update_71762[0];
  assign array_update_71772[1] = add_71713 == 32'h0000_0001 ? array_update_71769 : array_update_71762[1];
  assign array_update_71772[2] = add_71713 == 32'h0000_0002 ? array_update_71769 : array_update_71762[2];
  assign array_update_71772[3] = add_71713 == 32'h0000_0003 ? array_update_71769 : array_update_71762[3];
  assign array_update_71772[4] = add_71713 == 32'h0000_0004 ? array_update_71769 : array_update_71762[4];
  assign array_update_71772[5] = add_71713 == 32'h0000_0005 ? array_update_71769 : array_update_71762[5];
  assign array_update_71772[6] = add_71713 == 32'h0000_0006 ? array_update_71769 : array_update_71762[6];
  assign array_update_71772[7] = add_71713 == 32'h0000_0007 ? array_update_71769 : array_update_71762[7];
  assign array_update_71772[8] = add_71713 == 32'h0000_0008 ? array_update_71769 : array_update_71762[8];
  assign array_update_71772[9] = add_71713 == 32'h0000_0009 ? array_update_71769 : array_update_71762[9];
  assign array_index_71774 = array_update_71770[add_71711 > 32'h0000_0009 ? 4'h9 : add_71711[3:0]];
  assign add_71775 = add_71765 + 32'h0000_0001;
  assign array_index_71776 = array_update_71772[add_71713 > 32'h0000_0009 ? 4'h9 : add_71713[3:0]];
  assign add_71777 = add_71767 + 32'h0000_0001;
  assign array_update_71778[0] = add_71775 == 32'h0000_0000 ? TestBlock__A_op76 : array_index_71774[0];
  assign array_update_71778[1] = add_71775 == 32'h0000_0001 ? TestBlock__A_op76 : array_index_71774[1];
  assign array_update_71778[2] = add_71775 == 32'h0000_0002 ? TestBlock__A_op76 : array_index_71774[2];
  assign array_update_71778[3] = add_71775 == 32'h0000_0003 ? TestBlock__A_op76 : array_index_71774[3];
  assign array_update_71778[4] = add_71775 == 32'h0000_0004 ? TestBlock__A_op76 : array_index_71774[4];
  assign array_update_71778[5] = add_71775 == 32'h0000_0005 ? TestBlock__A_op76 : array_index_71774[5];
  assign array_update_71778[6] = add_71775 == 32'h0000_0006 ? TestBlock__A_op76 : array_index_71774[6];
  assign array_update_71778[7] = add_71775 == 32'h0000_0007 ? TestBlock__A_op76 : array_index_71774[7];
  assign array_update_71778[8] = add_71775 == 32'h0000_0008 ? TestBlock__A_op76 : array_index_71774[8];
  assign array_update_71778[9] = add_71775 == 32'h0000_0009 ? TestBlock__A_op76 : array_index_71774[9];
  assign array_update_71779[0] = add_71777 == 32'h0000_0000 ? TestBlock__B_op76 : array_index_71776[0];
  assign array_update_71779[1] = add_71777 == 32'h0000_0001 ? TestBlock__B_op76 : array_index_71776[1];
  assign array_update_71779[2] = add_71777 == 32'h0000_0002 ? TestBlock__B_op76 : array_index_71776[2];
  assign array_update_71779[3] = add_71777 == 32'h0000_0003 ? TestBlock__B_op76 : array_index_71776[3];
  assign array_update_71779[4] = add_71777 == 32'h0000_0004 ? TestBlock__B_op76 : array_index_71776[4];
  assign array_update_71779[5] = add_71777 == 32'h0000_0005 ? TestBlock__B_op76 : array_index_71776[5];
  assign array_update_71779[6] = add_71777 == 32'h0000_0006 ? TestBlock__B_op76 : array_index_71776[6];
  assign array_update_71779[7] = add_71777 == 32'h0000_0007 ? TestBlock__B_op76 : array_index_71776[7];
  assign array_update_71779[8] = add_71777 == 32'h0000_0008 ? TestBlock__B_op76 : array_index_71776[8];
  assign array_update_71779[9] = add_71777 == 32'h0000_0009 ? TestBlock__B_op76 : array_index_71776[9];
  assign array_update_71780[0] = add_71711 == 32'h0000_0000 ? array_update_71778 : array_update_71770[0];
  assign array_update_71780[1] = add_71711 == 32'h0000_0001 ? array_update_71778 : array_update_71770[1];
  assign array_update_71780[2] = add_71711 == 32'h0000_0002 ? array_update_71778 : array_update_71770[2];
  assign array_update_71780[3] = add_71711 == 32'h0000_0003 ? array_update_71778 : array_update_71770[3];
  assign array_update_71780[4] = add_71711 == 32'h0000_0004 ? array_update_71778 : array_update_71770[4];
  assign array_update_71780[5] = add_71711 == 32'h0000_0005 ? array_update_71778 : array_update_71770[5];
  assign array_update_71780[6] = add_71711 == 32'h0000_0006 ? array_update_71778 : array_update_71770[6];
  assign array_update_71780[7] = add_71711 == 32'h0000_0007 ? array_update_71778 : array_update_71770[7];
  assign array_update_71780[8] = add_71711 == 32'h0000_0008 ? array_update_71778 : array_update_71770[8];
  assign array_update_71780[9] = add_71711 == 32'h0000_0009 ? array_update_71778 : array_update_71770[9];
  assign array_update_71782[0] = add_71713 == 32'h0000_0000 ? array_update_71779 : array_update_71772[0];
  assign array_update_71782[1] = add_71713 == 32'h0000_0001 ? array_update_71779 : array_update_71772[1];
  assign array_update_71782[2] = add_71713 == 32'h0000_0002 ? array_update_71779 : array_update_71772[2];
  assign array_update_71782[3] = add_71713 == 32'h0000_0003 ? array_update_71779 : array_update_71772[3];
  assign array_update_71782[4] = add_71713 == 32'h0000_0004 ? array_update_71779 : array_update_71772[4];
  assign array_update_71782[5] = add_71713 == 32'h0000_0005 ? array_update_71779 : array_update_71772[5];
  assign array_update_71782[6] = add_71713 == 32'h0000_0006 ? array_update_71779 : array_update_71772[6];
  assign array_update_71782[7] = add_71713 == 32'h0000_0007 ? array_update_71779 : array_update_71772[7];
  assign array_update_71782[8] = add_71713 == 32'h0000_0008 ? array_update_71779 : array_update_71772[8];
  assign array_update_71782[9] = add_71713 == 32'h0000_0009 ? array_update_71779 : array_update_71772[9];
  assign array_index_71784 = array_update_71780[add_71711 > 32'h0000_0009 ? 4'h9 : add_71711[3:0]];
  assign add_71785 = add_71775 + 32'h0000_0001;
  assign array_index_71786 = array_update_71782[add_71713 > 32'h0000_0009 ? 4'h9 : add_71713[3:0]];
  assign add_71787 = add_71777 + 32'h0000_0001;
  assign array_update_71788[0] = add_71785 == 32'h0000_0000 ? TestBlock__A_op77 : array_index_71784[0];
  assign array_update_71788[1] = add_71785 == 32'h0000_0001 ? TestBlock__A_op77 : array_index_71784[1];
  assign array_update_71788[2] = add_71785 == 32'h0000_0002 ? TestBlock__A_op77 : array_index_71784[2];
  assign array_update_71788[3] = add_71785 == 32'h0000_0003 ? TestBlock__A_op77 : array_index_71784[3];
  assign array_update_71788[4] = add_71785 == 32'h0000_0004 ? TestBlock__A_op77 : array_index_71784[4];
  assign array_update_71788[5] = add_71785 == 32'h0000_0005 ? TestBlock__A_op77 : array_index_71784[5];
  assign array_update_71788[6] = add_71785 == 32'h0000_0006 ? TestBlock__A_op77 : array_index_71784[6];
  assign array_update_71788[7] = add_71785 == 32'h0000_0007 ? TestBlock__A_op77 : array_index_71784[7];
  assign array_update_71788[8] = add_71785 == 32'h0000_0008 ? TestBlock__A_op77 : array_index_71784[8];
  assign array_update_71788[9] = add_71785 == 32'h0000_0009 ? TestBlock__A_op77 : array_index_71784[9];
  assign array_update_71789[0] = add_71787 == 32'h0000_0000 ? TestBlock__B_op77 : array_index_71786[0];
  assign array_update_71789[1] = add_71787 == 32'h0000_0001 ? TestBlock__B_op77 : array_index_71786[1];
  assign array_update_71789[2] = add_71787 == 32'h0000_0002 ? TestBlock__B_op77 : array_index_71786[2];
  assign array_update_71789[3] = add_71787 == 32'h0000_0003 ? TestBlock__B_op77 : array_index_71786[3];
  assign array_update_71789[4] = add_71787 == 32'h0000_0004 ? TestBlock__B_op77 : array_index_71786[4];
  assign array_update_71789[5] = add_71787 == 32'h0000_0005 ? TestBlock__B_op77 : array_index_71786[5];
  assign array_update_71789[6] = add_71787 == 32'h0000_0006 ? TestBlock__B_op77 : array_index_71786[6];
  assign array_update_71789[7] = add_71787 == 32'h0000_0007 ? TestBlock__B_op77 : array_index_71786[7];
  assign array_update_71789[8] = add_71787 == 32'h0000_0008 ? TestBlock__B_op77 : array_index_71786[8];
  assign array_update_71789[9] = add_71787 == 32'h0000_0009 ? TestBlock__B_op77 : array_index_71786[9];
  assign array_update_71790[0] = add_71711 == 32'h0000_0000 ? array_update_71788 : array_update_71780[0];
  assign array_update_71790[1] = add_71711 == 32'h0000_0001 ? array_update_71788 : array_update_71780[1];
  assign array_update_71790[2] = add_71711 == 32'h0000_0002 ? array_update_71788 : array_update_71780[2];
  assign array_update_71790[3] = add_71711 == 32'h0000_0003 ? array_update_71788 : array_update_71780[3];
  assign array_update_71790[4] = add_71711 == 32'h0000_0004 ? array_update_71788 : array_update_71780[4];
  assign array_update_71790[5] = add_71711 == 32'h0000_0005 ? array_update_71788 : array_update_71780[5];
  assign array_update_71790[6] = add_71711 == 32'h0000_0006 ? array_update_71788 : array_update_71780[6];
  assign array_update_71790[7] = add_71711 == 32'h0000_0007 ? array_update_71788 : array_update_71780[7];
  assign array_update_71790[8] = add_71711 == 32'h0000_0008 ? array_update_71788 : array_update_71780[8];
  assign array_update_71790[9] = add_71711 == 32'h0000_0009 ? array_update_71788 : array_update_71780[9];
  assign array_update_71792[0] = add_71713 == 32'h0000_0000 ? array_update_71789 : array_update_71782[0];
  assign array_update_71792[1] = add_71713 == 32'h0000_0001 ? array_update_71789 : array_update_71782[1];
  assign array_update_71792[2] = add_71713 == 32'h0000_0002 ? array_update_71789 : array_update_71782[2];
  assign array_update_71792[3] = add_71713 == 32'h0000_0003 ? array_update_71789 : array_update_71782[3];
  assign array_update_71792[4] = add_71713 == 32'h0000_0004 ? array_update_71789 : array_update_71782[4];
  assign array_update_71792[5] = add_71713 == 32'h0000_0005 ? array_update_71789 : array_update_71782[5];
  assign array_update_71792[6] = add_71713 == 32'h0000_0006 ? array_update_71789 : array_update_71782[6];
  assign array_update_71792[7] = add_71713 == 32'h0000_0007 ? array_update_71789 : array_update_71782[7];
  assign array_update_71792[8] = add_71713 == 32'h0000_0008 ? array_update_71789 : array_update_71782[8];
  assign array_update_71792[9] = add_71713 == 32'h0000_0009 ? array_update_71789 : array_update_71782[9];
  assign array_index_71794 = array_update_71790[add_71711 > 32'h0000_0009 ? 4'h9 : add_71711[3:0]];
  assign add_71795 = add_71785 + 32'h0000_0001;
  assign array_index_71796 = array_update_71792[add_71713 > 32'h0000_0009 ? 4'h9 : add_71713[3:0]];
  assign add_71797 = add_71787 + 32'h0000_0001;
  assign array_update_71798[0] = add_71795 == 32'h0000_0000 ? TestBlock__A_op78 : array_index_71794[0];
  assign array_update_71798[1] = add_71795 == 32'h0000_0001 ? TestBlock__A_op78 : array_index_71794[1];
  assign array_update_71798[2] = add_71795 == 32'h0000_0002 ? TestBlock__A_op78 : array_index_71794[2];
  assign array_update_71798[3] = add_71795 == 32'h0000_0003 ? TestBlock__A_op78 : array_index_71794[3];
  assign array_update_71798[4] = add_71795 == 32'h0000_0004 ? TestBlock__A_op78 : array_index_71794[4];
  assign array_update_71798[5] = add_71795 == 32'h0000_0005 ? TestBlock__A_op78 : array_index_71794[5];
  assign array_update_71798[6] = add_71795 == 32'h0000_0006 ? TestBlock__A_op78 : array_index_71794[6];
  assign array_update_71798[7] = add_71795 == 32'h0000_0007 ? TestBlock__A_op78 : array_index_71794[7];
  assign array_update_71798[8] = add_71795 == 32'h0000_0008 ? TestBlock__A_op78 : array_index_71794[8];
  assign array_update_71798[9] = add_71795 == 32'h0000_0009 ? TestBlock__A_op78 : array_index_71794[9];
  assign array_update_71799[0] = add_71797 == 32'h0000_0000 ? TestBlock__B_op78 : array_index_71796[0];
  assign array_update_71799[1] = add_71797 == 32'h0000_0001 ? TestBlock__B_op78 : array_index_71796[1];
  assign array_update_71799[2] = add_71797 == 32'h0000_0002 ? TestBlock__B_op78 : array_index_71796[2];
  assign array_update_71799[3] = add_71797 == 32'h0000_0003 ? TestBlock__B_op78 : array_index_71796[3];
  assign array_update_71799[4] = add_71797 == 32'h0000_0004 ? TestBlock__B_op78 : array_index_71796[4];
  assign array_update_71799[5] = add_71797 == 32'h0000_0005 ? TestBlock__B_op78 : array_index_71796[5];
  assign array_update_71799[6] = add_71797 == 32'h0000_0006 ? TestBlock__B_op78 : array_index_71796[6];
  assign array_update_71799[7] = add_71797 == 32'h0000_0007 ? TestBlock__B_op78 : array_index_71796[7];
  assign array_update_71799[8] = add_71797 == 32'h0000_0008 ? TestBlock__B_op78 : array_index_71796[8];
  assign array_update_71799[9] = add_71797 == 32'h0000_0009 ? TestBlock__B_op78 : array_index_71796[9];
  assign array_update_71800[0] = add_71711 == 32'h0000_0000 ? array_update_71798 : array_update_71790[0];
  assign array_update_71800[1] = add_71711 == 32'h0000_0001 ? array_update_71798 : array_update_71790[1];
  assign array_update_71800[2] = add_71711 == 32'h0000_0002 ? array_update_71798 : array_update_71790[2];
  assign array_update_71800[3] = add_71711 == 32'h0000_0003 ? array_update_71798 : array_update_71790[3];
  assign array_update_71800[4] = add_71711 == 32'h0000_0004 ? array_update_71798 : array_update_71790[4];
  assign array_update_71800[5] = add_71711 == 32'h0000_0005 ? array_update_71798 : array_update_71790[5];
  assign array_update_71800[6] = add_71711 == 32'h0000_0006 ? array_update_71798 : array_update_71790[6];
  assign array_update_71800[7] = add_71711 == 32'h0000_0007 ? array_update_71798 : array_update_71790[7];
  assign array_update_71800[8] = add_71711 == 32'h0000_0008 ? array_update_71798 : array_update_71790[8];
  assign array_update_71800[9] = add_71711 == 32'h0000_0009 ? array_update_71798 : array_update_71790[9];
  assign array_update_71802[0] = add_71713 == 32'h0000_0000 ? array_update_71799 : array_update_71792[0];
  assign array_update_71802[1] = add_71713 == 32'h0000_0001 ? array_update_71799 : array_update_71792[1];
  assign array_update_71802[2] = add_71713 == 32'h0000_0002 ? array_update_71799 : array_update_71792[2];
  assign array_update_71802[3] = add_71713 == 32'h0000_0003 ? array_update_71799 : array_update_71792[3];
  assign array_update_71802[4] = add_71713 == 32'h0000_0004 ? array_update_71799 : array_update_71792[4];
  assign array_update_71802[5] = add_71713 == 32'h0000_0005 ? array_update_71799 : array_update_71792[5];
  assign array_update_71802[6] = add_71713 == 32'h0000_0006 ? array_update_71799 : array_update_71792[6];
  assign array_update_71802[7] = add_71713 == 32'h0000_0007 ? array_update_71799 : array_update_71792[7];
  assign array_update_71802[8] = add_71713 == 32'h0000_0008 ? array_update_71799 : array_update_71792[8];
  assign array_update_71802[9] = add_71713 == 32'h0000_0009 ? array_update_71799 : array_update_71792[9];
  assign array_index_71804 = array_update_71800[add_71711 > 32'h0000_0009 ? 4'h9 : add_71711[3:0]];
  assign add_71805 = add_71795 + 32'h0000_0001;
  assign array_index_71806 = array_update_71802[add_71713 > 32'h0000_0009 ? 4'h9 : add_71713[3:0]];
  assign add_71807 = add_71797 + 32'h0000_0001;
  assign array_update_71808[0] = add_71805 == 32'h0000_0000 ? TestBlock__A_op79 : array_index_71804[0];
  assign array_update_71808[1] = add_71805 == 32'h0000_0001 ? TestBlock__A_op79 : array_index_71804[1];
  assign array_update_71808[2] = add_71805 == 32'h0000_0002 ? TestBlock__A_op79 : array_index_71804[2];
  assign array_update_71808[3] = add_71805 == 32'h0000_0003 ? TestBlock__A_op79 : array_index_71804[3];
  assign array_update_71808[4] = add_71805 == 32'h0000_0004 ? TestBlock__A_op79 : array_index_71804[4];
  assign array_update_71808[5] = add_71805 == 32'h0000_0005 ? TestBlock__A_op79 : array_index_71804[5];
  assign array_update_71808[6] = add_71805 == 32'h0000_0006 ? TestBlock__A_op79 : array_index_71804[6];
  assign array_update_71808[7] = add_71805 == 32'h0000_0007 ? TestBlock__A_op79 : array_index_71804[7];
  assign array_update_71808[8] = add_71805 == 32'h0000_0008 ? TestBlock__A_op79 : array_index_71804[8];
  assign array_update_71808[9] = add_71805 == 32'h0000_0009 ? TestBlock__A_op79 : array_index_71804[9];
  assign array_update_71810[0] = add_71807 == 32'h0000_0000 ? TestBlock__B_op79 : array_index_71806[0];
  assign array_update_71810[1] = add_71807 == 32'h0000_0001 ? TestBlock__B_op79 : array_index_71806[1];
  assign array_update_71810[2] = add_71807 == 32'h0000_0002 ? TestBlock__B_op79 : array_index_71806[2];
  assign array_update_71810[3] = add_71807 == 32'h0000_0003 ? TestBlock__B_op79 : array_index_71806[3];
  assign array_update_71810[4] = add_71807 == 32'h0000_0004 ? TestBlock__B_op79 : array_index_71806[4];
  assign array_update_71810[5] = add_71807 == 32'h0000_0005 ? TestBlock__B_op79 : array_index_71806[5];
  assign array_update_71810[6] = add_71807 == 32'h0000_0006 ? TestBlock__B_op79 : array_index_71806[6];
  assign array_update_71810[7] = add_71807 == 32'h0000_0007 ? TestBlock__B_op79 : array_index_71806[7];
  assign array_update_71810[8] = add_71807 == 32'h0000_0008 ? TestBlock__B_op79 : array_index_71806[8];
  assign array_update_71810[9] = add_71807 == 32'h0000_0009 ? TestBlock__B_op79 : array_index_71806[9];
  assign array_update_71812[0] = add_71711 == 32'h0000_0000 ? array_update_71808 : array_update_71800[0];
  assign array_update_71812[1] = add_71711 == 32'h0000_0001 ? array_update_71808 : array_update_71800[1];
  assign array_update_71812[2] = add_71711 == 32'h0000_0002 ? array_update_71808 : array_update_71800[2];
  assign array_update_71812[3] = add_71711 == 32'h0000_0003 ? array_update_71808 : array_update_71800[3];
  assign array_update_71812[4] = add_71711 == 32'h0000_0004 ? array_update_71808 : array_update_71800[4];
  assign array_update_71812[5] = add_71711 == 32'h0000_0005 ? array_update_71808 : array_update_71800[5];
  assign array_update_71812[6] = add_71711 == 32'h0000_0006 ? array_update_71808 : array_update_71800[6];
  assign array_update_71812[7] = add_71711 == 32'h0000_0007 ? array_update_71808 : array_update_71800[7];
  assign array_update_71812[8] = add_71711 == 32'h0000_0008 ? array_update_71808 : array_update_71800[8];
  assign array_update_71812[9] = add_71711 == 32'h0000_0009 ? array_update_71808 : array_update_71800[9];
  assign add_71813 = add_71711 + 32'h0000_0001;
  assign array_update_71814[0] = add_71713 == 32'h0000_0000 ? array_update_71810 : array_update_71802[0];
  assign array_update_71814[1] = add_71713 == 32'h0000_0001 ? array_update_71810 : array_update_71802[1];
  assign array_update_71814[2] = add_71713 == 32'h0000_0002 ? array_update_71810 : array_update_71802[2];
  assign array_update_71814[3] = add_71713 == 32'h0000_0003 ? array_update_71810 : array_update_71802[3];
  assign array_update_71814[4] = add_71713 == 32'h0000_0004 ? array_update_71810 : array_update_71802[4];
  assign array_update_71814[5] = add_71713 == 32'h0000_0005 ? array_update_71810 : array_update_71802[5];
  assign array_update_71814[6] = add_71713 == 32'h0000_0006 ? array_update_71810 : array_update_71802[6];
  assign array_update_71814[7] = add_71713 == 32'h0000_0007 ? array_update_71810 : array_update_71802[7];
  assign array_update_71814[8] = add_71713 == 32'h0000_0008 ? array_update_71810 : array_update_71802[8];
  assign array_update_71814[9] = add_71713 == 32'h0000_0009 ? array_update_71810 : array_update_71802[9];
  assign add_71815 = add_71713 + 32'h0000_0001;
  assign array_index_71816 = array_update_71812[add_71813 > 32'h0000_0009 ? 4'h9 : add_71813[3:0]];
  assign literal_71817 = 32'h0000_0000;
  assign array_index_71818 = array_update_71814[add_71815 > 32'h0000_0009 ? 4'h9 : add_71815[3:0]];
  assign literal_71819 = 32'h0000_0000;
  assign array_update_71820[0] = literal_71817 == 32'h0000_0000 ? TestBlock__A_op80 : array_index_71816[0];
  assign array_update_71820[1] = literal_71817 == 32'h0000_0001 ? TestBlock__A_op80 : array_index_71816[1];
  assign array_update_71820[2] = literal_71817 == 32'h0000_0002 ? TestBlock__A_op80 : array_index_71816[2];
  assign array_update_71820[3] = literal_71817 == 32'h0000_0003 ? TestBlock__A_op80 : array_index_71816[3];
  assign array_update_71820[4] = literal_71817 == 32'h0000_0004 ? TestBlock__A_op80 : array_index_71816[4];
  assign array_update_71820[5] = literal_71817 == 32'h0000_0005 ? TestBlock__A_op80 : array_index_71816[5];
  assign array_update_71820[6] = literal_71817 == 32'h0000_0006 ? TestBlock__A_op80 : array_index_71816[6];
  assign array_update_71820[7] = literal_71817 == 32'h0000_0007 ? TestBlock__A_op80 : array_index_71816[7];
  assign array_update_71820[8] = literal_71817 == 32'h0000_0008 ? TestBlock__A_op80 : array_index_71816[8];
  assign array_update_71820[9] = literal_71817 == 32'h0000_0009 ? TestBlock__A_op80 : array_index_71816[9];
  assign array_update_71821[0] = literal_71819 == 32'h0000_0000 ? TestBlock__B_op80 : array_index_71818[0];
  assign array_update_71821[1] = literal_71819 == 32'h0000_0001 ? TestBlock__B_op80 : array_index_71818[1];
  assign array_update_71821[2] = literal_71819 == 32'h0000_0002 ? TestBlock__B_op80 : array_index_71818[2];
  assign array_update_71821[3] = literal_71819 == 32'h0000_0003 ? TestBlock__B_op80 : array_index_71818[3];
  assign array_update_71821[4] = literal_71819 == 32'h0000_0004 ? TestBlock__B_op80 : array_index_71818[4];
  assign array_update_71821[5] = literal_71819 == 32'h0000_0005 ? TestBlock__B_op80 : array_index_71818[5];
  assign array_update_71821[6] = literal_71819 == 32'h0000_0006 ? TestBlock__B_op80 : array_index_71818[6];
  assign array_update_71821[7] = literal_71819 == 32'h0000_0007 ? TestBlock__B_op80 : array_index_71818[7];
  assign array_update_71821[8] = literal_71819 == 32'h0000_0008 ? TestBlock__B_op80 : array_index_71818[8];
  assign array_update_71821[9] = literal_71819 == 32'h0000_0009 ? TestBlock__B_op80 : array_index_71818[9];
  assign array_update_71822[0] = add_71813 == 32'h0000_0000 ? array_update_71820 : array_update_71812[0];
  assign array_update_71822[1] = add_71813 == 32'h0000_0001 ? array_update_71820 : array_update_71812[1];
  assign array_update_71822[2] = add_71813 == 32'h0000_0002 ? array_update_71820 : array_update_71812[2];
  assign array_update_71822[3] = add_71813 == 32'h0000_0003 ? array_update_71820 : array_update_71812[3];
  assign array_update_71822[4] = add_71813 == 32'h0000_0004 ? array_update_71820 : array_update_71812[4];
  assign array_update_71822[5] = add_71813 == 32'h0000_0005 ? array_update_71820 : array_update_71812[5];
  assign array_update_71822[6] = add_71813 == 32'h0000_0006 ? array_update_71820 : array_update_71812[6];
  assign array_update_71822[7] = add_71813 == 32'h0000_0007 ? array_update_71820 : array_update_71812[7];
  assign array_update_71822[8] = add_71813 == 32'h0000_0008 ? array_update_71820 : array_update_71812[8];
  assign array_update_71822[9] = add_71813 == 32'h0000_0009 ? array_update_71820 : array_update_71812[9];
  assign array_update_71824[0] = add_71815 == 32'h0000_0000 ? array_update_71821 : array_update_71814[0];
  assign array_update_71824[1] = add_71815 == 32'h0000_0001 ? array_update_71821 : array_update_71814[1];
  assign array_update_71824[2] = add_71815 == 32'h0000_0002 ? array_update_71821 : array_update_71814[2];
  assign array_update_71824[3] = add_71815 == 32'h0000_0003 ? array_update_71821 : array_update_71814[3];
  assign array_update_71824[4] = add_71815 == 32'h0000_0004 ? array_update_71821 : array_update_71814[4];
  assign array_update_71824[5] = add_71815 == 32'h0000_0005 ? array_update_71821 : array_update_71814[5];
  assign array_update_71824[6] = add_71815 == 32'h0000_0006 ? array_update_71821 : array_update_71814[6];
  assign array_update_71824[7] = add_71815 == 32'h0000_0007 ? array_update_71821 : array_update_71814[7];
  assign array_update_71824[8] = add_71815 == 32'h0000_0008 ? array_update_71821 : array_update_71814[8];
  assign array_update_71824[9] = add_71815 == 32'h0000_0009 ? array_update_71821 : array_update_71814[9];
  assign array_index_71826 = array_update_71822[add_71813 > 32'h0000_0009 ? 4'h9 : add_71813[3:0]];
  assign add_71827 = literal_71817 + 32'h0000_0001;
  assign array_index_71828 = array_update_71824[add_71815 > 32'h0000_0009 ? 4'h9 : add_71815[3:0]];
  assign add_71829 = literal_71819 + 32'h0000_0001;
  assign array_update_71830[0] = add_71827 == 32'h0000_0000 ? TestBlock__A_op81 : array_index_71826[0];
  assign array_update_71830[1] = add_71827 == 32'h0000_0001 ? TestBlock__A_op81 : array_index_71826[1];
  assign array_update_71830[2] = add_71827 == 32'h0000_0002 ? TestBlock__A_op81 : array_index_71826[2];
  assign array_update_71830[3] = add_71827 == 32'h0000_0003 ? TestBlock__A_op81 : array_index_71826[3];
  assign array_update_71830[4] = add_71827 == 32'h0000_0004 ? TestBlock__A_op81 : array_index_71826[4];
  assign array_update_71830[5] = add_71827 == 32'h0000_0005 ? TestBlock__A_op81 : array_index_71826[5];
  assign array_update_71830[6] = add_71827 == 32'h0000_0006 ? TestBlock__A_op81 : array_index_71826[6];
  assign array_update_71830[7] = add_71827 == 32'h0000_0007 ? TestBlock__A_op81 : array_index_71826[7];
  assign array_update_71830[8] = add_71827 == 32'h0000_0008 ? TestBlock__A_op81 : array_index_71826[8];
  assign array_update_71830[9] = add_71827 == 32'h0000_0009 ? TestBlock__A_op81 : array_index_71826[9];
  assign array_update_71831[0] = add_71829 == 32'h0000_0000 ? TestBlock__B_op81 : array_index_71828[0];
  assign array_update_71831[1] = add_71829 == 32'h0000_0001 ? TestBlock__B_op81 : array_index_71828[1];
  assign array_update_71831[2] = add_71829 == 32'h0000_0002 ? TestBlock__B_op81 : array_index_71828[2];
  assign array_update_71831[3] = add_71829 == 32'h0000_0003 ? TestBlock__B_op81 : array_index_71828[3];
  assign array_update_71831[4] = add_71829 == 32'h0000_0004 ? TestBlock__B_op81 : array_index_71828[4];
  assign array_update_71831[5] = add_71829 == 32'h0000_0005 ? TestBlock__B_op81 : array_index_71828[5];
  assign array_update_71831[6] = add_71829 == 32'h0000_0006 ? TestBlock__B_op81 : array_index_71828[6];
  assign array_update_71831[7] = add_71829 == 32'h0000_0007 ? TestBlock__B_op81 : array_index_71828[7];
  assign array_update_71831[8] = add_71829 == 32'h0000_0008 ? TestBlock__B_op81 : array_index_71828[8];
  assign array_update_71831[9] = add_71829 == 32'h0000_0009 ? TestBlock__B_op81 : array_index_71828[9];
  assign array_update_71832[0] = add_71813 == 32'h0000_0000 ? array_update_71830 : array_update_71822[0];
  assign array_update_71832[1] = add_71813 == 32'h0000_0001 ? array_update_71830 : array_update_71822[1];
  assign array_update_71832[2] = add_71813 == 32'h0000_0002 ? array_update_71830 : array_update_71822[2];
  assign array_update_71832[3] = add_71813 == 32'h0000_0003 ? array_update_71830 : array_update_71822[3];
  assign array_update_71832[4] = add_71813 == 32'h0000_0004 ? array_update_71830 : array_update_71822[4];
  assign array_update_71832[5] = add_71813 == 32'h0000_0005 ? array_update_71830 : array_update_71822[5];
  assign array_update_71832[6] = add_71813 == 32'h0000_0006 ? array_update_71830 : array_update_71822[6];
  assign array_update_71832[7] = add_71813 == 32'h0000_0007 ? array_update_71830 : array_update_71822[7];
  assign array_update_71832[8] = add_71813 == 32'h0000_0008 ? array_update_71830 : array_update_71822[8];
  assign array_update_71832[9] = add_71813 == 32'h0000_0009 ? array_update_71830 : array_update_71822[9];
  assign array_update_71834[0] = add_71815 == 32'h0000_0000 ? array_update_71831 : array_update_71824[0];
  assign array_update_71834[1] = add_71815 == 32'h0000_0001 ? array_update_71831 : array_update_71824[1];
  assign array_update_71834[2] = add_71815 == 32'h0000_0002 ? array_update_71831 : array_update_71824[2];
  assign array_update_71834[3] = add_71815 == 32'h0000_0003 ? array_update_71831 : array_update_71824[3];
  assign array_update_71834[4] = add_71815 == 32'h0000_0004 ? array_update_71831 : array_update_71824[4];
  assign array_update_71834[5] = add_71815 == 32'h0000_0005 ? array_update_71831 : array_update_71824[5];
  assign array_update_71834[6] = add_71815 == 32'h0000_0006 ? array_update_71831 : array_update_71824[6];
  assign array_update_71834[7] = add_71815 == 32'h0000_0007 ? array_update_71831 : array_update_71824[7];
  assign array_update_71834[8] = add_71815 == 32'h0000_0008 ? array_update_71831 : array_update_71824[8];
  assign array_update_71834[9] = add_71815 == 32'h0000_0009 ? array_update_71831 : array_update_71824[9];
  assign array_index_71836 = array_update_71832[add_71813 > 32'h0000_0009 ? 4'h9 : add_71813[3:0]];
  assign add_71837 = add_71827 + 32'h0000_0001;
  assign array_index_71838 = array_update_71834[add_71815 > 32'h0000_0009 ? 4'h9 : add_71815[3:0]];
  assign add_71839 = add_71829 + 32'h0000_0001;
  assign array_update_71840[0] = add_71837 == 32'h0000_0000 ? TestBlock__A_op82 : array_index_71836[0];
  assign array_update_71840[1] = add_71837 == 32'h0000_0001 ? TestBlock__A_op82 : array_index_71836[1];
  assign array_update_71840[2] = add_71837 == 32'h0000_0002 ? TestBlock__A_op82 : array_index_71836[2];
  assign array_update_71840[3] = add_71837 == 32'h0000_0003 ? TestBlock__A_op82 : array_index_71836[3];
  assign array_update_71840[4] = add_71837 == 32'h0000_0004 ? TestBlock__A_op82 : array_index_71836[4];
  assign array_update_71840[5] = add_71837 == 32'h0000_0005 ? TestBlock__A_op82 : array_index_71836[5];
  assign array_update_71840[6] = add_71837 == 32'h0000_0006 ? TestBlock__A_op82 : array_index_71836[6];
  assign array_update_71840[7] = add_71837 == 32'h0000_0007 ? TestBlock__A_op82 : array_index_71836[7];
  assign array_update_71840[8] = add_71837 == 32'h0000_0008 ? TestBlock__A_op82 : array_index_71836[8];
  assign array_update_71840[9] = add_71837 == 32'h0000_0009 ? TestBlock__A_op82 : array_index_71836[9];
  assign array_update_71841[0] = add_71839 == 32'h0000_0000 ? TestBlock__B_op82 : array_index_71838[0];
  assign array_update_71841[1] = add_71839 == 32'h0000_0001 ? TestBlock__B_op82 : array_index_71838[1];
  assign array_update_71841[2] = add_71839 == 32'h0000_0002 ? TestBlock__B_op82 : array_index_71838[2];
  assign array_update_71841[3] = add_71839 == 32'h0000_0003 ? TestBlock__B_op82 : array_index_71838[3];
  assign array_update_71841[4] = add_71839 == 32'h0000_0004 ? TestBlock__B_op82 : array_index_71838[4];
  assign array_update_71841[5] = add_71839 == 32'h0000_0005 ? TestBlock__B_op82 : array_index_71838[5];
  assign array_update_71841[6] = add_71839 == 32'h0000_0006 ? TestBlock__B_op82 : array_index_71838[6];
  assign array_update_71841[7] = add_71839 == 32'h0000_0007 ? TestBlock__B_op82 : array_index_71838[7];
  assign array_update_71841[8] = add_71839 == 32'h0000_0008 ? TestBlock__B_op82 : array_index_71838[8];
  assign array_update_71841[9] = add_71839 == 32'h0000_0009 ? TestBlock__B_op82 : array_index_71838[9];
  assign array_update_71842[0] = add_71813 == 32'h0000_0000 ? array_update_71840 : array_update_71832[0];
  assign array_update_71842[1] = add_71813 == 32'h0000_0001 ? array_update_71840 : array_update_71832[1];
  assign array_update_71842[2] = add_71813 == 32'h0000_0002 ? array_update_71840 : array_update_71832[2];
  assign array_update_71842[3] = add_71813 == 32'h0000_0003 ? array_update_71840 : array_update_71832[3];
  assign array_update_71842[4] = add_71813 == 32'h0000_0004 ? array_update_71840 : array_update_71832[4];
  assign array_update_71842[5] = add_71813 == 32'h0000_0005 ? array_update_71840 : array_update_71832[5];
  assign array_update_71842[6] = add_71813 == 32'h0000_0006 ? array_update_71840 : array_update_71832[6];
  assign array_update_71842[7] = add_71813 == 32'h0000_0007 ? array_update_71840 : array_update_71832[7];
  assign array_update_71842[8] = add_71813 == 32'h0000_0008 ? array_update_71840 : array_update_71832[8];
  assign array_update_71842[9] = add_71813 == 32'h0000_0009 ? array_update_71840 : array_update_71832[9];
  assign array_update_71844[0] = add_71815 == 32'h0000_0000 ? array_update_71841 : array_update_71834[0];
  assign array_update_71844[1] = add_71815 == 32'h0000_0001 ? array_update_71841 : array_update_71834[1];
  assign array_update_71844[2] = add_71815 == 32'h0000_0002 ? array_update_71841 : array_update_71834[2];
  assign array_update_71844[3] = add_71815 == 32'h0000_0003 ? array_update_71841 : array_update_71834[3];
  assign array_update_71844[4] = add_71815 == 32'h0000_0004 ? array_update_71841 : array_update_71834[4];
  assign array_update_71844[5] = add_71815 == 32'h0000_0005 ? array_update_71841 : array_update_71834[5];
  assign array_update_71844[6] = add_71815 == 32'h0000_0006 ? array_update_71841 : array_update_71834[6];
  assign array_update_71844[7] = add_71815 == 32'h0000_0007 ? array_update_71841 : array_update_71834[7];
  assign array_update_71844[8] = add_71815 == 32'h0000_0008 ? array_update_71841 : array_update_71834[8];
  assign array_update_71844[9] = add_71815 == 32'h0000_0009 ? array_update_71841 : array_update_71834[9];
  assign array_index_71846 = array_update_71842[add_71813 > 32'h0000_0009 ? 4'h9 : add_71813[3:0]];
  assign add_71847 = add_71837 + 32'h0000_0001;
  assign array_index_71848 = array_update_71844[add_71815 > 32'h0000_0009 ? 4'h9 : add_71815[3:0]];
  assign add_71849 = add_71839 + 32'h0000_0001;
  assign array_update_71850[0] = add_71847 == 32'h0000_0000 ? TestBlock__A_op83 : array_index_71846[0];
  assign array_update_71850[1] = add_71847 == 32'h0000_0001 ? TestBlock__A_op83 : array_index_71846[1];
  assign array_update_71850[2] = add_71847 == 32'h0000_0002 ? TestBlock__A_op83 : array_index_71846[2];
  assign array_update_71850[3] = add_71847 == 32'h0000_0003 ? TestBlock__A_op83 : array_index_71846[3];
  assign array_update_71850[4] = add_71847 == 32'h0000_0004 ? TestBlock__A_op83 : array_index_71846[4];
  assign array_update_71850[5] = add_71847 == 32'h0000_0005 ? TestBlock__A_op83 : array_index_71846[5];
  assign array_update_71850[6] = add_71847 == 32'h0000_0006 ? TestBlock__A_op83 : array_index_71846[6];
  assign array_update_71850[7] = add_71847 == 32'h0000_0007 ? TestBlock__A_op83 : array_index_71846[7];
  assign array_update_71850[8] = add_71847 == 32'h0000_0008 ? TestBlock__A_op83 : array_index_71846[8];
  assign array_update_71850[9] = add_71847 == 32'h0000_0009 ? TestBlock__A_op83 : array_index_71846[9];
  assign array_update_71851[0] = add_71849 == 32'h0000_0000 ? TestBlock__B_op83 : array_index_71848[0];
  assign array_update_71851[1] = add_71849 == 32'h0000_0001 ? TestBlock__B_op83 : array_index_71848[1];
  assign array_update_71851[2] = add_71849 == 32'h0000_0002 ? TestBlock__B_op83 : array_index_71848[2];
  assign array_update_71851[3] = add_71849 == 32'h0000_0003 ? TestBlock__B_op83 : array_index_71848[3];
  assign array_update_71851[4] = add_71849 == 32'h0000_0004 ? TestBlock__B_op83 : array_index_71848[4];
  assign array_update_71851[5] = add_71849 == 32'h0000_0005 ? TestBlock__B_op83 : array_index_71848[5];
  assign array_update_71851[6] = add_71849 == 32'h0000_0006 ? TestBlock__B_op83 : array_index_71848[6];
  assign array_update_71851[7] = add_71849 == 32'h0000_0007 ? TestBlock__B_op83 : array_index_71848[7];
  assign array_update_71851[8] = add_71849 == 32'h0000_0008 ? TestBlock__B_op83 : array_index_71848[8];
  assign array_update_71851[9] = add_71849 == 32'h0000_0009 ? TestBlock__B_op83 : array_index_71848[9];
  assign array_update_71852[0] = add_71813 == 32'h0000_0000 ? array_update_71850 : array_update_71842[0];
  assign array_update_71852[1] = add_71813 == 32'h0000_0001 ? array_update_71850 : array_update_71842[1];
  assign array_update_71852[2] = add_71813 == 32'h0000_0002 ? array_update_71850 : array_update_71842[2];
  assign array_update_71852[3] = add_71813 == 32'h0000_0003 ? array_update_71850 : array_update_71842[3];
  assign array_update_71852[4] = add_71813 == 32'h0000_0004 ? array_update_71850 : array_update_71842[4];
  assign array_update_71852[5] = add_71813 == 32'h0000_0005 ? array_update_71850 : array_update_71842[5];
  assign array_update_71852[6] = add_71813 == 32'h0000_0006 ? array_update_71850 : array_update_71842[6];
  assign array_update_71852[7] = add_71813 == 32'h0000_0007 ? array_update_71850 : array_update_71842[7];
  assign array_update_71852[8] = add_71813 == 32'h0000_0008 ? array_update_71850 : array_update_71842[8];
  assign array_update_71852[9] = add_71813 == 32'h0000_0009 ? array_update_71850 : array_update_71842[9];
  assign array_update_71854[0] = add_71815 == 32'h0000_0000 ? array_update_71851 : array_update_71844[0];
  assign array_update_71854[1] = add_71815 == 32'h0000_0001 ? array_update_71851 : array_update_71844[1];
  assign array_update_71854[2] = add_71815 == 32'h0000_0002 ? array_update_71851 : array_update_71844[2];
  assign array_update_71854[3] = add_71815 == 32'h0000_0003 ? array_update_71851 : array_update_71844[3];
  assign array_update_71854[4] = add_71815 == 32'h0000_0004 ? array_update_71851 : array_update_71844[4];
  assign array_update_71854[5] = add_71815 == 32'h0000_0005 ? array_update_71851 : array_update_71844[5];
  assign array_update_71854[6] = add_71815 == 32'h0000_0006 ? array_update_71851 : array_update_71844[6];
  assign array_update_71854[7] = add_71815 == 32'h0000_0007 ? array_update_71851 : array_update_71844[7];
  assign array_update_71854[8] = add_71815 == 32'h0000_0008 ? array_update_71851 : array_update_71844[8];
  assign array_update_71854[9] = add_71815 == 32'h0000_0009 ? array_update_71851 : array_update_71844[9];
  assign array_index_71856 = array_update_71852[add_71813 > 32'h0000_0009 ? 4'h9 : add_71813[3:0]];
  assign add_71857 = add_71847 + 32'h0000_0001;
  assign array_index_71858 = array_update_71854[add_71815 > 32'h0000_0009 ? 4'h9 : add_71815[3:0]];
  assign add_71859 = add_71849 + 32'h0000_0001;
  assign array_update_71860[0] = add_71857 == 32'h0000_0000 ? TestBlock__A_op84 : array_index_71856[0];
  assign array_update_71860[1] = add_71857 == 32'h0000_0001 ? TestBlock__A_op84 : array_index_71856[1];
  assign array_update_71860[2] = add_71857 == 32'h0000_0002 ? TestBlock__A_op84 : array_index_71856[2];
  assign array_update_71860[3] = add_71857 == 32'h0000_0003 ? TestBlock__A_op84 : array_index_71856[3];
  assign array_update_71860[4] = add_71857 == 32'h0000_0004 ? TestBlock__A_op84 : array_index_71856[4];
  assign array_update_71860[5] = add_71857 == 32'h0000_0005 ? TestBlock__A_op84 : array_index_71856[5];
  assign array_update_71860[6] = add_71857 == 32'h0000_0006 ? TestBlock__A_op84 : array_index_71856[6];
  assign array_update_71860[7] = add_71857 == 32'h0000_0007 ? TestBlock__A_op84 : array_index_71856[7];
  assign array_update_71860[8] = add_71857 == 32'h0000_0008 ? TestBlock__A_op84 : array_index_71856[8];
  assign array_update_71860[9] = add_71857 == 32'h0000_0009 ? TestBlock__A_op84 : array_index_71856[9];
  assign array_update_71861[0] = add_71859 == 32'h0000_0000 ? TestBlock__B_op84 : array_index_71858[0];
  assign array_update_71861[1] = add_71859 == 32'h0000_0001 ? TestBlock__B_op84 : array_index_71858[1];
  assign array_update_71861[2] = add_71859 == 32'h0000_0002 ? TestBlock__B_op84 : array_index_71858[2];
  assign array_update_71861[3] = add_71859 == 32'h0000_0003 ? TestBlock__B_op84 : array_index_71858[3];
  assign array_update_71861[4] = add_71859 == 32'h0000_0004 ? TestBlock__B_op84 : array_index_71858[4];
  assign array_update_71861[5] = add_71859 == 32'h0000_0005 ? TestBlock__B_op84 : array_index_71858[5];
  assign array_update_71861[6] = add_71859 == 32'h0000_0006 ? TestBlock__B_op84 : array_index_71858[6];
  assign array_update_71861[7] = add_71859 == 32'h0000_0007 ? TestBlock__B_op84 : array_index_71858[7];
  assign array_update_71861[8] = add_71859 == 32'h0000_0008 ? TestBlock__B_op84 : array_index_71858[8];
  assign array_update_71861[9] = add_71859 == 32'h0000_0009 ? TestBlock__B_op84 : array_index_71858[9];
  assign array_update_71862[0] = add_71813 == 32'h0000_0000 ? array_update_71860 : array_update_71852[0];
  assign array_update_71862[1] = add_71813 == 32'h0000_0001 ? array_update_71860 : array_update_71852[1];
  assign array_update_71862[2] = add_71813 == 32'h0000_0002 ? array_update_71860 : array_update_71852[2];
  assign array_update_71862[3] = add_71813 == 32'h0000_0003 ? array_update_71860 : array_update_71852[3];
  assign array_update_71862[4] = add_71813 == 32'h0000_0004 ? array_update_71860 : array_update_71852[4];
  assign array_update_71862[5] = add_71813 == 32'h0000_0005 ? array_update_71860 : array_update_71852[5];
  assign array_update_71862[6] = add_71813 == 32'h0000_0006 ? array_update_71860 : array_update_71852[6];
  assign array_update_71862[7] = add_71813 == 32'h0000_0007 ? array_update_71860 : array_update_71852[7];
  assign array_update_71862[8] = add_71813 == 32'h0000_0008 ? array_update_71860 : array_update_71852[8];
  assign array_update_71862[9] = add_71813 == 32'h0000_0009 ? array_update_71860 : array_update_71852[9];
  assign array_update_71864[0] = add_71815 == 32'h0000_0000 ? array_update_71861 : array_update_71854[0];
  assign array_update_71864[1] = add_71815 == 32'h0000_0001 ? array_update_71861 : array_update_71854[1];
  assign array_update_71864[2] = add_71815 == 32'h0000_0002 ? array_update_71861 : array_update_71854[2];
  assign array_update_71864[3] = add_71815 == 32'h0000_0003 ? array_update_71861 : array_update_71854[3];
  assign array_update_71864[4] = add_71815 == 32'h0000_0004 ? array_update_71861 : array_update_71854[4];
  assign array_update_71864[5] = add_71815 == 32'h0000_0005 ? array_update_71861 : array_update_71854[5];
  assign array_update_71864[6] = add_71815 == 32'h0000_0006 ? array_update_71861 : array_update_71854[6];
  assign array_update_71864[7] = add_71815 == 32'h0000_0007 ? array_update_71861 : array_update_71854[7];
  assign array_update_71864[8] = add_71815 == 32'h0000_0008 ? array_update_71861 : array_update_71854[8];
  assign array_update_71864[9] = add_71815 == 32'h0000_0009 ? array_update_71861 : array_update_71854[9];
  assign array_index_71866 = array_update_71862[add_71813 > 32'h0000_0009 ? 4'h9 : add_71813[3:0]];
  assign add_71867 = add_71857 + 32'h0000_0001;
  assign array_index_71868 = array_update_71864[add_71815 > 32'h0000_0009 ? 4'h9 : add_71815[3:0]];
  assign add_71869 = add_71859 + 32'h0000_0001;
  assign array_update_71870[0] = add_71867 == 32'h0000_0000 ? TestBlock__A_op85 : array_index_71866[0];
  assign array_update_71870[1] = add_71867 == 32'h0000_0001 ? TestBlock__A_op85 : array_index_71866[1];
  assign array_update_71870[2] = add_71867 == 32'h0000_0002 ? TestBlock__A_op85 : array_index_71866[2];
  assign array_update_71870[3] = add_71867 == 32'h0000_0003 ? TestBlock__A_op85 : array_index_71866[3];
  assign array_update_71870[4] = add_71867 == 32'h0000_0004 ? TestBlock__A_op85 : array_index_71866[4];
  assign array_update_71870[5] = add_71867 == 32'h0000_0005 ? TestBlock__A_op85 : array_index_71866[5];
  assign array_update_71870[6] = add_71867 == 32'h0000_0006 ? TestBlock__A_op85 : array_index_71866[6];
  assign array_update_71870[7] = add_71867 == 32'h0000_0007 ? TestBlock__A_op85 : array_index_71866[7];
  assign array_update_71870[8] = add_71867 == 32'h0000_0008 ? TestBlock__A_op85 : array_index_71866[8];
  assign array_update_71870[9] = add_71867 == 32'h0000_0009 ? TestBlock__A_op85 : array_index_71866[9];
  assign array_update_71871[0] = add_71869 == 32'h0000_0000 ? TestBlock__B_op85 : array_index_71868[0];
  assign array_update_71871[1] = add_71869 == 32'h0000_0001 ? TestBlock__B_op85 : array_index_71868[1];
  assign array_update_71871[2] = add_71869 == 32'h0000_0002 ? TestBlock__B_op85 : array_index_71868[2];
  assign array_update_71871[3] = add_71869 == 32'h0000_0003 ? TestBlock__B_op85 : array_index_71868[3];
  assign array_update_71871[4] = add_71869 == 32'h0000_0004 ? TestBlock__B_op85 : array_index_71868[4];
  assign array_update_71871[5] = add_71869 == 32'h0000_0005 ? TestBlock__B_op85 : array_index_71868[5];
  assign array_update_71871[6] = add_71869 == 32'h0000_0006 ? TestBlock__B_op85 : array_index_71868[6];
  assign array_update_71871[7] = add_71869 == 32'h0000_0007 ? TestBlock__B_op85 : array_index_71868[7];
  assign array_update_71871[8] = add_71869 == 32'h0000_0008 ? TestBlock__B_op85 : array_index_71868[8];
  assign array_update_71871[9] = add_71869 == 32'h0000_0009 ? TestBlock__B_op85 : array_index_71868[9];
  assign array_update_71872[0] = add_71813 == 32'h0000_0000 ? array_update_71870 : array_update_71862[0];
  assign array_update_71872[1] = add_71813 == 32'h0000_0001 ? array_update_71870 : array_update_71862[1];
  assign array_update_71872[2] = add_71813 == 32'h0000_0002 ? array_update_71870 : array_update_71862[2];
  assign array_update_71872[3] = add_71813 == 32'h0000_0003 ? array_update_71870 : array_update_71862[3];
  assign array_update_71872[4] = add_71813 == 32'h0000_0004 ? array_update_71870 : array_update_71862[4];
  assign array_update_71872[5] = add_71813 == 32'h0000_0005 ? array_update_71870 : array_update_71862[5];
  assign array_update_71872[6] = add_71813 == 32'h0000_0006 ? array_update_71870 : array_update_71862[6];
  assign array_update_71872[7] = add_71813 == 32'h0000_0007 ? array_update_71870 : array_update_71862[7];
  assign array_update_71872[8] = add_71813 == 32'h0000_0008 ? array_update_71870 : array_update_71862[8];
  assign array_update_71872[9] = add_71813 == 32'h0000_0009 ? array_update_71870 : array_update_71862[9];
  assign array_update_71874[0] = add_71815 == 32'h0000_0000 ? array_update_71871 : array_update_71864[0];
  assign array_update_71874[1] = add_71815 == 32'h0000_0001 ? array_update_71871 : array_update_71864[1];
  assign array_update_71874[2] = add_71815 == 32'h0000_0002 ? array_update_71871 : array_update_71864[2];
  assign array_update_71874[3] = add_71815 == 32'h0000_0003 ? array_update_71871 : array_update_71864[3];
  assign array_update_71874[4] = add_71815 == 32'h0000_0004 ? array_update_71871 : array_update_71864[4];
  assign array_update_71874[5] = add_71815 == 32'h0000_0005 ? array_update_71871 : array_update_71864[5];
  assign array_update_71874[6] = add_71815 == 32'h0000_0006 ? array_update_71871 : array_update_71864[6];
  assign array_update_71874[7] = add_71815 == 32'h0000_0007 ? array_update_71871 : array_update_71864[7];
  assign array_update_71874[8] = add_71815 == 32'h0000_0008 ? array_update_71871 : array_update_71864[8];
  assign array_update_71874[9] = add_71815 == 32'h0000_0009 ? array_update_71871 : array_update_71864[9];
  assign array_index_71876 = array_update_71872[add_71813 > 32'h0000_0009 ? 4'h9 : add_71813[3:0]];
  assign add_71877 = add_71867 + 32'h0000_0001;
  assign array_index_71878 = array_update_71874[add_71815 > 32'h0000_0009 ? 4'h9 : add_71815[3:0]];
  assign add_71879 = add_71869 + 32'h0000_0001;
  assign array_update_71880[0] = add_71877 == 32'h0000_0000 ? TestBlock__A_op86 : array_index_71876[0];
  assign array_update_71880[1] = add_71877 == 32'h0000_0001 ? TestBlock__A_op86 : array_index_71876[1];
  assign array_update_71880[2] = add_71877 == 32'h0000_0002 ? TestBlock__A_op86 : array_index_71876[2];
  assign array_update_71880[3] = add_71877 == 32'h0000_0003 ? TestBlock__A_op86 : array_index_71876[3];
  assign array_update_71880[4] = add_71877 == 32'h0000_0004 ? TestBlock__A_op86 : array_index_71876[4];
  assign array_update_71880[5] = add_71877 == 32'h0000_0005 ? TestBlock__A_op86 : array_index_71876[5];
  assign array_update_71880[6] = add_71877 == 32'h0000_0006 ? TestBlock__A_op86 : array_index_71876[6];
  assign array_update_71880[7] = add_71877 == 32'h0000_0007 ? TestBlock__A_op86 : array_index_71876[7];
  assign array_update_71880[8] = add_71877 == 32'h0000_0008 ? TestBlock__A_op86 : array_index_71876[8];
  assign array_update_71880[9] = add_71877 == 32'h0000_0009 ? TestBlock__A_op86 : array_index_71876[9];
  assign array_update_71881[0] = add_71879 == 32'h0000_0000 ? TestBlock__B_op86 : array_index_71878[0];
  assign array_update_71881[1] = add_71879 == 32'h0000_0001 ? TestBlock__B_op86 : array_index_71878[1];
  assign array_update_71881[2] = add_71879 == 32'h0000_0002 ? TestBlock__B_op86 : array_index_71878[2];
  assign array_update_71881[3] = add_71879 == 32'h0000_0003 ? TestBlock__B_op86 : array_index_71878[3];
  assign array_update_71881[4] = add_71879 == 32'h0000_0004 ? TestBlock__B_op86 : array_index_71878[4];
  assign array_update_71881[5] = add_71879 == 32'h0000_0005 ? TestBlock__B_op86 : array_index_71878[5];
  assign array_update_71881[6] = add_71879 == 32'h0000_0006 ? TestBlock__B_op86 : array_index_71878[6];
  assign array_update_71881[7] = add_71879 == 32'h0000_0007 ? TestBlock__B_op86 : array_index_71878[7];
  assign array_update_71881[8] = add_71879 == 32'h0000_0008 ? TestBlock__B_op86 : array_index_71878[8];
  assign array_update_71881[9] = add_71879 == 32'h0000_0009 ? TestBlock__B_op86 : array_index_71878[9];
  assign array_update_71882[0] = add_71813 == 32'h0000_0000 ? array_update_71880 : array_update_71872[0];
  assign array_update_71882[1] = add_71813 == 32'h0000_0001 ? array_update_71880 : array_update_71872[1];
  assign array_update_71882[2] = add_71813 == 32'h0000_0002 ? array_update_71880 : array_update_71872[2];
  assign array_update_71882[3] = add_71813 == 32'h0000_0003 ? array_update_71880 : array_update_71872[3];
  assign array_update_71882[4] = add_71813 == 32'h0000_0004 ? array_update_71880 : array_update_71872[4];
  assign array_update_71882[5] = add_71813 == 32'h0000_0005 ? array_update_71880 : array_update_71872[5];
  assign array_update_71882[6] = add_71813 == 32'h0000_0006 ? array_update_71880 : array_update_71872[6];
  assign array_update_71882[7] = add_71813 == 32'h0000_0007 ? array_update_71880 : array_update_71872[7];
  assign array_update_71882[8] = add_71813 == 32'h0000_0008 ? array_update_71880 : array_update_71872[8];
  assign array_update_71882[9] = add_71813 == 32'h0000_0009 ? array_update_71880 : array_update_71872[9];
  assign array_update_71884[0] = add_71815 == 32'h0000_0000 ? array_update_71881 : array_update_71874[0];
  assign array_update_71884[1] = add_71815 == 32'h0000_0001 ? array_update_71881 : array_update_71874[1];
  assign array_update_71884[2] = add_71815 == 32'h0000_0002 ? array_update_71881 : array_update_71874[2];
  assign array_update_71884[3] = add_71815 == 32'h0000_0003 ? array_update_71881 : array_update_71874[3];
  assign array_update_71884[4] = add_71815 == 32'h0000_0004 ? array_update_71881 : array_update_71874[4];
  assign array_update_71884[5] = add_71815 == 32'h0000_0005 ? array_update_71881 : array_update_71874[5];
  assign array_update_71884[6] = add_71815 == 32'h0000_0006 ? array_update_71881 : array_update_71874[6];
  assign array_update_71884[7] = add_71815 == 32'h0000_0007 ? array_update_71881 : array_update_71874[7];
  assign array_update_71884[8] = add_71815 == 32'h0000_0008 ? array_update_71881 : array_update_71874[8];
  assign array_update_71884[9] = add_71815 == 32'h0000_0009 ? array_update_71881 : array_update_71874[9];
  assign array_index_71886 = array_update_71882[add_71813 > 32'h0000_0009 ? 4'h9 : add_71813[3:0]];
  assign add_71887 = add_71877 + 32'h0000_0001;
  assign array_index_71888 = array_update_71884[add_71815 > 32'h0000_0009 ? 4'h9 : add_71815[3:0]];
  assign add_71889 = add_71879 + 32'h0000_0001;
  assign array_update_71890[0] = add_71887 == 32'h0000_0000 ? TestBlock__A_op87 : array_index_71886[0];
  assign array_update_71890[1] = add_71887 == 32'h0000_0001 ? TestBlock__A_op87 : array_index_71886[1];
  assign array_update_71890[2] = add_71887 == 32'h0000_0002 ? TestBlock__A_op87 : array_index_71886[2];
  assign array_update_71890[3] = add_71887 == 32'h0000_0003 ? TestBlock__A_op87 : array_index_71886[3];
  assign array_update_71890[4] = add_71887 == 32'h0000_0004 ? TestBlock__A_op87 : array_index_71886[4];
  assign array_update_71890[5] = add_71887 == 32'h0000_0005 ? TestBlock__A_op87 : array_index_71886[5];
  assign array_update_71890[6] = add_71887 == 32'h0000_0006 ? TestBlock__A_op87 : array_index_71886[6];
  assign array_update_71890[7] = add_71887 == 32'h0000_0007 ? TestBlock__A_op87 : array_index_71886[7];
  assign array_update_71890[8] = add_71887 == 32'h0000_0008 ? TestBlock__A_op87 : array_index_71886[8];
  assign array_update_71890[9] = add_71887 == 32'h0000_0009 ? TestBlock__A_op87 : array_index_71886[9];
  assign array_update_71891[0] = add_71889 == 32'h0000_0000 ? TestBlock__B_op87 : array_index_71888[0];
  assign array_update_71891[1] = add_71889 == 32'h0000_0001 ? TestBlock__B_op87 : array_index_71888[1];
  assign array_update_71891[2] = add_71889 == 32'h0000_0002 ? TestBlock__B_op87 : array_index_71888[2];
  assign array_update_71891[3] = add_71889 == 32'h0000_0003 ? TestBlock__B_op87 : array_index_71888[3];
  assign array_update_71891[4] = add_71889 == 32'h0000_0004 ? TestBlock__B_op87 : array_index_71888[4];
  assign array_update_71891[5] = add_71889 == 32'h0000_0005 ? TestBlock__B_op87 : array_index_71888[5];
  assign array_update_71891[6] = add_71889 == 32'h0000_0006 ? TestBlock__B_op87 : array_index_71888[6];
  assign array_update_71891[7] = add_71889 == 32'h0000_0007 ? TestBlock__B_op87 : array_index_71888[7];
  assign array_update_71891[8] = add_71889 == 32'h0000_0008 ? TestBlock__B_op87 : array_index_71888[8];
  assign array_update_71891[9] = add_71889 == 32'h0000_0009 ? TestBlock__B_op87 : array_index_71888[9];
  assign array_update_71892[0] = add_71813 == 32'h0000_0000 ? array_update_71890 : array_update_71882[0];
  assign array_update_71892[1] = add_71813 == 32'h0000_0001 ? array_update_71890 : array_update_71882[1];
  assign array_update_71892[2] = add_71813 == 32'h0000_0002 ? array_update_71890 : array_update_71882[2];
  assign array_update_71892[3] = add_71813 == 32'h0000_0003 ? array_update_71890 : array_update_71882[3];
  assign array_update_71892[4] = add_71813 == 32'h0000_0004 ? array_update_71890 : array_update_71882[4];
  assign array_update_71892[5] = add_71813 == 32'h0000_0005 ? array_update_71890 : array_update_71882[5];
  assign array_update_71892[6] = add_71813 == 32'h0000_0006 ? array_update_71890 : array_update_71882[6];
  assign array_update_71892[7] = add_71813 == 32'h0000_0007 ? array_update_71890 : array_update_71882[7];
  assign array_update_71892[8] = add_71813 == 32'h0000_0008 ? array_update_71890 : array_update_71882[8];
  assign array_update_71892[9] = add_71813 == 32'h0000_0009 ? array_update_71890 : array_update_71882[9];
  assign array_update_71894[0] = add_71815 == 32'h0000_0000 ? array_update_71891 : array_update_71884[0];
  assign array_update_71894[1] = add_71815 == 32'h0000_0001 ? array_update_71891 : array_update_71884[1];
  assign array_update_71894[2] = add_71815 == 32'h0000_0002 ? array_update_71891 : array_update_71884[2];
  assign array_update_71894[3] = add_71815 == 32'h0000_0003 ? array_update_71891 : array_update_71884[3];
  assign array_update_71894[4] = add_71815 == 32'h0000_0004 ? array_update_71891 : array_update_71884[4];
  assign array_update_71894[5] = add_71815 == 32'h0000_0005 ? array_update_71891 : array_update_71884[5];
  assign array_update_71894[6] = add_71815 == 32'h0000_0006 ? array_update_71891 : array_update_71884[6];
  assign array_update_71894[7] = add_71815 == 32'h0000_0007 ? array_update_71891 : array_update_71884[7];
  assign array_update_71894[8] = add_71815 == 32'h0000_0008 ? array_update_71891 : array_update_71884[8];
  assign array_update_71894[9] = add_71815 == 32'h0000_0009 ? array_update_71891 : array_update_71884[9];
  assign array_index_71896 = array_update_71892[add_71813 > 32'h0000_0009 ? 4'h9 : add_71813[3:0]];
  assign add_71897 = add_71887 + 32'h0000_0001;
  assign array_index_71898 = array_update_71894[add_71815 > 32'h0000_0009 ? 4'h9 : add_71815[3:0]];
  assign add_71899 = add_71889 + 32'h0000_0001;
  assign array_update_71900[0] = add_71897 == 32'h0000_0000 ? TestBlock__A_op88 : array_index_71896[0];
  assign array_update_71900[1] = add_71897 == 32'h0000_0001 ? TestBlock__A_op88 : array_index_71896[1];
  assign array_update_71900[2] = add_71897 == 32'h0000_0002 ? TestBlock__A_op88 : array_index_71896[2];
  assign array_update_71900[3] = add_71897 == 32'h0000_0003 ? TestBlock__A_op88 : array_index_71896[3];
  assign array_update_71900[4] = add_71897 == 32'h0000_0004 ? TestBlock__A_op88 : array_index_71896[4];
  assign array_update_71900[5] = add_71897 == 32'h0000_0005 ? TestBlock__A_op88 : array_index_71896[5];
  assign array_update_71900[6] = add_71897 == 32'h0000_0006 ? TestBlock__A_op88 : array_index_71896[6];
  assign array_update_71900[7] = add_71897 == 32'h0000_0007 ? TestBlock__A_op88 : array_index_71896[7];
  assign array_update_71900[8] = add_71897 == 32'h0000_0008 ? TestBlock__A_op88 : array_index_71896[8];
  assign array_update_71900[9] = add_71897 == 32'h0000_0009 ? TestBlock__A_op88 : array_index_71896[9];
  assign array_update_71901[0] = add_71899 == 32'h0000_0000 ? TestBlock__B_op88 : array_index_71898[0];
  assign array_update_71901[1] = add_71899 == 32'h0000_0001 ? TestBlock__B_op88 : array_index_71898[1];
  assign array_update_71901[2] = add_71899 == 32'h0000_0002 ? TestBlock__B_op88 : array_index_71898[2];
  assign array_update_71901[3] = add_71899 == 32'h0000_0003 ? TestBlock__B_op88 : array_index_71898[3];
  assign array_update_71901[4] = add_71899 == 32'h0000_0004 ? TestBlock__B_op88 : array_index_71898[4];
  assign array_update_71901[5] = add_71899 == 32'h0000_0005 ? TestBlock__B_op88 : array_index_71898[5];
  assign array_update_71901[6] = add_71899 == 32'h0000_0006 ? TestBlock__B_op88 : array_index_71898[6];
  assign array_update_71901[7] = add_71899 == 32'h0000_0007 ? TestBlock__B_op88 : array_index_71898[7];
  assign array_update_71901[8] = add_71899 == 32'h0000_0008 ? TestBlock__B_op88 : array_index_71898[8];
  assign array_update_71901[9] = add_71899 == 32'h0000_0009 ? TestBlock__B_op88 : array_index_71898[9];
  assign array_update_71902[0] = add_71813 == 32'h0000_0000 ? array_update_71900 : array_update_71892[0];
  assign array_update_71902[1] = add_71813 == 32'h0000_0001 ? array_update_71900 : array_update_71892[1];
  assign array_update_71902[2] = add_71813 == 32'h0000_0002 ? array_update_71900 : array_update_71892[2];
  assign array_update_71902[3] = add_71813 == 32'h0000_0003 ? array_update_71900 : array_update_71892[3];
  assign array_update_71902[4] = add_71813 == 32'h0000_0004 ? array_update_71900 : array_update_71892[4];
  assign array_update_71902[5] = add_71813 == 32'h0000_0005 ? array_update_71900 : array_update_71892[5];
  assign array_update_71902[6] = add_71813 == 32'h0000_0006 ? array_update_71900 : array_update_71892[6];
  assign array_update_71902[7] = add_71813 == 32'h0000_0007 ? array_update_71900 : array_update_71892[7];
  assign array_update_71902[8] = add_71813 == 32'h0000_0008 ? array_update_71900 : array_update_71892[8];
  assign array_update_71902[9] = add_71813 == 32'h0000_0009 ? array_update_71900 : array_update_71892[9];
  assign array_update_71904[0] = add_71815 == 32'h0000_0000 ? array_update_71901 : array_update_71894[0];
  assign array_update_71904[1] = add_71815 == 32'h0000_0001 ? array_update_71901 : array_update_71894[1];
  assign array_update_71904[2] = add_71815 == 32'h0000_0002 ? array_update_71901 : array_update_71894[2];
  assign array_update_71904[3] = add_71815 == 32'h0000_0003 ? array_update_71901 : array_update_71894[3];
  assign array_update_71904[4] = add_71815 == 32'h0000_0004 ? array_update_71901 : array_update_71894[4];
  assign array_update_71904[5] = add_71815 == 32'h0000_0005 ? array_update_71901 : array_update_71894[5];
  assign array_update_71904[6] = add_71815 == 32'h0000_0006 ? array_update_71901 : array_update_71894[6];
  assign array_update_71904[7] = add_71815 == 32'h0000_0007 ? array_update_71901 : array_update_71894[7];
  assign array_update_71904[8] = add_71815 == 32'h0000_0008 ? array_update_71901 : array_update_71894[8];
  assign array_update_71904[9] = add_71815 == 32'h0000_0009 ? array_update_71901 : array_update_71894[9];
  assign array_index_71906 = array_update_71902[add_71813 > 32'h0000_0009 ? 4'h9 : add_71813[3:0]];
  assign add_71907 = add_71897 + 32'h0000_0001;
  assign array_index_71908 = array_update_71904[add_71815 > 32'h0000_0009 ? 4'h9 : add_71815[3:0]];
  assign add_71909 = add_71899 + 32'h0000_0001;
  assign array_update_71910[0] = add_71907 == 32'h0000_0000 ? TestBlock__A_op89 : array_index_71906[0];
  assign array_update_71910[1] = add_71907 == 32'h0000_0001 ? TestBlock__A_op89 : array_index_71906[1];
  assign array_update_71910[2] = add_71907 == 32'h0000_0002 ? TestBlock__A_op89 : array_index_71906[2];
  assign array_update_71910[3] = add_71907 == 32'h0000_0003 ? TestBlock__A_op89 : array_index_71906[3];
  assign array_update_71910[4] = add_71907 == 32'h0000_0004 ? TestBlock__A_op89 : array_index_71906[4];
  assign array_update_71910[5] = add_71907 == 32'h0000_0005 ? TestBlock__A_op89 : array_index_71906[5];
  assign array_update_71910[6] = add_71907 == 32'h0000_0006 ? TestBlock__A_op89 : array_index_71906[6];
  assign array_update_71910[7] = add_71907 == 32'h0000_0007 ? TestBlock__A_op89 : array_index_71906[7];
  assign array_update_71910[8] = add_71907 == 32'h0000_0008 ? TestBlock__A_op89 : array_index_71906[8];
  assign array_update_71910[9] = add_71907 == 32'h0000_0009 ? TestBlock__A_op89 : array_index_71906[9];
  assign array_update_71912[0] = add_71909 == 32'h0000_0000 ? TestBlock__B_op89 : array_index_71908[0];
  assign array_update_71912[1] = add_71909 == 32'h0000_0001 ? TestBlock__B_op89 : array_index_71908[1];
  assign array_update_71912[2] = add_71909 == 32'h0000_0002 ? TestBlock__B_op89 : array_index_71908[2];
  assign array_update_71912[3] = add_71909 == 32'h0000_0003 ? TestBlock__B_op89 : array_index_71908[3];
  assign array_update_71912[4] = add_71909 == 32'h0000_0004 ? TestBlock__B_op89 : array_index_71908[4];
  assign array_update_71912[5] = add_71909 == 32'h0000_0005 ? TestBlock__B_op89 : array_index_71908[5];
  assign array_update_71912[6] = add_71909 == 32'h0000_0006 ? TestBlock__B_op89 : array_index_71908[6];
  assign array_update_71912[7] = add_71909 == 32'h0000_0007 ? TestBlock__B_op89 : array_index_71908[7];
  assign array_update_71912[8] = add_71909 == 32'h0000_0008 ? TestBlock__B_op89 : array_index_71908[8];
  assign array_update_71912[9] = add_71909 == 32'h0000_0009 ? TestBlock__B_op89 : array_index_71908[9];
  assign array_update_71914[0] = add_71813 == 32'h0000_0000 ? array_update_71910 : array_update_71902[0];
  assign array_update_71914[1] = add_71813 == 32'h0000_0001 ? array_update_71910 : array_update_71902[1];
  assign array_update_71914[2] = add_71813 == 32'h0000_0002 ? array_update_71910 : array_update_71902[2];
  assign array_update_71914[3] = add_71813 == 32'h0000_0003 ? array_update_71910 : array_update_71902[3];
  assign array_update_71914[4] = add_71813 == 32'h0000_0004 ? array_update_71910 : array_update_71902[4];
  assign array_update_71914[5] = add_71813 == 32'h0000_0005 ? array_update_71910 : array_update_71902[5];
  assign array_update_71914[6] = add_71813 == 32'h0000_0006 ? array_update_71910 : array_update_71902[6];
  assign array_update_71914[7] = add_71813 == 32'h0000_0007 ? array_update_71910 : array_update_71902[7];
  assign array_update_71914[8] = add_71813 == 32'h0000_0008 ? array_update_71910 : array_update_71902[8];
  assign array_update_71914[9] = add_71813 == 32'h0000_0009 ? array_update_71910 : array_update_71902[9];
  assign add_71915 = add_71813 + 32'h0000_0001;
  assign array_update_71916[0] = add_71815 == 32'h0000_0000 ? array_update_71912 : array_update_71904[0];
  assign array_update_71916[1] = add_71815 == 32'h0000_0001 ? array_update_71912 : array_update_71904[1];
  assign array_update_71916[2] = add_71815 == 32'h0000_0002 ? array_update_71912 : array_update_71904[2];
  assign array_update_71916[3] = add_71815 == 32'h0000_0003 ? array_update_71912 : array_update_71904[3];
  assign array_update_71916[4] = add_71815 == 32'h0000_0004 ? array_update_71912 : array_update_71904[4];
  assign array_update_71916[5] = add_71815 == 32'h0000_0005 ? array_update_71912 : array_update_71904[5];
  assign array_update_71916[6] = add_71815 == 32'h0000_0006 ? array_update_71912 : array_update_71904[6];
  assign array_update_71916[7] = add_71815 == 32'h0000_0007 ? array_update_71912 : array_update_71904[7];
  assign array_update_71916[8] = add_71815 == 32'h0000_0008 ? array_update_71912 : array_update_71904[8];
  assign array_update_71916[9] = add_71815 == 32'h0000_0009 ? array_update_71912 : array_update_71904[9];
  assign add_71917 = add_71815 + 32'h0000_0001;
  assign array_index_71918 = array_update_71914[add_71915 > 32'h0000_0009 ? 4'h9 : add_71915[3:0]];
  assign literal_71919 = 32'h0000_0000;
  assign array_index_71920 = array_update_71916[add_71917 > 32'h0000_0009 ? 4'h9 : add_71917[3:0]];
  assign literal_71921 = 32'h0000_0000;
  assign array_update_71922[0] = literal_71919 == 32'h0000_0000 ? TestBlock__A_op90 : array_index_71918[0];
  assign array_update_71922[1] = literal_71919 == 32'h0000_0001 ? TestBlock__A_op90 : array_index_71918[1];
  assign array_update_71922[2] = literal_71919 == 32'h0000_0002 ? TestBlock__A_op90 : array_index_71918[2];
  assign array_update_71922[3] = literal_71919 == 32'h0000_0003 ? TestBlock__A_op90 : array_index_71918[3];
  assign array_update_71922[4] = literal_71919 == 32'h0000_0004 ? TestBlock__A_op90 : array_index_71918[4];
  assign array_update_71922[5] = literal_71919 == 32'h0000_0005 ? TestBlock__A_op90 : array_index_71918[5];
  assign array_update_71922[6] = literal_71919 == 32'h0000_0006 ? TestBlock__A_op90 : array_index_71918[6];
  assign array_update_71922[7] = literal_71919 == 32'h0000_0007 ? TestBlock__A_op90 : array_index_71918[7];
  assign array_update_71922[8] = literal_71919 == 32'h0000_0008 ? TestBlock__A_op90 : array_index_71918[8];
  assign array_update_71922[9] = literal_71919 == 32'h0000_0009 ? TestBlock__A_op90 : array_index_71918[9];
  assign array_update_71923[0] = literal_71921 == 32'h0000_0000 ? TestBlock__B_op90 : array_index_71920[0];
  assign array_update_71923[1] = literal_71921 == 32'h0000_0001 ? TestBlock__B_op90 : array_index_71920[1];
  assign array_update_71923[2] = literal_71921 == 32'h0000_0002 ? TestBlock__B_op90 : array_index_71920[2];
  assign array_update_71923[3] = literal_71921 == 32'h0000_0003 ? TestBlock__B_op90 : array_index_71920[3];
  assign array_update_71923[4] = literal_71921 == 32'h0000_0004 ? TestBlock__B_op90 : array_index_71920[4];
  assign array_update_71923[5] = literal_71921 == 32'h0000_0005 ? TestBlock__B_op90 : array_index_71920[5];
  assign array_update_71923[6] = literal_71921 == 32'h0000_0006 ? TestBlock__B_op90 : array_index_71920[6];
  assign array_update_71923[7] = literal_71921 == 32'h0000_0007 ? TestBlock__B_op90 : array_index_71920[7];
  assign array_update_71923[8] = literal_71921 == 32'h0000_0008 ? TestBlock__B_op90 : array_index_71920[8];
  assign array_update_71923[9] = literal_71921 == 32'h0000_0009 ? TestBlock__B_op90 : array_index_71920[9];
  assign array_update_71924[0] = add_71915 == 32'h0000_0000 ? array_update_71922 : array_update_71914[0];
  assign array_update_71924[1] = add_71915 == 32'h0000_0001 ? array_update_71922 : array_update_71914[1];
  assign array_update_71924[2] = add_71915 == 32'h0000_0002 ? array_update_71922 : array_update_71914[2];
  assign array_update_71924[3] = add_71915 == 32'h0000_0003 ? array_update_71922 : array_update_71914[3];
  assign array_update_71924[4] = add_71915 == 32'h0000_0004 ? array_update_71922 : array_update_71914[4];
  assign array_update_71924[5] = add_71915 == 32'h0000_0005 ? array_update_71922 : array_update_71914[5];
  assign array_update_71924[6] = add_71915 == 32'h0000_0006 ? array_update_71922 : array_update_71914[6];
  assign array_update_71924[7] = add_71915 == 32'h0000_0007 ? array_update_71922 : array_update_71914[7];
  assign array_update_71924[8] = add_71915 == 32'h0000_0008 ? array_update_71922 : array_update_71914[8];
  assign array_update_71924[9] = add_71915 == 32'h0000_0009 ? array_update_71922 : array_update_71914[9];
  assign array_update_71926[0] = add_71917 == 32'h0000_0000 ? array_update_71923 : array_update_71916[0];
  assign array_update_71926[1] = add_71917 == 32'h0000_0001 ? array_update_71923 : array_update_71916[1];
  assign array_update_71926[2] = add_71917 == 32'h0000_0002 ? array_update_71923 : array_update_71916[2];
  assign array_update_71926[3] = add_71917 == 32'h0000_0003 ? array_update_71923 : array_update_71916[3];
  assign array_update_71926[4] = add_71917 == 32'h0000_0004 ? array_update_71923 : array_update_71916[4];
  assign array_update_71926[5] = add_71917 == 32'h0000_0005 ? array_update_71923 : array_update_71916[5];
  assign array_update_71926[6] = add_71917 == 32'h0000_0006 ? array_update_71923 : array_update_71916[6];
  assign array_update_71926[7] = add_71917 == 32'h0000_0007 ? array_update_71923 : array_update_71916[7];
  assign array_update_71926[8] = add_71917 == 32'h0000_0008 ? array_update_71923 : array_update_71916[8];
  assign array_update_71926[9] = add_71917 == 32'h0000_0009 ? array_update_71923 : array_update_71916[9];
  assign array_index_71928 = array_update_71924[add_71915 > 32'h0000_0009 ? 4'h9 : add_71915[3:0]];
  assign add_71929 = literal_71919 + 32'h0000_0001;
  assign array_index_71930 = array_update_71926[add_71917 > 32'h0000_0009 ? 4'h9 : add_71917[3:0]];
  assign add_71931 = literal_71921 + 32'h0000_0001;
  assign array_update_71932[0] = add_71929 == 32'h0000_0000 ? TestBlock__A_op91 : array_index_71928[0];
  assign array_update_71932[1] = add_71929 == 32'h0000_0001 ? TestBlock__A_op91 : array_index_71928[1];
  assign array_update_71932[2] = add_71929 == 32'h0000_0002 ? TestBlock__A_op91 : array_index_71928[2];
  assign array_update_71932[3] = add_71929 == 32'h0000_0003 ? TestBlock__A_op91 : array_index_71928[3];
  assign array_update_71932[4] = add_71929 == 32'h0000_0004 ? TestBlock__A_op91 : array_index_71928[4];
  assign array_update_71932[5] = add_71929 == 32'h0000_0005 ? TestBlock__A_op91 : array_index_71928[5];
  assign array_update_71932[6] = add_71929 == 32'h0000_0006 ? TestBlock__A_op91 : array_index_71928[6];
  assign array_update_71932[7] = add_71929 == 32'h0000_0007 ? TestBlock__A_op91 : array_index_71928[7];
  assign array_update_71932[8] = add_71929 == 32'h0000_0008 ? TestBlock__A_op91 : array_index_71928[8];
  assign array_update_71932[9] = add_71929 == 32'h0000_0009 ? TestBlock__A_op91 : array_index_71928[9];
  assign array_update_71933[0] = add_71931 == 32'h0000_0000 ? TestBlock__B_op91 : array_index_71930[0];
  assign array_update_71933[1] = add_71931 == 32'h0000_0001 ? TestBlock__B_op91 : array_index_71930[1];
  assign array_update_71933[2] = add_71931 == 32'h0000_0002 ? TestBlock__B_op91 : array_index_71930[2];
  assign array_update_71933[3] = add_71931 == 32'h0000_0003 ? TestBlock__B_op91 : array_index_71930[3];
  assign array_update_71933[4] = add_71931 == 32'h0000_0004 ? TestBlock__B_op91 : array_index_71930[4];
  assign array_update_71933[5] = add_71931 == 32'h0000_0005 ? TestBlock__B_op91 : array_index_71930[5];
  assign array_update_71933[6] = add_71931 == 32'h0000_0006 ? TestBlock__B_op91 : array_index_71930[6];
  assign array_update_71933[7] = add_71931 == 32'h0000_0007 ? TestBlock__B_op91 : array_index_71930[7];
  assign array_update_71933[8] = add_71931 == 32'h0000_0008 ? TestBlock__B_op91 : array_index_71930[8];
  assign array_update_71933[9] = add_71931 == 32'h0000_0009 ? TestBlock__B_op91 : array_index_71930[9];
  assign array_update_71934[0] = add_71915 == 32'h0000_0000 ? array_update_71932 : array_update_71924[0];
  assign array_update_71934[1] = add_71915 == 32'h0000_0001 ? array_update_71932 : array_update_71924[1];
  assign array_update_71934[2] = add_71915 == 32'h0000_0002 ? array_update_71932 : array_update_71924[2];
  assign array_update_71934[3] = add_71915 == 32'h0000_0003 ? array_update_71932 : array_update_71924[3];
  assign array_update_71934[4] = add_71915 == 32'h0000_0004 ? array_update_71932 : array_update_71924[4];
  assign array_update_71934[5] = add_71915 == 32'h0000_0005 ? array_update_71932 : array_update_71924[5];
  assign array_update_71934[6] = add_71915 == 32'h0000_0006 ? array_update_71932 : array_update_71924[6];
  assign array_update_71934[7] = add_71915 == 32'h0000_0007 ? array_update_71932 : array_update_71924[7];
  assign array_update_71934[8] = add_71915 == 32'h0000_0008 ? array_update_71932 : array_update_71924[8];
  assign array_update_71934[9] = add_71915 == 32'h0000_0009 ? array_update_71932 : array_update_71924[9];
  assign array_update_71936[0] = add_71917 == 32'h0000_0000 ? array_update_71933 : array_update_71926[0];
  assign array_update_71936[1] = add_71917 == 32'h0000_0001 ? array_update_71933 : array_update_71926[1];
  assign array_update_71936[2] = add_71917 == 32'h0000_0002 ? array_update_71933 : array_update_71926[2];
  assign array_update_71936[3] = add_71917 == 32'h0000_0003 ? array_update_71933 : array_update_71926[3];
  assign array_update_71936[4] = add_71917 == 32'h0000_0004 ? array_update_71933 : array_update_71926[4];
  assign array_update_71936[5] = add_71917 == 32'h0000_0005 ? array_update_71933 : array_update_71926[5];
  assign array_update_71936[6] = add_71917 == 32'h0000_0006 ? array_update_71933 : array_update_71926[6];
  assign array_update_71936[7] = add_71917 == 32'h0000_0007 ? array_update_71933 : array_update_71926[7];
  assign array_update_71936[8] = add_71917 == 32'h0000_0008 ? array_update_71933 : array_update_71926[8];
  assign array_update_71936[9] = add_71917 == 32'h0000_0009 ? array_update_71933 : array_update_71926[9];
  assign array_index_71938 = array_update_71934[add_71915 > 32'h0000_0009 ? 4'h9 : add_71915[3:0]];
  assign add_71939 = add_71929 + 32'h0000_0001;
  assign array_index_71940 = array_update_71936[add_71917 > 32'h0000_0009 ? 4'h9 : add_71917[3:0]];
  assign add_71941 = add_71931 + 32'h0000_0001;
  assign array_update_71942[0] = add_71939 == 32'h0000_0000 ? TestBlock__A_op92 : array_index_71938[0];
  assign array_update_71942[1] = add_71939 == 32'h0000_0001 ? TestBlock__A_op92 : array_index_71938[1];
  assign array_update_71942[2] = add_71939 == 32'h0000_0002 ? TestBlock__A_op92 : array_index_71938[2];
  assign array_update_71942[3] = add_71939 == 32'h0000_0003 ? TestBlock__A_op92 : array_index_71938[3];
  assign array_update_71942[4] = add_71939 == 32'h0000_0004 ? TestBlock__A_op92 : array_index_71938[4];
  assign array_update_71942[5] = add_71939 == 32'h0000_0005 ? TestBlock__A_op92 : array_index_71938[5];
  assign array_update_71942[6] = add_71939 == 32'h0000_0006 ? TestBlock__A_op92 : array_index_71938[6];
  assign array_update_71942[7] = add_71939 == 32'h0000_0007 ? TestBlock__A_op92 : array_index_71938[7];
  assign array_update_71942[8] = add_71939 == 32'h0000_0008 ? TestBlock__A_op92 : array_index_71938[8];
  assign array_update_71942[9] = add_71939 == 32'h0000_0009 ? TestBlock__A_op92 : array_index_71938[9];
  assign array_update_71943[0] = add_71941 == 32'h0000_0000 ? TestBlock__B_op92 : array_index_71940[0];
  assign array_update_71943[1] = add_71941 == 32'h0000_0001 ? TestBlock__B_op92 : array_index_71940[1];
  assign array_update_71943[2] = add_71941 == 32'h0000_0002 ? TestBlock__B_op92 : array_index_71940[2];
  assign array_update_71943[3] = add_71941 == 32'h0000_0003 ? TestBlock__B_op92 : array_index_71940[3];
  assign array_update_71943[4] = add_71941 == 32'h0000_0004 ? TestBlock__B_op92 : array_index_71940[4];
  assign array_update_71943[5] = add_71941 == 32'h0000_0005 ? TestBlock__B_op92 : array_index_71940[5];
  assign array_update_71943[6] = add_71941 == 32'h0000_0006 ? TestBlock__B_op92 : array_index_71940[6];
  assign array_update_71943[7] = add_71941 == 32'h0000_0007 ? TestBlock__B_op92 : array_index_71940[7];
  assign array_update_71943[8] = add_71941 == 32'h0000_0008 ? TestBlock__B_op92 : array_index_71940[8];
  assign array_update_71943[9] = add_71941 == 32'h0000_0009 ? TestBlock__B_op92 : array_index_71940[9];
  assign array_update_71944[0] = add_71915 == 32'h0000_0000 ? array_update_71942 : array_update_71934[0];
  assign array_update_71944[1] = add_71915 == 32'h0000_0001 ? array_update_71942 : array_update_71934[1];
  assign array_update_71944[2] = add_71915 == 32'h0000_0002 ? array_update_71942 : array_update_71934[2];
  assign array_update_71944[3] = add_71915 == 32'h0000_0003 ? array_update_71942 : array_update_71934[3];
  assign array_update_71944[4] = add_71915 == 32'h0000_0004 ? array_update_71942 : array_update_71934[4];
  assign array_update_71944[5] = add_71915 == 32'h0000_0005 ? array_update_71942 : array_update_71934[5];
  assign array_update_71944[6] = add_71915 == 32'h0000_0006 ? array_update_71942 : array_update_71934[6];
  assign array_update_71944[7] = add_71915 == 32'h0000_0007 ? array_update_71942 : array_update_71934[7];
  assign array_update_71944[8] = add_71915 == 32'h0000_0008 ? array_update_71942 : array_update_71934[8];
  assign array_update_71944[9] = add_71915 == 32'h0000_0009 ? array_update_71942 : array_update_71934[9];
  assign array_update_71946[0] = add_71917 == 32'h0000_0000 ? array_update_71943 : array_update_71936[0];
  assign array_update_71946[1] = add_71917 == 32'h0000_0001 ? array_update_71943 : array_update_71936[1];
  assign array_update_71946[2] = add_71917 == 32'h0000_0002 ? array_update_71943 : array_update_71936[2];
  assign array_update_71946[3] = add_71917 == 32'h0000_0003 ? array_update_71943 : array_update_71936[3];
  assign array_update_71946[4] = add_71917 == 32'h0000_0004 ? array_update_71943 : array_update_71936[4];
  assign array_update_71946[5] = add_71917 == 32'h0000_0005 ? array_update_71943 : array_update_71936[5];
  assign array_update_71946[6] = add_71917 == 32'h0000_0006 ? array_update_71943 : array_update_71936[6];
  assign array_update_71946[7] = add_71917 == 32'h0000_0007 ? array_update_71943 : array_update_71936[7];
  assign array_update_71946[8] = add_71917 == 32'h0000_0008 ? array_update_71943 : array_update_71936[8];
  assign array_update_71946[9] = add_71917 == 32'h0000_0009 ? array_update_71943 : array_update_71936[9];
  assign array_index_71948 = array_update_71944[add_71915 > 32'h0000_0009 ? 4'h9 : add_71915[3:0]];
  assign add_71949 = add_71939 + 32'h0000_0001;
  assign array_index_71950 = array_update_71946[add_71917 > 32'h0000_0009 ? 4'h9 : add_71917[3:0]];
  assign add_71951 = add_71941 + 32'h0000_0001;
  assign array_update_71952[0] = add_71949 == 32'h0000_0000 ? TestBlock__A_op93 : array_index_71948[0];
  assign array_update_71952[1] = add_71949 == 32'h0000_0001 ? TestBlock__A_op93 : array_index_71948[1];
  assign array_update_71952[2] = add_71949 == 32'h0000_0002 ? TestBlock__A_op93 : array_index_71948[2];
  assign array_update_71952[3] = add_71949 == 32'h0000_0003 ? TestBlock__A_op93 : array_index_71948[3];
  assign array_update_71952[4] = add_71949 == 32'h0000_0004 ? TestBlock__A_op93 : array_index_71948[4];
  assign array_update_71952[5] = add_71949 == 32'h0000_0005 ? TestBlock__A_op93 : array_index_71948[5];
  assign array_update_71952[6] = add_71949 == 32'h0000_0006 ? TestBlock__A_op93 : array_index_71948[6];
  assign array_update_71952[7] = add_71949 == 32'h0000_0007 ? TestBlock__A_op93 : array_index_71948[7];
  assign array_update_71952[8] = add_71949 == 32'h0000_0008 ? TestBlock__A_op93 : array_index_71948[8];
  assign array_update_71952[9] = add_71949 == 32'h0000_0009 ? TestBlock__A_op93 : array_index_71948[9];
  assign array_update_71953[0] = add_71951 == 32'h0000_0000 ? TestBlock__B_op93 : array_index_71950[0];
  assign array_update_71953[1] = add_71951 == 32'h0000_0001 ? TestBlock__B_op93 : array_index_71950[1];
  assign array_update_71953[2] = add_71951 == 32'h0000_0002 ? TestBlock__B_op93 : array_index_71950[2];
  assign array_update_71953[3] = add_71951 == 32'h0000_0003 ? TestBlock__B_op93 : array_index_71950[3];
  assign array_update_71953[4] = add_71951 == 32'h0000_0004 ? TestBlock__B_op93 : array_index_71950[4];
  assign array_update_71953[5] = add_71951 == 32'h0000_0005 ? TestBlock__B_op93 : array_index_71950[5];
  assign array_update_71953[6] = add_71951 == 32'h0000_0006 ? TestBlock__B_op93 : array_index_71950[6];
  assign array_update_71953[7] = add_71951 == 32'h0000_0007 ? TestBlock__B_op93 : array_index_71950[7];
  assign array_update_71953[8] = add_71951 == 32'h0000_0008 ? TestBlock__B_op93 : array_index_71950[8];
  assign array_update_71953[9] = add_71951 == 32'h0000_0009 ? TestBlock__B_op93 : array_index_71950[9];
  assign array_update_71954[0] = add_71915 == 32'h0000_0000 ? array_update_71952 : array_update_71944[0];
  assign array_update_71954[1] = add_71915 == 32'h0000_0001 ? array_update_71952 : array_update_71944[1];
  assign array_update_71954[2] = add_71915 == 32'h0000_0002 ? array_update_71952 : array_update_71944[2];
  assign array_update_71954[3] = add_71915 == 32'h0000_0003 ? array_update_71952 : array_update_71944[3];
  assign array_update_71954[4] = add_71915 == 32'h0000_0004 ? array_update_71952 : array_update_71944[4];
  assign array_update_71954[5] = add_71915 == 32'h0000_0005 ? array_update_71952 : array_update_71944[5];
  assign array_update_71954[6] = add_71915 == 32'h0000_0006 ? array_update_71952 : array_update_71944[6];
  assign array_update_71954[7] = add_71915 == 32'h0000_0007 ? array_update_71952 : array_update_71944[7];
  assign array_update_71954[8] = add_71915 == 32'h0000_0008 ? array_update_71952 : array_update_71944[8];
  assign array_update_71954[9] = add_71915 == 32'h0000_0009 ? array_update_71952 : array_update_71944[9];
  assign array_update_71956[0] = add_71917 == 32'h0000_0000 ? array_update_71953 : array_update_71946[0];
  assign array_update_71956[1] = add_71917 == 32'h0000_0001 ? array_update_71953 : array_update_71946[1];
  assign array_update_71956[2] = add_71917 == 32'h0000_0002 ? array_update_71953 : array_update_71946[2];
  assign array_update_71956[3] = add_71917 == 32'h0000_0003 ? array_update_71953 : array_update_71946[3];
  assign array_update_71956[4] = add_71917 == 32'h0000_0004 ? array_update_71953 : array_update_71946[4];
  assign array_update_71956[5] = add_71917 == 32'h0000_0005 ? array_update_71953 : array_update_71946[5];
  assign array_update_71956[6] = add_71917 == 32'h0000_0006 ? array_update_71953 : array_update_71946[6];
  assign array_update_71956[7] = add_71917 == 32'h0000_0007 ? array_update_71953 : array_update_71946[7];
  assign array_update_71956[8] = add_71917 == 32'h0000_0008 ? array_update_71953 : array_update_71946[8];
  assign array_update_71956[9] = add_71917 == 32'h0000_0009 ? array_update_71953 : array_update_71946[9];
  assign array_index_71958 = array_update_71954[add_71915 > 32'h0000_0009 ? 4'h9 : add_71915[3:0]];
  assign add_71959 = add_71949 + 32'h0000_0001;
  assign array_index_71960 = array_update_71956[add_71917 > 32'h0000_0009 ? 4'h9 : add_71917[3:0]];
  assign add_71961 = add_71951 + 32'h0000_0001;
  assign array_update_71962[0] = add_71959 == 32'h0000_0000 ? TestBlock__A_op94 : array_index_71958[0];
  assign array_update_71962[1] = add_71959 == 32'h0000_0001 ? TestBlock__A_op94 : array_index_71958[1];
  assign array_update_71962[2] = add_71959 == 32'h0000_0002 ? TestBlock__A_op94 : array_index_71958[2];
  assign array_update_71962[3] = add_71959 == 32'h0000_0003 ? TestBlock__A_op94 : array_index_71958[3];
  assign array_update_71962[4] = add_71959 == 32'h0000_0004 ? TestBlock__A_op94 : array_index_71958[4];
  assign array_update_71962[5] = add_71959 == 32'h0000_0005 ? TestBlock__A_op94 : array_index_71958[5];
  assign array_update_71962[6] = add_71959 == 32'h0000_0006 ? TestBlock__A_op94 : array_index_71958[6];
  assign array_update_71962[7] = add_71959 == 32'h0000_0007 ? TestBlock__A_op94 : array_index_71958[7];
  assign array_update_71962[8] = add_71959 == 32'h0000_0008 ? TestBlock__A_op94 : array_index_71958[8];
  assign array_update_71962[9] = add_71959 == 32'h0000_0009 ? TestBlock__A_op94 : array_index_71958[9];
  assign array_update_71963[0] = add_71961 == 32'h0000_0000 ? TestBlock__B_op94 : array_index_71960[0];
  assign array_update_71963[1] = add_71961 == 32'h0000_0001 ? TestBlock__B_op94 : array_index_71960[1];
  assign array_update_71963[2] = add_71961 == 32'h0000_0002 ? TestBlock__B_op94 : array_index_71960[2];
  assign array_update_71963[3] = add_71961 == 32'h0000_0003 ? TestBlock__B_op94 : array_index_71960[3];
  assign array_update_71963[4] = add_71961 == 32'h0000_0004 ? TestBlock__B_op94 : array_index_71960[4];
  assign array_update_71963[5] = add_71961 == 32'h0000_0005 ? TestBlock__B_op94 : array_index_71960[5];
  assign array_update_71963[6] = add_71961 == 32'h0000_0006 ? TestBlock__B_op94 : array_index_71960[6];
  assign array_update_71963[7] = add_71961 == 32'h0000_0007 ? TestBlock__B_op94 : array_index_71960[7];
  assign array_update_71963[8] = add_71961 == 32'h0000_0008 ? TestBlock__B_op94 : array_index_71960[8];
  assign array_update_71963[9] = add_71961 == 32'h0000_0009 ? TestBlock__B_op94 : array_index_71960[9];
  assign array_update_71964[0] = add_71915 == 32'h0000_0000 ? array_update_71962 : array_update_71954[0];
  assign array_update_71964[1] = add_71915 == 32'h0000_0001 ? array_update_71962 : array_update_71954[1];
  assign array_update_71964[2] = add_71915 == 32'h0000_0002 ? array_update_71962 : array_update_71954[2];
  assign array_update_71964[3] = add_71915 == 32'h0000_0003 ? array_update_71962 : array_update_71954[3];
  assign array_update_71964[4] = add_71915 == 32'h0000_0004 ? array_update_71962 : array_update_71954[4];
  assign array_update_71964[5] = add_71915 == 32'h0000_0005 ? array_update_71962 : array_update_71954[5];
  assign array_update_71964[6] = add_71915 == 32'h0000_0006 ? array_update_71962 : array_update_71954[6];
  assign array_update_71964[7] = add_71915 == 32'h0000_0007 ? array_update_71962 : array_update_71954[7];
  assign array_update_71964[8] = add_71915 == 32'h0000_0008 ? array_update_71962 : array_update_71954[8];
  assign array_update_71964[9] = add_71915 == 32'h0000_0009 ? array_update_71962 : array_update_71954[9];
  assign array_update_71966[0] = add_71917 == 32'h0000_0000 ? array_update_71963 : array_update_71956[0];
  assign array_update_71966[1] = add_71917 == 32'h0000_0001 ? array_update_71963 : array_update_71956[1];
  assign array_update_71966[2] = add_71917 == 32'h0000_0002 ? array_update_71963 : array_update_71956[2];
  assign array_update_71966[3] = add_71917 == 32'h0000_0003 ? array_update_71963 : array_update_71956[3];
  assign array_update_71966[4] = add_71917 == 32'h0000_0004 ? array_update_71963 : array_update_71956[4];
  assign array_update_71966[5] = add_71917 == 32'h0000_0005 ? array_update_71963 : array_update_71956[5];
  assign array_update_71966[6] = add_71917 == 32'h0000_0006 ? array_update_71963 : array_update_71956[6];
  assign array_update_71966[7] = add_71917 == 32'h0000_0007 ? array_update_71963 : array_update_71956[7];
  assign array_update_71966[8] = add_71917 == 32'h0000_0008 ? array_update_71963 : array_update_71956[8];
  assign array_update_71966[9] = add_71917 == 32'h0000_0009 ? array_update_71963 : array_update_71956[9];
  assign array_index_71968 = array_update_71964[add_71915 > 32'h0000_0009 ? 4'h9 : add_71915[3:0]];
  assign add_71969 = add_71959 + 32'h0000_0001;
  assign array_index_71970 = array_update_71966[add_71917 > 32'h0000_0009 ? 4'h9 : add_71917[3:0]];
  assign add_71971 = add_71961 + 32'h0000_0001;
  assign array_update_71972[0] = add_71969 == 32'h0000_0000 ? TestBlock__A_op95 : array_index_71968[0];
  assign array_update_71972[1] = add_71969 == 32'h0000_0001 ? TestBlock__A_op95 : array_index_71968[1];
  assign array_update_71972[2] = add_71969 == 32'h0000_0002 ? TestBlock__A_op95 : array_index_71968[2];
  assign array_update_71972[3] = add_71969 == 32'h0000_0003 ? TestBlock__A_op95 : array_index_71968[3];
  assign array_update_71972[4] = add_71969 == 32'h0000_0004 ? TestBlock__A_op95 : array_index_71968[4];
  assign array_update_71972[5] = add_71969 == 32'h0000_0005 ? TestBlock__A_op95 : array_index_71968[5];
  assign array_update_71972[6] = add_71969 == 32'h0000_0006 ? TestBlock__A_op95 : array_index_71968[6];
  assign array_update_71972[7] = add_71969 == 32'h0000_0007 ? TestBlock__A_op95 : array_index_71968[7];
  assign array_update_71972[8] = add_71969 == 32'h0000_0008 ? TestBlock__A_op95 : array_index_71968[8];
  assign array_update_71972[9] = add_71969 == 32'h0000_0009 ? TestBlock__A_op95 : array_index_71968[9];
  assign array_update_71973[0] = add_71971 == 32'h0000_0000 ? TestBlock__B_op95 : array_index_71970[0];
  assign array_update_71973[1] = add_71971 == 32'h0000_0001 ? TestBlock__B_op95 : array_index_71970[1];
  assign array_update_71973[2] = add_71971 == 32'h0000_0002 ? TestBlock__B_op95 : array_index_71970[2];
  assign array_update_71973[3] = add_71971 == 32'h0000_0003 ? TestBlock__B_op95 : array_index_71970[3];
  assign array_update_71973[4] = add_71971 == 32'h0000_0004 ? TestBlock__B_op95 : array_index_71970[4];
  assign array_update_71973[5] = add_71971 == 32'h0000_0005 ? TestBlock__B_op95 : array_index_71970[5];
  assign array_update_71973[6] = add_71971 == 32'h0000_0006 ? TestBlock__B_op95 : array_index_71970[6];
  assign array_update_71973[7] = add_71971 == 32'h0000_0007 ? TestBlock__B_op95 : array_index_71970[7];
  assign array_update_71973[8] = add_71971 == 32'h0000_0008 ? TestBlock__B_op95 : array_index_71970[8];
  assign array_update_71973[9] = add_71971 == 32'h0000_0009 ? TestBlock__B_op95 : array_index_71970[9];
  assign array_update_71974[0] = add_71915 == 32'h0000_0000 ? array_update_71972 : array_update_71964[0];
  assign array_update_71974[1] = add_71915 == 32'h0000_0001 ? array_update_71972 : array_update_71964[1];
  assign array_update_71974[2] = add_71915 == 32'h0000_0002 ? array_update_71972 : array_update_71964[2];
  assign array_update_71974[3] = add_71915 == 32'h0000_0003 ? array_update_71972 : array_update_71964[3];
  assign array_update_71974[4] = add_71915 == 32'h0000_0004 ? array_update_71972 : array_update_71964[4];
  assign array_update_71974[5] = add_71915 == 32'h0000_0005 ? array_update_71972 : array_update_71964[5];
  assign array_update_71974[6] = add_71915 == 32'h0000_0006 ? array_update_71972 : array_update_71964[6];
  assign array_update_71974[7] = add_71915 == 32'h0000_0007 ? array_update_71972 : array_update_71964[7];
  assign array_update_71974[8] = add_71915 == 32'h0000_0008 ? array_update_71972 : array_update_71964[8];
  assign array_update_71974[9] = add_71915 == 32'h0000_0009 ? array_update_71972 : array_update_71964[9];
  assign array_update_71976[0] = add_71917 == 32'h0000_0000 ? array_update_71973 : array_update_71966[0];
  assign array_update_71976[1] = add_71917 == 32'h0000_0001 ? array_update_71973 : array_update_71966[1];
  assign array_update_71976[2] = add_71917 == 32'h0000_0002 ? array_update_71973 : array_update_71966[2];
  assign array_update_71976[3] = add_71917 == 32'h0000_0003 ? array_update_71973 : array_update_71966[3];
  assign array_update_71976[4] = add_71917 == 32'h0000_0004 ? array_update_71973 : array_update_71966[4];
  assign array_update_71976[5] = add_71917 == 32'h0000_0005 ? array_update_71973 : array_update_71966[5];
  assign array_update_71976[6] = add_71917 == 32'h0000_0006 ? array_update_71973 : array_update_71966[6];
  assign array_update_71976[7] = add_71917 == 32'h0000_0007 ? array_update_71973 : array_update_71966[7];
  assign array_update_71976[8] = add_71917 == 32'h0000_0008 ? array_update_71973 : array_update_71966[8];
  assign array_update_71976[9] = add_71917 == 32'h0000_0009 ? array_update_71973 : array_update_71966[9];
  assign array_index_71978 = array_update_71974[add_71915 > 32'h0000_0009 ? 4'h9 : add_71915[3:0]];
  assign add_71979 = add_71969 + 32'h0000_0001;
  assign array_index_71980 = array_update_71976[add_71917 > 32'h0000_0009 ? 4'h9 : add_71917[3:0]];
  assign add_71981 = add_71971 + 32'h0000_0001;
  assign array_update_71982[0] = add_71979 == 32'h0000_0000 ? TestBlock__A_op96 : array_index_71978[0];
  assign array_update_71982[1] = add_71979 == 32'h0000_0001 ? TestBlock__A_op96 : array_index_71978[1];
  assign array_update_71982[2] = add_71979 == 32'h0000_0002 ? TestBlock__A_op96 : array_index_71978[2];
  assign array_update_71982[3] = add_71979 == 32'h0000_0003 ? TestBlock__A_op96 : array_index_71978[3];
  assign array_update_71982[4] = add_71979 == 32'h0000_0004 ? TestBlock__A_op96 : array_index_71978[4];
  assign array_update_71982[5] = add_71979 == 32'h0000_0005 ? TestBlock__A_op96 : array_index_71978[5];
  assign array_update_71982[6] = add_71979 == 32'h0000_0006 ? TestBlock__A_op96 : array_index_71978[6];
  assign array_update_71982[7] = add_71979 == 32'h0000_0007 ? TestBlock__A_op96 : array_index_71978[7];
  assign array_update_71982[8] = add_71979 == 32'h0000_0008 ? TestBlock__A_op96 : array_index_71978[8];
  assign array_update_71982[9] = add_71979 == 32'h0000_0009 ? TestBlock__A_op96 : array_index_71978[9];
  assign array_update_71983[0] = add_71981 == 32'h0000_0000 ? TestBlock__B_op96 : array_index_71980[0];
  assign array_update_71983[1] = add_71981 == 32'h0000_0001 ? TestBlock__B_op96 : array_index_71980[1];
  assign array_update_71983[2] = add_71981 == 32'h0000_0002 ? TestBlock__B_op96 : array_index_71980[2];
  assign array_update_71983[3] = add_71981 == 32'h0000_0003 ? TestBlock__B_op96 : array_index_71980[3];
  assign array_update_71983[4] = add_71981 == 32'h0000_0004 ? TestBlock__B_op96 : array_index_71980[4];
  assign array_update_71983[5] = add_71981 == 32'h0000_0005 ? TestBlock__B_op96 : array_index_71980[5];
  assign array_update_71983[6] = add_71981 == 32'h0000_0006 ? TestBlock__B_op96 : array_index_71980[6];
  assign array_update_71983[7] = add_71981 == 32'h0000_0007 ? TestBlock__B_op96 : array_index_71980[7];
  assign array_update_71983[8] = add_71981 == 32'h0000_0008 ? TestBlock__B_op96 : array_index_71980[8];
  assign array_update_71983[9] = add_71981 == 32'h0000_0009 ? TestBlock__B_op96 : array_index_71980[9];
  assign array_update_71984[0] = add_71915 == 32'h0000_0000 ? array_update_71982 : array_update_71974[0];
  assign array_update_71984[1] = add_71915 == 32'h0000_0001 ? array_update_71982 : array_update_71974[1];
  assign array_update_71984[2] = add_71915 == 32'h0000_0002 ? array_update_71982 : array_update_71974[2];
  assign array_update_71984[3] = add_71915 == 32'h0000_0003 ? array_update_71982 : array_update_71974[3];
  assign array_update_71984[4] = add_71915 == 32'h0000_0004 ? array_update_71982 : array_update_71974[4];
  assign array_update_71984[5] = add_71915 == 32'h0000_0005 ? array_update_71982 : array_update_71974[5];
  assign array_update_71984[6] = add_71915 == 32'h0000_0006 ? array_update_71982 : array_update_71974[6];
  assign array_update_71984[7] = add_71915 == 32'h0000_0007 ? array_update_71982 : array_update_71974[7];
  assign array_update_71984[8] = add_71915 == 32'h0000_0008 ? array_update_71982 : array_update_71974[8];
  assign array_update_71984[9] = add_71915 == 32'h0000_0009 ? array_update_71982 : array_update_71974[9];
  assign array_update_71986[0] = add_71917 == 32'h0000_0000 ? array_update_71983 : array_update_71976[0];
  assign array_update_71986[1] = add_71917 == 32'h0000_0001 ? array_update_71983 : array_update_71976[1];
  assign array_update_71986[2] = add_71917 == 32'h0000_0002 ? array_update_71983 : array_update_71976[2];
  assign array_update_71986[3] = add_71917 == 32'h0000_0003 ? array_update_71983 : array_update_71976[3];
  assign array_update_71986[4] = add_71917 == 32'h0000_0004 ? array_update_71983 : array_update_71976[4];
  assign array_update_71986[5] = add_71917 == 32'h0000_0005 ? array_update_71983 : array_update_71976[5];
  assign array_update_71986[6] = add_71917 == 32'h0000_0006 ? array_update_71983 : array_update_71976[6];
  assign array_update_71986[7] = add_71917 == 32'h0000_0007 ? array_update_71983 : array_update_71976[7];
  assign array_update_71986[8] = add_71917 == 32'h0000_0008 ? array_update_71983 : array_update_71976[8];
  assign array_update_71986[9] = add_71917 == 32'h0000_0009 ? array_update_71983 : array_update_71976[9];
  assign array_index_71988 = array_update_71984[add_71915 > 32'h0000_0009 ? 4'h9 : add_71915[3:0]];
  assign add_71989 = add_71979 + 32'h0000_0001;
  assign array_index_71990 = array_update_71986[add_71917 > 32'h0000_0009 ? 4'h9 : add_71917[3:0]];
  assign add_71991 = add_71981 + 32'h0000_0001;
  assign array_update_71992[0] = add_71989 == 32'h0000_0000 ? TestBlock__A_op97 : array_index_71988[0];
  assign array_update_71992[1] = add_71989 == 32'h0000_0001 ? TestBlock__A_op97 : array_index_71988[1];
  assign array_update_71992[2] = add_71989 == 32'h0000_0002 ? TestBlock__A_op97 : array_index_71988[2];
  assign array_update_71992[3] = add_71989 == 32'h0000_0003 ? TestBlock__A_op97 : array_index_71988[3];
  assign array_update_71992[4] = add_71989 == 32'h0000_0004 ? TestBlock__A_op97 : array_index_71988[4];
  assign array_update_71992[5] = add_71989 == 32'h0000_0005 ? TestBlock__A_op97 : array_index_71988[5];
  assign array_update_71992[6] = add_71989 == 32'h0000_0006 ? TestBlock__A_op97 : array_index_71988[6];
  assign array_update_71992[7] = add_71989 == 32'h0000_0007 ? TestBlock__A_op97 : array_index_71988[7];
  assign array_update_71992[8] = add_71989 == 32'h0000_0008 ? TestBlock__A_op97 : array_index_71988[8];
  assign array_update_71992[9] = add_71989 == 32'h0000_0009 ? TestBlock__A_op97 : array_index_71988[9];
  assign array_update_71993[0] = add_71991 == 32'h0000_0000 ? TestBlock__B_op97 : array_index_71990[0];
  assign array_update_71993[1] = add_71991 == 32'h0000_0001 ? TestBlock__B_op97 : array_index_71990[1];
  assign array_update_71993[2] = add_71991 == 32'h0000_0002 ? TestBlock__B_op97 : array_index_71990[2];
  assign array_update_71993[3] = add_71991 == 32'h0000_0003 ? TestBlock__B_op97 : array_index_71990[3];
  assign array_update_71993[4] = add_71991 == 32'h0000_0004 ? TestBlock__B_op97 : array_index_71990[4];
  assign array_update_71993[5] = add_71991 == 32'h0000_0005 ? TestBlock__B_op97 : array_index_71990[5];
  assign array_update_71993[6] = add_71991 == 32'h0000_0006 ? TestBlock__B_op97 : array_index_71990[6];
  assign array_update_71993[7] = add_71991 == 32'h0000_0007 ? TestBlock__B_op97 : array_index_71990[7];
  assign array_update_71993[8] = add_71991 == 32'h0000_0008 ? TestBlock__B_op97 : array_index_71990[8];
  assign array_update_71993[9] = add_71991 == 32'h0000_0009 ? TestBlock__B_op97 : array_index_71990[9];
  assign array_update_71994[0] = add_71915 == 32'h0000_0000 ? array_update_71992 : array_update_71984[0];
  assign array_update_71994[1] = add_71915 == 32'h0000_0001 ? array_update_71992 : array_update_71984[1];
  assign array_update_71994[2] = add_71915 == 32'h0000_0002 ? array_update_71992 : array_update_71984[2];
  assign array_update_71994[3] = add_71915 == 32'h0000_0003 ? array_update_71992 : array_update_71984[3];
  assign array_update_71994[4] = add_71915 == 32'h0000_0004 ? array_update_71992 : array_update_71984[4];
  assign array_update_71994[5] = add_71915 == 32'h0000_0005 ? array_update_71992 : array_update_71984[5];
  assign array_update_71994[6] = add_71915 == 32'h0000_0006 ? array_update_71992 : array_update_71984[6];
  assign array_update_71994[7] = add_71915 == 32'h0000_0007 ? array_update_71992 : array_update_71984[7];
  assign array_update_71994[8] = add_71915 == 32'h0000_0008 ? array_update_71992 : array_update_71984[8];
  assign array_update_71994[9] = add_71915 == 32'h0000_0009 ? array_update_71992 : array_update_71984[9];
  assign array_update_71996[0] = add_71917 == 32'h0000_0000 ? array_update_71993 : array_update_71986[0];
  assign array_update_71996[1] = add_71917 == 32'h0000_0001 ? array_update_71993 : array_update_71986[1];
  assign array_update_71996[2] = add_71917 == 32'h0000_0002 ? array_update_71993 : array_update_71986[2];
  assign array_update_71996[3] = add_71917 == 32'h0000_0003 ? array_update_71993 : array_update_71986[3];
  assign array_update_71996[4] = add_71917 == 32'h0000_0004 ? array_update_71993 : array_update_71986[4];
  assign array_update_71996[5] = add_71917 == 32'h0000_0005 ? array_update_71993 : array_update_71986[5];
  assign array_update_71996[6] = add_71917 == 32'h0000_0006 ? array_update_71993 : array_update_71986[6];
  assign array_update_71996[7] = add_71917 == 32'h0000_0007 ? array_update_71993 : array_update_71986[7];
  assign array_update_71996[8] = add_71917 == 32'h0000_0008 ? array_update_71993 : array_update_71986[8];
  assign array_update_71996[9] = add_71917 == 32'h0000_0009 ? array_update_71993 : array_update_71986[9];
  assign array_index_71998 = array_update_71994[add_71915 > 32'h0000_0009 ? 4'h9 : add_71915[3:0]];
  assign add_71999 = add_71989 + 32'h0000_0001;
  assign array_index_72000 = array_update_71996[add_71917 > 32'h0000_0009 ? 4'h9 : add_71917[3:0]];
  assign add_72001 = add_71991 + 32'h0000_0001;
  assign array_update_72002[0] = add_71999 == 32'h0000_0000 ? TestBlock__A_op98 : array_index_71998[0];
  assign array_update_72002[1] = add_71999 == 32'h0000_0001 ? TestBlock__A_op98 : array_index_71998[1];
  assign array_update_72002[2] = add_71999 == 32'h0000_0002 ? TestBlock__A_op98 : array_index_71998[2];
  assign array_update_72002[3] = add_71999 == 32'h0000_0003 ? TestBlock__A_op98 : array_index_71998[3];
  assign array_update_72002[4] = add_71999 == 32'h0000_0004 ? TestBlock__A_op98 : array_index_71998[4];
  assign array_update_72002[5] = add_71999 == 32'h0000_0005 ? TestBlock__A_op98 : array_index_71998[5];
  assign array_update_72002[6] = add_71999 == 32'h0000_0006 ? TestBlock__A_op98 : array_index_71998[6];
  assign array_update_72002[7] = add_71999 == 32'h0000_0007 ? TestBlock__A_op98 : array_index_71998[7];
  assign array_update_72002[8] = add_71999 == 32'h0000_0008 ? TestBlock__A_op98 : array_index_71998[8];
  assign array_update_72002[9] = add_71999 == 32'h0000_0009 ? TestBlock__A_op98 : array_index_71998[9];
  assign array_update_72003[0] = add_72001 == 32'h0000_0000 ? TestBlock__B_op98 : array_index_72000[0];
  assign array_update_72003[1] = add_72001 == 32'h0000_0001 ? TestBlock__B_op98 : array_index_72000[1];
  assign array_update_72003[2] = add_72001 == 32'h0000_0002 ? TestBlock__B_op98 : array_index_72000[2];
  assign array_update_72003[3] = add_72001 == 32'h0000_0003 ? TestBlock__B_op98 : array_index_72000[3];
  assign array_update_72003[4] = add_72001 == 32'h0000_0004 ? TestBlock__B_op98 : array_index_72000[4];
  assign array_update_72003[5] = add_72001 == 32'h0000_0005 ? TestBlock__B_op98 : array_index_72000[5];
  assign array_update_72003[6] = add_72001 == 32'h0000_0006 ? TestBlock__B_op98 : array_index_72000[6];
  assign array_update_72003[7] = add_72001 == 32'h0000_0007 ? TestBlock__B_op98 : array_index_72000[7];
  assign array_update_72003[8] = add_72001 == 32'h0000_0008 ? TestBlock__B_op98 : array_index_72000[8];
  assign array_update_72003[9] = add_72001 == 32'h0000_0009 ? TestBlock__B_op98 : array_index_72000[9];
  assign array_update_72004[0] = add_71915 == 32'h0000_0000 ? array_update_72002 : array_update_71994[0];
  assign array_update_72004[1] = add_71915 == 32'h0000_0001 ? array_update_72002 : array_update_71994[1];
  assign array_update_72004[2] = add_71915 == 32'h0000_0002 ? array_update_72002 : array_update_71994[2];
  assign array_update_72004[3] = add_71915 == 32'h0000_0003 ? array_update_72002 : array_update_71994[3];
  assign array_update_72004[4] = add_71915 == 32'h0000_0004 ? array_update_72002 : array_update_71994[4];
  assign array_update_72004[5] = add_71915 == 32'h0000_0005 ? array_update_72002 : array_update_71994[5];
  assign array_update_72004[6] = add_71915 == 32'h0000_0006 ? array_update_72002 : array_update_71994[6];
  assign array_update_72004[7] = add_71915 == 32'h0000_0007 ? array_update_72002 : array_update_71994[7];
  assign array_update_72004[8] = add_71915 == 32'h0000_0008 ? array_update_72002 : array_update_71994[8];
  assign array_update_72004[9] = add_71915 == 32'h0000_0009 ? array_update_72002 : array_update_71994[9];
  assign array_update_72006[0] = add_71917 == 32'h0000_0000 ? array_update_72003 : array_update_71996[0];
  assign array_update_72006[1] = add_71917 == 32'h0000_0001 ? array_update_72003 : array_update_71996[1];
  assign array_update_72006[2] = add_71917 == 32'h0000_0002 ? array_update_72003 : array_update_71996[2];
  assign array_update_72006[3] = add_71917 == 32'h0000_0003 ? array_update_72003 : array_update_71996[3];
  assign array_update_72006[4] = add_71917 == 32'h0000_0004 ? array_update_72003 : array_update_71996[4];
  assign array_update_72006[5] = add_71917 == 32'h0000_0005 ? array_update_72003 : array_update_71996[5];
  assign array_update_72006[6] = add_71917 == 32'h0000_0006 ? array_update_72003 : array_update_71996[6];
  assign array_update_72006[7] = add_71917 == 32'h0000_0007 ? array_update_72003 : array_update_71996[7];
  assign array_update_72006[8] = add_71917 == 32'h0000_0008 ? array_update_72003 : array_update_71996[8];
  assign array_update_72006[9] = add_71917 == 32'h0000_0009 ? array_update_72003 : array_update_71996[9];
  assign literal_72009 = 32'h0000_0000;
  assign array_index_72010 = array_update_72004[add_71915 > 32'h0000_0009 ? 4'h9 : add_71915[3:0]];
  assign add_72011 = add_71999 + 32'h0000_0001;
  assign array_index_72012 = array_update_72006[add_71917 > 32'h0000_0009 ? 4'h9 : add_71917[3:0]];
  assign add_72013 = add_72001 + 32'h0000_0001;
  assign array_index_72014 = literal_72008[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign literal_72016 = 32'h0000_0000;
  assign array_update_72017[0] = add_72011 == 32'h0000_0000 ? TestBlock__A_op99 : array_index_72010[0];
  assign array_update_72017[1] = add_72011 == 32'h0000_0001 ? TestBlock__A_op99 : array_index_72010[1];
  assign array_update_72017[2] = add_72011 == 32'h0000_0002 ? TestBlock__A_op99 : array_index_72010[2];
  assign array_update_72017[3] = add_72011 == 32'h0000_0003 ? TestBlock__A_op99 : array_index_72010[3];
  assign array_update_72017[4] = add_72011 == 32'h0000_0004 ? TestBlock__A_op99 : array_index_72010[4];
  assign array_update_72017[5] = add_72011 == 32'h0000_0005 ? TestBlock__A_op99 : array_index_72010[5];
  assign array_update_72017[6] = add_72011 == 32'h0000_0006 ? TestBlock__A_op99 : array_index_72010[6];
  assign array_update_72017[7] = add_72011 == 32'h0000_0007 ? TestBlock__A_op99 : array_index_72010[7];
  assign array_update_72017[8] = add_72011 == 32'h0000_0008 ? TestBlock__A_op99 : array_index_72010[8];
  assign array_update_72017[9] = add_72011 == 32'h0000_0009 ? TestBlock__A_op99 : array_index_72010[9];
  assign array_update_72018[0] = add_72013 == 32'h0000_0000 ? TestBlock__B_op99 : array_index_72012[0];
  assign array_update_72018[1] = add_72013 == 32'h0000_0001 ? TestBlock__B_op99 : array_index_72012[1];
  assign array_update_72018[2] = add_72013 == 32'h0000_0002 ? TestBlock__B_op99 : array_index_72012[2];
  assign array_update_72018[3] = add_72013 == 32'h0000_0003 ? TestBlock__B_op99 : array_index_72012[3];
  assign array_update_72018[4] = add_72013 == 32'h0000_0004 ? TestBlock__B_op99 : array_index_72012[4];
  assign array_update_72018[5] = add_72013 == 32'h0000_0005 ? TestBlock__B_op99 : array_index_72012[5];
  assign array_update_72018[6] = add_72013 == 32'h0000_0006 ? TestBlock__B_op99 : array_index_72012[6];
  assign array_update_72018[7] = add_72013 == 32'h0000_0007 ? TestBlock__B_op99 : array_index_72012[7];
  assign array_update_72018[8] = add_72013 == 32'h0000_0008 ? TestBlock__B_op99 : array_index_72012[8];
  assign array_update_72018[9] = add_72013 == 32'h0000_0009 ? TestBlock__B_op99 : array_index_72012[9];
  assign array_update_72019[0] = literal_72016 == 32'h0000_0000 ? 32'h0000_0000 : array_index_72014[0];
  assign array_update_72019[1] = literal_72016 == 32'h0000_0001 ? 32'h0000_0000 : array_index_72014[1];
  assign array_update_72019[2] = literal_72016 == 32'h0000_0002 ? 32'h0000_0000 : array_index_72014[2];
  assign array_update_72019[3] = literal_72016 == 32'h0000_0003 ? 32'h0000_0000 : array_index_72014[3];
  assign array_update_72019[4] = literal_72016 == 32'h0000_0004 ? 32'h0000_0000 : array_index_72014[4];
  assign array_update_72019[5] = literal_72016 == 32'h0000_0005 ? 32'h0000_0000 : array_index_72014[5];
  assign array_update_72019[6] = literal_72016 == 32'h0000_0006 ? 32'h0000_0000 : array_index_72014[6];
  assign array_update_72019[7] = literal_72016 == 32'h0000_0007 ? 32'h0000_0000 : array_index_72014[7];
  assign array_update_72019[8] = literal_72016 == 32'h0000_0008 ? 32'h0000_0000 : array_index_72014[8];
  assign array_update_72019[9] = literal_72016 == 32'h0000_0009 ? 32'h0000_0000 : array_index_72014[9];
  assign array_update_72020[0] = add_71915 == 32'h0000_0000 ? array_update_72017 : array_update_72004[0];
  assign array_update_72020[1] = add_71915 == 32'h0000_0001 ? array_update_72017 : array_update_72004[1];
  assign array_update_72020[2] = add_71915 == 32'h0000_0002 ? array_update_72017 : array_update_72004[2];
  assign array_update_72020[3] = add_71915 == 32'h0000_0003 ? array_update_72017 : array_update_72004[3];
  assign array_update_72020[4] = add_71915 == 32'h0000_0004 ? array_update_72017 : array_update_72004[4];
  assign array_update_72020[5] = add_71915 == 32'h0000_0005 ? array_update_72017 : array_update_72004[5];
  assign array_update_72020[6] = add_71915 == 32'h0000_0006 ? array_update_72017 : array_update_72004[6];
  assign array_update_72020[7] = add_71915 == 32'h0000_0007 ? array_update_72017 : array_update_72004[7];
  assign array_update_72020[8] = add_71915 == 32'h0000_0008 ? array_update_72017 : array_update_72004[8];
  assign array_update_72020[9] = add_71915 == 32'h0000_0009 ? array_update_72017 : array_update_72004[9];
  assign array_update_72021[0] = add_71917 == 32'h0000_0000 ? array_update_72018 : array_update_72006[0];
  assign array_update_72021[1] = add_71917 == 32'h0000_0001 ? array_update_72018 : array_update_72006[1];
  assign array_update_72021[2] = add_71917 == 32'h0000_0002 ? array_update_72018 : array_update_72006[2];
  assign array_update_72021[3] = add_71917 == 32'h0000_0003 ? array_update_72018 : array_update_72006[3];
  assign array_update_72021[4] = add_71917 == 32'h0000_0004 ? array_update_72018 : array_update_72006[4];
  assign array_update_72021[5] = add_71917 == 32'h0000_0005 ? array_update_72018 : array_update_72006[5];
  assign array_update_72021[6] = add_71917 == 32'h0000_0006 ? array_update_72018 : array_update_72006[6];
  assign array_update_72021[7] = add_71917 == 32'h0000_0007 ? array_update_72018 : array_update_72006[7];
  assign array_update_72021[8] = add_71917 == 32'h0000_0008 ? array_update_72018 : array_update_72006[8];
  assign array_update_72021[9] = add_71917 == 32'h0000_0009 ? array_update_72018 : array_update_72006[9];
  assign literal_72022 = 32'h0000_0000;
  assign array_update_72023[0] = literal_72009 == 32'h0000_0000 ? array_update_72019 : literal_72008[0];
  assign array_update_72023[1] = literal_72009 == 32'h0000_0001 ? array_update_72019 : literal_72008[1];
  assign array_update_72023[2] = literal_72009 == 32'h0000_0002 ? array_update_72019 : literal_72008[2];
  assign array_update_72023[3] = literal_72009 == 32'h0000_0003 ? array_update_72019 : literal_72008[3];
  assign array_update_72023[4] = literal_72009 == 32'h0000_0004 ? array_update_72019 : literal_72008[4];
  assign array_update_72023[5] = literal_72009 == 32'h0000_0005 ? array_update_72019 : literal_72008[5];
  assign array_update_72023[6] = literal_72009 == 32'h0000_0006 ? array_update_72019 : literal_72008[6];
  assign array_update_72023[7] = literal_72009 == 32'h0000_0007 ? array_update_72019 : literal_72008[7];
  assign array_update_72023[8] = literal_72009 == 32'h0000_0008 ? array_update_72019 : literal_72008[8];
  assign array_update_72023[9] = literal_72009 == 32'h0000_0009 ? array_update_72019 : literal_72008[9];
  assign array_index_72024 = array_update_72020[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign array_index_72025 = array_update_72021[literal_72022 > 32'h0000_0009 ? 4'h9 : literal_72022[3:0]];
  assign array_index_72026 = array_update_72023[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_72030 = smul32b_32b_x_32b(array_index_72024[literal_72022 > 32'h0000_0009 ? 4'h9 : literal_72022[3:0]], array_index_72025[literal_72016 > 32'h0000_0009 ? 4'h9 : literal_72016[3:0]]);
  assign add_72032 = array_index_72026[literal_72016 > 32'h0000_0009 ? 4'h9 : literal_72016[3:0]] + smul_72030;
  assign array_update_72034[0] = literal_72016 == 32'h0000_0000 ? add_72032 : array_index_72026[0];
  assign array_update_72034[1] = literal_72016 == 32'h0000_0001 ? add_72032 : array_index_72026[1];
  assign array_update_72034[2] = literal_72016 == 32'h0000_0002 ? add_72032 : array_index_72026[2];
  assign array_update_72034[3] = literal_72016 == 32'h0000_0003 ? add_72032 : array_index_72026[3];
  assign array_update_72034[4] = literal_72016 == 32'h0000_0004 ? add_72032 : array_index_72026[4];
  assign array_update_72034[5] = literal_72016 == 32'h0000_0005 ? add_72032 : array_index_72026[5];
  assign array_update_72034[6] = literal_72016 == 32'h0000_0006 ? add_72032 : array_index_72026[6];
  assign array_update_72034[7] = literal_72016 == 32'h0000_0007 ? add_72032 : array_index_72026[7];
  assign array_update_72034[8] = literal_72016 == 32'h0000_0008 ? add_72032 : array_index_72026[8];
  assign array_update_72034[9] = literal_72016 == 32'h0000_0009 ? add_72032 : array_index_72026[9];
  assign add_72035 = literal_72022 + 32'h0000_0001;
  assign array_update_72036[0] = literal_72009 == 32'h0000_0000 ? array_update_72034 : array_update_72023[0];
  assign array_update_72036[1] = literal_72009 == 32'h0000_0001 ? array_update_72034 : array_update_72023[1];
  assign array_update_72036[2] = literal_72009 == 32'h0000_0002 ? array_update_72034 : array_update_72023[2];
  assign array_update_72036[3] = literal_72009 == 32'h0000_0003 ? array_update_72034 : array_update_72023[3];
  assign array_update_72036[4] = literal_72009 == 32'h0000_0004 ? array_update_72034 : array_update_72023[4];
  assign array_update_72036[5] = literal_72009 == 32'h0000_0005 ? array_update_72034 : array_update_72023[5];
  assign array_update_72036[6] = literal_72009 == 32'h0000_0006 ? array_update_72034 : array_update_72023[6];
  assign array_update_72036[7] = literal_72009 == 32'h0000_0007 ? array_update_72034 : array_update_72023[7];
  assign array_update_72036[8] = literal_72009 == 32'h0000_0008 ? array_update_72034 : array_update_72023[8];
  assign array_update_72036[9] = literal_72009 == 32'h0000_0009 ? array_update_72034 : array_update_72023[9];
  assign array_index_72038 = array_update_72021[add_72035 > 32'h0000_0009 ? 4'h9 : add_72035[3:0]];
  assign array_index_72039 = array_update_72036[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_72043 = smul32b_32b_x_32b(array_index_72024[add_72035 > 32'h0000_0009 ? 4'h9 : add_72035[3:0]], array_index_72038[literal_72016 > 32'h0000_0009 ? 4'h9 : literal_72016[3:0]]);
  assign add_72045 = array_index_72039[literal_72016 > 32'h0000_0009 ? 4'h9 : literal_72016[3:0]] + smul_72043;
  assign array_update_72047[0] = literal_72016 == 32'h0000_0000 ? add_72045 : array_index_72039[0];
  assign array_update_72047[1] = literal_72016 == 32'h0000_0001 ? add_72045 : array_index_72039[1];
  assign array_update_72047[2] = literal_72016 == 32'h0000_0002 ? add_72045 : array_index_72039[2];
  assign array_update_72047[3] = literal_72016 == 32'h0000_0003 ? add_72045 : array_index_72039[3];
  assign array_update_72047[4] = literal_72016 == 32'h0000_0004 ? add_72045 : array_index_72039[4];
  assign array_update_72047[5] = literal_72016 == 32'h0000_0005 ? add_72045 : array_index_72039[5];
  assign array_update_72047[6] = literal_72016 == 32'h0000_0006 ? add_72045 : array_index_72039[6];
  assign array_update_72047[7] = literal_72016 == 32'h0000_0007 ? add_72045 : array_index_72039[7];
  assign array_update_72047[8] = literal_72016 == 32'h0000_0008 ? add_72045 : array_index_72039[8];
  assign array_update_72047[9] = literal_72016 == 32'h0000_0009 ? add_72045 : array_index_72039[9];
  assign add_72048 = add_72035 + 32'h0000_0001;
  assign array_update_72049[0] = literal_72009 == 32'h0000_0000 ? array_update_72047 : array_update_72036[0];
  assign array_update_72049[1] = literal_72009 == 32'h0000_0001 ? array_update_72047 : array_update_72036[1];
  assign array_update_72049[2] = literal_72009 == 32'h0000_0002 ? array_update_72047 : array_update_72036[2];
  assign array_update_72049[3] = literal_72009 == 32'h0000_0003 ? array_update_72047 : array_update_72036[3];
  assign array_update_72049[4] = literal_72009 == 32'h0000_0004 ? array_update_72047 : array_update_72036[4];
  assign array_update_72049[5] = literal_72009 == 32'h0000_0005 ? array_update_72047 : array_update_72036[5];
  assign array_update_72049[6] = literal_72009 == 32'h0000_0006 ? array_update_72047 : array_update_72036[6];
  assign array_update_72049[7] = literal_72009 == 32'h0000_0007 ? array_update_72047 : array_update_72036[7];
  assign array_update_72049[8] = literal_72009 == 32'h0000_0008 ? array_update_72047 : array_update_72036[8];
  assign array_update_72049[9] = literal_72009 == 32'h0000_0009 ? array_update_72047 : array_update_72036[9];
  assign array_index_72051 = array_update_72021[add_72048 > 32'h0000_0009 ? 4'h9 : add_72048[3:0]];
  assign array_index_72052 = array_update_72049[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_72056 = smul32b_32b_x_32b(array_index_72024[add_72048 > 32'h0000_0009 ? 4'h9 : add_72048[3:0]], array_index_72051[literal_72016 > 32'h0000_0009 ? 4'h9 : literal_72016[3:0]]);
  assign add_72058 = array_index_72052[literal_72016 > 32'h0000_0009 ? 4'h9 : literal_72016[3:0]] + smul_72056;
  assign array_update_72060[0] = literal_72016 == 32'h0000_0000 ? add_72058 : array_index_72052[0];
  assign array_update_72060[1] = literal_72016 == 32'h0000_0001 ? add_72058 : array_index_72052[1];
  assign array_update_72060[2] = literal_72016 == 32'h0000_0002 ? add_72058 : array_index_72052[2];
  assign array_update_72060[3] = literal_72016 == 32'h0000_0003 ? add_72058 : array_index_72052[3];
  assign array_update_72060[4] = literal_72016 == 32'h0000_0004 ? add_72058 : array_index_72052[4];
  assign array_update_72060[5] = literal_72016 == 32'h0000_0005 ? add_72058 : array_index_72052[5];
  assign array_update_72060[6] = literal_72016 == 32'h0000_0006 ? add_72058 : array_index_72052[6];
  assign array_update_72060[7] = literal_72016 == 32'h0000_0007 ? add_72058 : array_index_72052[7];
  assign array_update_72060[8] = literal_72016 == 32'h0000_0008 ? add_72058 : array_index_72052[8];
  assign array_update_72060[9] = literal_72016 == 32'h0000_0009 ? add_72058 : array_index_72052[9];
  assign add_72061 = add_72048 + 32'h0000_0001;
  assign array_update_72062[0] = literal_72009 == 32'h0000_0000 ? array_update_72060 : array_update_72049[0];
  assign array_update_72062[1] = literal_72009 == 32'h0000_0001 ? array_update_72060 : array_update_72049[1];
  assign array_update_72062[2] = literal_72009 == 32'h0000_0002 ? array_update_72060 : array_update_72049[2];
  assign array_update_72062[3] = literal_72009 == 32'h0000_0003 ? array_update_72060 : array_update_72049[3];
  assign array_update_72062[4] = literal_72009 == 32'h0000_0004 ? array_update_72060 : array_update_72049[4];
  assign array_update_72062[5] = literal_72009 == 32'h0000_0005 ? array_update_72060 : array_update_72049[5];
  assign array_update_72062[6] = literal_72009 == 32'h0000_0006 ? array_update_72060 : array_update_72049[6];
  assign array_update_72062[7] = literal_72009 == 32'h0000_0007 ? array_update_72060 : array_update_72049[7];
  assign array_update_72062[8] = literal_72009 == 32'h0000_0008 ? array_update_72060 : array_update_72049[8];
  assign array_update_72062[9] = literal_72009 == 32'h0000_0009 ? array_update_72060 : array_update_72049[9];
  assign array_index_72064 = array_update_72021[add_72061 > 32'h0000_0009 ? 4'h9 : add_72061[3:0]];
  assign array_index_72065 = array_update_72062[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_72069 = smul32b_32b_x_32b(array_index_72024[add_72061 > 32'h0000_0009 ? 4'h9 : add_72061[3:0]], array_index_72064[literal_72016 > 32'h0000_0009 ? 4'h9 : literal_72016[3:0]]);
  assign add_72071 = array_index_72065[literal_72016 > 32'h0000_0009 ? 4'h9 : literal_72016[3:0]] + smul_72069;
  assign array_update_72073[0] = literal_72016 == 32'h0000_0000 ? add_72071 : array_index_72065[0];
  assign array_update_72073[1] = literal_72016 == 32'h0000_0001 ? add_72071 : array_index_72065[1];
  assign array_update_72073[2] = literal_72016 == 32'h0000_0002 ? add_72071 : array_index_72065[2];
  assign array_update_72073[3] = literal_72016 == 32'h0000_0003 ? add_72071 : array_index_72065[3];
  assign array_update_72073[4] = literal_72016 == 32'h0000_0004 ? add_72071 : array_index_72065[4];
  assign array_update_72073[5] = literal_72016 == 32'h0000_0005 ? add_72071 : array_index_72065[5];
  assign array_update_72073[6] = literal_72016 == 32'h0000_0006 ? add_72071 : array_index_72065[6];
  assign array_update_72073[7] = literal_72016 == 32'h0000_0007 ? add_72071 : array_index_72065[7];
  assign array_update_72073[8] = literal_72016 == 32'h0000_0008 ? add_72071 : array_index_72065[8];
  assign array_update_72073[9] = literal_72016 == 32'h0000_0009 ? add_72071 : array_index_72065[9];
  assign add_72074 = add_72061 + 32'h0000_0001;
  assign array_update_72075[0] = literal_72009 == 32'h0000_0000 ? array_update_72073 : array_update_72062[0];
  assign array_update_72075[1] = literal_72009 == 32'h0000_0001 ? array_update_72073 : array_update_72062[1];
  assign array_update_72075[2] = literal_72009 == 32'h0000_0002 ? array_update_72073 : array_update_72062[2];
  assign array_update_72075[3] = literal_72009 == 32'h0000_0003 ? array_update_72073 : array_update_72062[3];
  assign array_update_72075[4] = literal_72009 == 32'h0000_0004 ? array_update_72073 : array_update_72062[4];
  assign array_update_72075[5] = literal_72009 == 32'h0000_0005 ? array_update_72073 : array_update_72062[5];
  assign array_update_72075[6] = literal_72009 == 32'h0000_0006 ? array_update_72073 : array_update_72062[6];
  assign array_update_72075[7] = literal_72009 == 32'h0000_0007 ? array_update_72073 : array_update_72062[7];
  assign array_update_72075[8] = literal_72009 == 32'h0000_0008 ? array_update_72073 : array_update_72062[8];
  assign array_update_72075[9] = literal_72009 == 32'h0000_0009 ? array_update_72073 : array_update_72062[9];
  assign array_index_72077 = array_update_72021[add_72074 > 32'h0000_0009 ? 4'h9 : add_72074[3:0]];
  assign array_index_72078 = array_update_72075[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_72082 = smul32b_32b_x_32b(array_index_72024[add_72074 > 32'h0000_0009 ? 4'h9 : add_72074[3:0]], array_index_72077[literal_72016 > 32'h0000_0009 ? 4'h9 : literal_72016[3:0]]);
  assign add_72084 = array_index_72078[literal_72016 > 32'h0000_0009 ? 4'h9 : literal_72016[3:0]] + smul_72082;
  assign array_update_72086[0] = literal_72016 == 32'h0000_0000 ? add_72084 : array_index_72078[0];
  assign array_update_72086[1] = literal_72016 == 32'h0000_0001 ? add_72084 : array_index_72078[1];
  assign array_update_72086[2] = literal_72016 == 32'h0000_0002 ? add_72084 : array_index_72078[2];
  assign array_update_72086[3] = literal_72016 == 32'h0000_0003 ? add_72084 : array_index_72078[3];
  assign array_update_72086[4] = literal_72016 == 32'h0000_0004 ? add_72084 : array_index_72078[4];
  assign array_update_72086[5] = literal_72016 == 32'h0000_0005 ? add_72084 : array_index_72078[5];
  assign array_update_72086[6] = literal_72016 == 32'h0000_0006 ? add_72084 : array_index_72078[6];
  assign array_update_72086[7] = literal_72016 == 32'h0000_0007 ? add_72084 : array_index_72078[7];
  assign array_update_72086[8] = literal_72016 == 32'h0000_0008 ? add_72084 : array_index_72078[8];
  assign array_update_72086[9] = literal_72016 == 32'h0000_0009 ? add_72084 : array_index_72078[9];
  assign add_72087 = add_72074 + 32'h0000_0001;
  assign array_update_72088[0] = literal_72009 == 32'h0000_0000 ? array_update_72086 : array_update_72075[0];
  assign array_update_72088[1] = literal_72009 == 32'h0000_0001 ? array_update_72086 : array_update_72075[1];
  assign array_update_72088[2] = literal_72009 == 32'h0000_0002 ? array_update_72086 : array_update_72075[2];
  assign array_update_72088[3] = literal_72009 == 32'h0000_0003 ? array_update_72086 : array_update_72075[3];
  assign array_update_72088[4] = literal_72009 == 32'h0000_0004 ? array_update_72086 : array_update_72075[4];
  assign array_update_72088[5] = literal_72009 == 32'h0000_0005 ? array_update_72086 : array_update_72075[5];
  assign array_update_72088[6] = literal_72009 == 32'h0000_0006 ? array_update_72086 : array_update_72075[6];
  assign array_update_72088[7] = literal_72009 == 32'h0000_0007 ? array_update_72086 : array_update_72075[7];
  assign array_update_72088[8] = literal_72009 == 32'h0000_0008 ? array_update_72086 : array_update_72075[8];
  assign array_update_72088[9] = literal_72009 == 32'h0000_0009 ? array_update_72086 : array_update_72075[9];
  assign array_index_72090 = array_update_72021[add_72087 > 32'h0000_0009 ? 4'h9 : add_72087[3:0]];
  assign array_index_72091 = array_update_72088[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_72095 = smul32b_32b_x_32b(array_index_72024[add_72087 > 32'h0000_0009 ? 4'h9 : add_72087[3:0]], array_index_72090[literal_72016 > 32'h0000_0009 ? 4'h9 : literal_72016[3:0]]);
  assign add_72097 = array_index_72091[literal_72016 > 32'h0000_0009 ? 4'h9 : literal_72016[3:0]] + smul_72095;
  assign array_update_72099[0] = literal_72016 == 32'h0000_0000 ? add_72097 : array_index_72091[0];
  assign array_update_72099[1] = literal_72016 == 32'h0000_0001 ? add_72097 : array_index_72091[1];
  assign array_update_72099[2] = literal_72016 == 32'h0000_0002 ? add_72097 : array_index_72091[2];
  assign array_update_72099[3] = literal_72016 == 32'h0000_0003 ? add_72097 : array_index_72091[3];
  assign array_update_72099[4] = literal_72016 == 32'h0000_0004 ? add_72097 : array_index_72091[4];
  assign array_update_72099[5] = literal_72016 == 32'h0000_0005 ? add_72097 : array_index_72091[5];
  assign array_update_72099[6] = literal_72016 == 32'h0000_0006 ? add_72097 : array_index_72091[6];
  assign array_update_72099[7] = literal_72016 == 32'h0000_0007 ? add_72097 : array_index_72091[7];
  assign array_update_72099[8] = literal_72016 == 32'h0000_0008 ? add_72097 : array_index_72091[8];
  assign array_update_72099[9] = literal_72016 == 32'h0000_0009 ? add_72097 : array_index_72091[9];
  assign add_72100 = add_72087 + 32'h0000_0001;
  assign array_update_72101[0] = literal_72009 == 32'h0000_0000 ? array_update_72099 : array_update_72088[0];
  assign array_update_72101[1] = literal_72009 == 32'h0000_0001 ? array_update_72099 : array_update_72088[1];
  assign array_update_72101[2] = literal_72009 == 32'h0000_0002 ? array_update_72099 : array_update_72088[2];
  assign array_update_72101[3] = literal_72009 == 32'h0000_0003 ? array_update_72099 : array_update_72088[3];
  assign array_update_72101[4] = literal_72009 == 32'h0000_0004 ? array_update_72099 : array_update_72088[4];
  assign array_update_72101[5] = literal_72009 == 32'h0000_0005 ? array_update_72099 : array_update_72088[5];
  assign array_update_72101[6] = literal_72009 == 32'h0000_0006 ? array_update_72099 : array_update_72088[6];
  assign array_update_72101[7] = literal_72009 == 32'h0000_0007 ? array_update_72099 : array_update_72088[7];
  assign array_update_72101[8] = literal_72009 == 32'h0000_0008 ? array_update_72099 : array_update_72088[8];
  assign array_update_72101[9] = literal_72009 == 32'h0000_0009 ? array_update_72099 : array_update_72088[9];
  assign array_index_72103 = array_update_72021[add_72100 > 32'h0000_0009 ? 4'h9 : add_72100[3:0]];
  assign array_index_72104 = array_update_72101[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_72108 = smul32b_32b_x_32b(array_index_72024[add_72100 > 32'h0000_0009 ? 4'h9 : add_72100[3:0]], array_index_72103[literal_72016 > 32'h0000_0009 ? 4'h9 : literal_72016[3:0]]);
  assign add_72110 = array_index_72104[literal_72016 > 32'h0000_0009 ? 4'h9 : literal_72016[3:0]] + smul_72108;
  assign array_update_72112[0] = literal_72016 == 32'h0000_0000 ? add_72110 : array_index_72104[0];
  assign array_update_72112[1] = literal_72016 == 32'h0000_0001 ? add_72110 : array_index_72104[1];
  assign array_update_72112[2] = literal_72016 == 32'h0000_0002 ? add_72110 : array_index_72104[2];
  assign array_update_72112[3] = literal_72016 == 32'h0000_0003 ? add_72110 : array_index_72104[3];
  assign array_update_72112[4] = literal_72016 == 32'h0000_0004 ? add_72110 : array_index_72104[4];
  assign array_update_72112[5] = literal_72016 == 32'h0000_0005 ? add_72110 : array_index_72104[5];
  assign array_update_72112[6] = literal_72016 == 32'h0000_0006 ? add_72110 : array_index_72104[6];
  assign array_update_72112[7] = literal_72016 == 32'h0000_0007 ? add_72110 : array_index_72104[7];
  assign array_update_72112[8] = literal_72016 == 32'h0000_0008 ? add_72110 : array_index_72104[8];
  assign array_update_72112[9] = literal_72016 == 32'h0000_0009 ? add_72110 : array_index_72104[9];
  assign add_72113 = add_72100 + 32'h0000_0001;
  assign array_update_72114[0] = literal_72009 == 32'h0000_0000 ? array_update_72112 : array_update_72101[0];
  assign array_update_72114[1] = literal_72009 == 32'h0000_0001 ? array_update_72112 : array_update_72101[1];
  assign array_update_72114[2] = literal_72009 == 32'h0000_0002 ? array_update_72112 : array_update_72101[2];
  assign array_update_72114[3] = literal_72009 == 32'h0000_0003 ? array_update_72112 : array_update_72101[3];
  assign array_update_72114[4] = literal_72009 == 32'h0000_0004 ? array_update_72112 : array_update_72101[4];
  assign array_update_72114[5] = literal_72009 == 32'h0000_0005 ? array_update_72112 : array_update_72101[5];
  assign array_update_72114[6] = literal_72009 == 32'h0000_0006 ? array_update_72112 : array_update_72101[6];
  assign array_update_72114[7] = literal_72009 == 32'h0000_0007 ? array_update_72112 : array_update_72101[7];
  assign array_update_72114[8] = literal_72009 == 32'h0000_0008 ? array_update_72112 : array_update_72101[8];
  assign array_update_72114[9] = literal_72009 == 32'h0000_0009 ? array_update_72112 : array_update_72101[9];
  assign array_index_72116 = array_update_72021[add_72113 > 32'h0000_0009 ? 4'h9 : add_72113[3:0]];
  assign array_index_72117 = array_update_72114[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_72121 = smul32b_32b_x_32b(array_index_72024[add_72113 > 32'h0000_0009 ? 4'h9 : add_72113[3:0]], array_index_72116[literal_72016 > 32'h0000_0009 ? 4'h9 : literal_72016[3:0]]);
  assign add_72123 = array_index_72117[literal_72016 > 32'h0000_0009 ? 4'h9 : literal_72016[3:0]] + smul_72121;
  assign array_update_72125[0] = literal_72016 == 32'h0000_0000 ? add_72123 : array_index_72117[0];
  assign array_update_72125[1] = literal_72016 == 32'h0000_0001 ? add_72123 : array_index_72117[1];
  assign array_update_72125[2] = literal_72016 == 32'h0000_0002 ? add_72123 : array_index_72117[2];
  assign array_update_72125[3] = literal_72016 == 32'h0000_0003 ? add_72123 : array_index_72117[3];
  assign array_update_72125[4] = literal_72016 == 32'h0000_0004 ? add_72123 : array_index_72117[4];
  assign array_update_72125[5] = literal_72016 == 32'h0000_0005 ? add_72123 : array_index_72117[5];
  assign array_update_72125[6] = literal_72016 == 32'h0000_0006 ? add_72123 : array_index_72117[6];
  assign array_update_72125[7] = literal_72016 == 32'h0000_0007 ? add_72123 : array_index_72117[7];
  assign array_update_72125[8] = literal_72016 == 32'h0000_0008 ? add_72123 : array_index_72117[8];
  assign array_update_72125[9] = literal_72016 == 32'h0000_0009 ? add_72123 : array_index_72117[9];
  assign add_72126 = add_72113 + 32'h0000_0001;
  assign array_update_72127[0] = literal_72009 == 32'h0000_0000 ? array_update_72125 : array_update_72114[0];
  assign array_update_72127[1] = literal_72009 == 32'h0000_0001 ? array_update_72125 : array_update_72114[1];
  assign array_update_72127[2] = literal_72009 == 32'h0000_0002 ? array_update_72125 : array_update_72114[2];
  assign array_update_72127[3] = literal_72009 == 32'h0000_0003 ? array_update_72125 : array_update_72114[3];
  assign array_update_72127[4] = literal_72009 == 32'h0000_0004 ? array_update_72125 : array_update_72114[4];
  assign array_update_72127[5] = literal_72009 == 32'h0000_0005 ? array_update_72125 : array_update_72114[5];
  assign array_update_72127[6] = literal_72009 == 32'h0000_0006 ? array_update_72125 : array_update_72114[6];
  assign array_update_72127[7] = literal_72009 == 32'h0000_0007 ? array_update_72125 : array_update_72114[7];
  assign array_update_72127[8] = literal_72009 == 32'h0000_0008 ? array_update_72125 : array_update_72114[8];
  assign array_update_72127[9] = literal_72009 == 32'h0000_0009 ? array_update_72125 : array_update_72114[9];
  assign array_index_72129 = array_update_72021[add_72126 > 32'h0000_0009 ? 4'h9 : add_72126[3:0]];
  assign array_index_72130 = array_update_72127[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_72134 = smul32b_32b_x_32b(array_index_72024[add_72126 > 32'h0000_0009 ? 4'h9 : add_72126[3:0]], array_index_72129[literal_72016 > 32'h0000_0009 ? 4'h9 : literal_72016[3:0]]);
  assign add_72136 = array_index_72130[literal_72016 > 32'h0000_0009 ? 4'h9 : literal_72016[3:0]] + smul_72134;
  assign array_update_72138[0] = literal_72016 == 32'h0000_0000 ? add_72136 : array_index_72130[0];
  assign array_update_72138[1] = literal_72016 == 32'h0000_0001 ? add_72136 : array_index_72130[1];
  assign array_update_72138[2] = literal_72016 == 32'h0000_0002 ? add_72136 : array_index_72130[2];
  assign array_update_72138[3] = literal_72016 == 32'h0000_0003 ? add_72136 : array_index_72130[3];
  assign array_update_72138[4] = literal_72016 == 32'h0000_0004 ? add_72136 : array_index_72130[4];
  assign array_update_72138[5] = literal_72016 == 32'h0000_0005 ? add_72136 : array_index_72130[5];
  assign array_update_72138[6] = literal_72016 == 32'h0000_0006 ? add_72136 : array_index_72130[6];
  assign array_update_72138[7] = literal_72016 == 32'h0000_0007 ? add_72136 : array_index_72130[7];
  assign array_update_72138[8] = literal_72016 == 32'h0000_0008 ? add_72136 : array_index_72130[8];
  assign array_update_72138[9] = literal_72016 == 32'h0000_0009 ? add_72136 : array_index_72130[9];
  assign add_72139 = add_72126 + 32'h0000_0001;
  assign array_update_72140[0] = literal_72009 == 32'h0000_0000 ? array_update_72138 : array_update_72127[0];
  assign array_update_72140[1] = literal_72009 == 32'h0000_0001 ? array_update_72138 : array_update_72127[1];
  assign array_update_72140[2] = literal_72009 == 32'h0000_0002 ? array_update_72138 : array_update_72127[2];
  assign array_update_72140[3] = literal_72009 == 32'h0000_0003 ? array_update_72138 : array_update_72127[3];
  assign array_update_72140[4] = literal_72009 == 32'h0000_0004 ? array_update_72138 : array_update_72127[4];
  assign array_update_72140[5] = literal_72009 == 32'h0000_0005 ? array_update_72138 : array_update_72127[5];
  assign array_update_72140[6] = literal_72009 == 32'h0000_0006 ? array_update_72138 : array_update_72127[6];
  assign array_update_72140[7] = literal_72009 == 32'h0000_0007 ? array_update_72138 : array_update_72127[7];
  assign array_update_72140[8] = literal_72009 == 32'h0000_0008 ? array_update_72138 : array_update_72127[8];
  assign array_update_72140[9] = literal_72009 == 32'h0000_0009 ? array_update_72138 : array_update_72127[9];
  assign array_index_72142 = array_update_72021[add_72139 > 32'h0000_0009 ? 4'h9 : add_72139[3:0]];
  assign array_index_72143 = array_update_72140[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_72147 = smul32b_32b_x_32b(array_index_72024[add_72139 > 32'h0000_0009 ? 4'h9 : add_72139[3:0]], array_index_72142[literal_72016 > 32'h0000_0009 ? 4'h9 : literal_72016[3:0]]);
  assign add_72149 = array_index_72143[literal_72016 > 32'h0000_0009 ? 4'h9 : literal_72016[3:0]] + smul_72147;
  assign array_update_72150[0] = literal_72016 == 32'h0000_0000 ? add_72149 : array_index_72143[0];
  assign array_update_72150[1] = literal_72016 == 32'h0000_0001 ? add_72149 : array_index_72143[1];
  assign array_update_72150[2] = literal_72016 == 32'h0000_0002 ? add_72149 : array_index_72143[2];
  assign array_update_72150[3] = literal_72016 == 32'h0000_0003 ? add_72149 : array_index_72143[3];
  assign array_update_72150[4] = literal_72016 == 32'h0000_0004 ? add_72149 : array_index_72143[4];
  assign array_update_72150[5] = literal_72016 == 32'h0000_0005 ? add_72149 : array_index_72143[5];
  assign array_update_72150[6] = literal_72016 == 32'h0000_0006 ? add_72149 : array_index_72143[6];
  assign array_update_72150[7] = literal_72016 == 32'h0000_0007 ? add_72149 : array_index_72143[7];
  assign array_update_72150[8] = literal_72016 == 32'h0000_0008 ? add_72149 : array_index_72143[8];
  assign array_update_72150[9] = literal_72016 == 32'h0000_0009 ? add_72149 : array_index_72143[9];
  assign array_update_72151[0] = literal_72009 == 32'h0000_0000 ? array_update_72150 : array_update_72140[0];
  assign array_update_72151[1] = literal_72009 == 32'h0000_0001 ? array_update_72150 : array_update_72140[1];
  assign array_update_72151[2] = literal_72009 == 32'h0000_0002 ? array_update_72150 : array_update_72140[2];
  assign array_update_72151[3] = literal_72009 == 32'h0000_0003 ? array_update_72150 : array_update_72140[3];
  assign array_update_72151[4] = literal_72009 == 32'h0000_0004 ? array_update_72150 : array_update_72140[4];
  assign array_update_72151[5] = literal_72009 == 32'h0000_0005 ? array_update_72150 : array_update_72140[5];
  assign array_update_72151[6] = literal_72009 == 32'h0000_0006 ? array_update_72150 : array_update_72140[6];
  assign array_update_72151[7] = literal_72009 == 32'h0000_0007 ? array_update_72150 : array_update_72140[7];
  assign array_update_72151[8] = literal_72009 == 32'h0000_0008 ? array_update_72150 : array_update_72140[8];
  assign array_update_72151[9] = literal_72009 == 32'h0000_0009 ? array_update_72150 : array_update_72140[9];
  assign array_index_72153 = array_update_72151[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign add_72155 = literal_72016 + 32'h0000_0001;
  assign array_update_72156[0] = add_72155 == 32'h0000_0000 ? 32'h0000_0000 : array_index_72153[0];
  assign array_update_72156[1] = add_72155 == 32'h0000_0001 ? 32'h0000_0000 : array_index_72153[1];
  assign array_update_72156[2] = add_72155 == 32'h0000_0002 ? 32'h0000_0000 : array_index_72153[2];
  assign array_update_72156[3] = add_72155 == 32'h0000_0003 ? 32'h0000_0000 : array_index_72153[3];
  assign array_update_72156[4] = add_72155 == 32'h0000_0004 ? 32'h0000_0000 : array_index_72153[4];
  assign array_update_72156[5] = add_72155 == 32'h0000_0005 ? 32'h0000_0000 : array_index_72153[5];
  assign array_update_72156[6] = add_72155 == 32'h0000_0006 ? 32'h0000_0000 : array_index_72153[6];
  assign array_update_72156[7] = add_72155 == 32'h0000_0007 ? 32'h0000_0000 : array_index_72153[7];
  assign array_update_72156[8] = add_72155 == 32'h0000_0008 ? 32'h0000_0000 : array_index_72153[8];
  assign array_update_72156[9] = add_72155 == 32'h0000_0009 ? 32'h0000_0000 : array_index_72153[9];
  assign literal_72157 = 32'h0000_0000;
  assign array_update_72158[0] = literal_72009 == 32'h0000_0000 ? array_update_72156 : array_update_72151[0];
  assign array_update_72158[1] = literal_72009 == 32'h0000_0001 ? array_update_72156 : array_update_72151[1];
  assign array_update_72158[2] = literal_72009 == 32'h0000_0002 ? array_update_72156 : array_update_72151[2];
  assign array_update_72158[3] = literal_72009 == 32'h0000_0003 ? array_update_72156 : array_update_72151[3];
  assign array_update_72158[4] = literal_72009 == 32'h0000_0004 ? array_update_72156 : array_update_72151[4];
  assign array_update_72158[5] = literal_72009 == 32'h0000_0005 ? array_update_72156 : array_update_72151[5];
  assign array_update_72158[6] = literal_72009 == 32'h0000_0006 ? array_update_72156 : array_update_72151[6];
  assign array_update_72158[7] = literal_72009 == 32'h0000_0007 ? array_update_72156 : array_update_72151[7];
  assign array_update_72158[8] = literal_72009 == 32'h0000_0008 ? array_update_72156 : array_update_72151[8];
  assign array_update_72158[9] = literal_72009 == 32'h0000_0009 ? array_update_72156 : array_update_72151[9];
  assign array_index_72160 = array_update_72021[literal_72157 > 32'h0000_0009 ? 4'h9 : literal_72157[3:0]];
  assign array_index_72161 = array_update_72158[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_72165 = smul32b_32b_x_32b(array_index_72024[literal_72157 > 32'h0000_0009 ? 4'h9 : literal_72157[3:0]], array_index_72160[add_72155 > 32'h0000_0009 ? 4'h9 : add_72155[3:0]]);
  assign add_72167 = array_index_72161[add_72155 > 32'h0000_0009 ? 4'h9 : add_72155[3:0]] + smul_72165;
  assign array_update_72169[0] = add_72155 == 32'h0000_0000 ? add_72167 : array_index_72161[0];
  assign array_update_72169[1] = add_72155 == 32'h0000_0001 ? add_72167 : array_index_72161[1];
  assign array_update_72169[2] = add_72155 == 32'h0000_0002 ? add_72167 : array_index_72161[2];
  assign array_update_72169[3] = add_72155 == 32'h0000_0003 ? add_72167 : array_index_72161[3];
  assign array_update_72169[4] = add_72155 == 32'h0000_0004 ? add_72167 : array_index_72161[4];
  assign array_update_72169[5] = add_72155 == 32'h0000_0005 ? add_72167 : array_index_72161[5];
  assign array_update_72169[6] = add_72155 == 32'h0000_0006 ? add_72167 : array_index_72161[6];
  assign array_update_72169[7] = add_72155 == 32'h0000_0007 ? add_72167 : array_index_72161[7];
  assign array_update_72169[8] = add_72155 == 32'h0000_0008 ? add_72167 : array_index_72161[8];
  assign array_update_72169[9] = add_72155 == 32'h0000_0009 ? add_72167 : array_index_72161[9];
  assign add_72170 = literal_72157 + 32'h0000_0001;
  assign array_update_72171[0] = literal_72009 == 32'h0000_0000 ? array_update_72169 : array_update_72158[0];
  assign array_update_72171[1] = literal_72009 == 32'h0000_0001 ? array_update_72169 : array_update_72158[1];
  assign array_update_72171[2] = literal_72009 == 32'h0000_0002 ? array_update_72169 : array_update_72158[2];
  assign array_update_72171[3] = literal_72009 == 32'h0000_0003 ? array_update_72169 : array_update_72158[3];
  assign array_update_72171[4] = literal_72009 == 32'h0000_0004 ? array_update_72169 : array_update_72158[4];
  assign array_update_72171[5] = literal_72009 == 32'h0000_0005 ? array_update_72169 : array_update_72158[5];
  assign array_update_72171[6] = literal_72009 == 32'h0000_0006 ? array_update_72169 : array_update_72158[6];
  assign array_update_72171[7] = literal_72009 == 32'h0000_0007 ? array_update_72169 : array_update_72158[7];
  assign array_update_72171[8] = literal_72009 == 32'h0000_0008 ? array_update_72169 : array_update_72158[8];
  assign array_update_72171[9] = literal_72009 == 32'h0000_0009 ? array_update_72169 : array_update_72158[9];
  assign array_index_72173 = array_update_72021[add_72170 > 32'h0000_0009 ? 4'h9 : add_72170[3:0]];
  assign array_index_72174 = array_update_72171[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_72178 = smul32b_32b_x_32b(array_index_72024[add_72170 > 32'h0000_0009 ? 4'h9 : add_72170[3:0]], array_index_72173[add_72155 > 32'h0000_0009 ? 4'h9 : add_72155[3:0]]);
  assign add_72180 = array_index_72174[add_72155 > 32'h0000_0009 ? 4'h9 : add_72155[3:0]] + smul_72178;
  assign array_update_72182[0] = add_72155 == 32'h0000_0000 ? add_72180 : array_index_72174[0];
  assign array_update_72182[1] = add_72155 == 32'h0000_0001 ? add_72180 : array_index_72174[1];
  assign array_update_72182[2] = add_72155 == 32'h0000_0002 ? add_72180 : array_index_72174[2];
  assign array_update_72182[3] = add_72155 == 32'h0000_0003 ? add_72180 : array_index_72174[3];
  assign array_update_72182[4] = add_72155 == 32'h0000_0004 ? add_72180 : array_index_72174[4];
  assign array_update_72182[5] = add_72155 == 32'h0000_0005 ? add_72180 : array_index_72174[5];
  assign array_update_72182[6] = add_72155 == 32'h0000_0006 ? add_72180 : array_index_72174[6];
  assign array_update_72182[7] = add_72155 == 32'h0000_0007 ? add_72180 : array_index_72174[7];
  assign array_update_72182[8] = add_72155 == 32'h0000_0008 ? add_72180 : array_index_72174[8];
  assign array_update_72182[9] = add_72155 == 32'h0000_0009 ? add_72180 : array_index_72174[9];
  assign add_72183 = add_72170 + 32'h0000_0001;
  assign array_update_72184[0] = literal_72009 == 32'h0000_0000 ? array_update_72182 : array_update_72171[0];
  assign array_update_72184[1] = literal_72009 == 32'h0000_0001 ? array_update_72182 : array_update_72171[1];
  assign array_update_72184[2] = literal_72009 == 32'h0000_0002 ? array_update_72182 : array_update_72171[2];
  assign array_update_72184[3] = literal_72009 == 32'h0000_0003 ? array_update_72182 : array_update_72171[3];
  assign array_update_72184[4] = literal_72009 == 32'h0000_0004 ? array_update_72182 : array_update_72171[4];
  assign array_update_72184[5] = literal_72009 == 32'h0000_0005 ? array_update_72182 : array_update_72171[5];
  assign array_update_72184[6] = literal_72009 == 32'h0000_0006 ? array_update_72182 : array_update_72171[6];
  assign array_update_72184[7] = literal_72009 == 32'h0000_0007 ? array_update_72182 : array_update_72171[7];
  assign array_update_72184[8] = literal_72009 == 32'h0000_0008 ? array_update_72182 : array_update_72171[8];
  assign array_update_72184[9] = literal_72009 == 32'h0000_0009 ? array_update_72182 : array_update_72171[9];
  assign array_index_72186 = array_update_72021[add_72183 > 32'h0000_0009 ? 4'h9 : add_72183[3:0]];
  assign array_index_72187 = array_update_72184[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_72191 = smul32b_32b_x_32b(array_index_72024[add_72183 > 32'h0000_0009 ? 4'h9 : add_72183[3:0]], array_index_72186[add_72155 > 32'h0000_0009 ? 4'h9 : add_72155[3:0]]);
  assign add_72193 = array_index_72187[add_72155 > 32'h0000_0009 ? 4'h9 : add_72155[3:0]] + smul_72191;
  assign array_update_72195[0] = add_72155 == 32'h0000_0000 ? add_72193 : array_index_72187[0];
  assign array_update_72195[1] = add_72155 == 32'h0000_0001 ? add_72193 : array_index_72187[1];
  assign array_update_72195[2] = add_72155 == 32'h0000_0002 ? add_72193 : array_index_72187[2];
  assign array_update_72195[3] = add_72155 == 32'h0000_0003 ? add_72193 : array_index_72187[3];
  assign array_update_72195[4] = add_72155 == 32'h0000_0004 ? add_72193 : array_index_72187[4];
  assign array_update_72195[5] = add_72155 == 32'h0000_0005 ? add_72193 : array_index_72187[5];
  assign array_update_72195[6] = add_72155 == 32'h0000_0006 ? add_72193 : array_index_72187[6];
  assign array_update_72195[7] = add_72155 == 32'h0000_0007 ? add_72193 : array_index_72187[7];
  assign array_update_72195[8] = add_72155 == 32'h0000_0008 ? add_72193 : array_index_72187[8];
  assign array_update_72195[9] = add_72155 == 32'h0000_0009 ? add_72193 : array_index_72187[9];
  assign add_72196 = add_72183 + 32'h0000_0001;
  assign array_update_72197[0] = literal_72009 == 32'h0000_0000 ? array_update_72195 : array_update_72184[0];
  assign array_update_72197[1] = literal_72009 == 32'h0000_0001 ? array_update_72195 : array_update_72184[1];
  assign array_update_72197[2] = literal_72009 == 32'h0000_0002 ? array_update_72195 : array_update_72184[2];
  assign array_update_72197[3] = literal_72009 == 32'h0000_0003 ? array_update_72195 : array_update_72184[3];
  assign array_update_72197[4] = literal_72009 == 32'h0000_0004 ? array_update_72195 : array_update_72184[4];
  assign array_update_72197[5] = literal_72009 == 32'h0000_0005 ? array_update_72195 : array_update_72184[5];
  assign array_update_72197[6] = literal_72009 == 32'h0000_0006 ? array_update_72195 : array_update_72184[6];
  assign array_update_72197[7] = literal_72009 == 32'h0000_0007 ? array_update_72195 : array_update_72184[7];
  assign array_update_72197[8] = literal_72009 == 32'h0000_0008 ? array_update_72195 : array_update_72184[8];
  assign array_update_72197[9] = literal_72009 == 32'h0000_0009 ? array_update_72195 : array_update_72184[9];
  assign array_index_72199 = array_update_72021[add_72196 > 32'h0000_0009 ? 4'h9 : add_72196[3:0]];
  assign array_index_72200 = array_update_72197[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_72204 = smul32b_32b_x_32b(array_index_72024[add_72196 > 32'h0000_0009 ? 4'h9 : add_72196[3:0]], array_index_72199[add_72155 > 32'h0000_0009 ? 4'h9 : add_72155[3:0]]);
  assign add_72206 = array_index_72200[add_72155 > 32'h0000_0009 ? 4'h9 : add_72155[3:0]] + smul_72204;
  assign array_update_72208[0] = add_72155 == 32'h0000_0000 ? add_72206 : array_index_72200[0];
  assign array_update_72208[1] = add_72155 == 32'h0000_0001 ? add_72206 : array_index_72200[1];
  assign array_update_72208[2] = add_72155 == 32'h0000_0002 ? add_72206 : array_index_72200[2];
  assign array_update_72208[3] = add_72155 == 32'h0000_0003 ? add_72206 : array_index_72200[3];
  assign array_update_72208[4] = add_72155 == 32'h0000_0004 ? add_72206 : array_index_72200[4];
  assign array_update_72208[5] = add_72155 == 32'h0000_0005 ? add_72206 : array_index_72200[5];
  assign array_update_72208[6] = add_72155 == 32'h0000_0006 ? add_72206 : array_index_72200[6];
  assign array_update_72208[7] = add_72155 == 32'h0000_0007 ? add_72206 : array_index_72200[7];
  assign array_update_72208[8] = add_72155 == 32'h0000_0008 ? add_72206 : array_index_72200[8];
  assign array_update_72208[9] = add_72155 == 32'h0000_0009 ? add_72206 : array_index_72200[9];
  assign add_72209 = add_72196 + 32'h0000_0001;
  assign array_update_72210[0] = literal_72009 == 32'h0000_0000 ? array_update_72208 : array_update_72197[0];
  assign array_update_72210[1] = literal_72009 == 32'h0000_0001 ? array_update_72208 : array_update_72197[1];
  assign array_update_72210[2] = literal_72009 == 32'h0000_0002 ? array_update_72208 : array_update_72197[2];
  assign array_update_72210[3] = literal_72009 == 32'h0000_0003 ? array_update_72208 : array_update_72197[3];
  assign array_update_72210[4] = literal_72009 == 32'h0000_0004 ? array_update_72208 : array_update_72197[4];
  assign array_update_72210[5] = literal_72009 == 32'h0000_0005 ? array_update_72208 : array_update_72197[5];
  assign array_update_72210[6] = literal_72009 == 32'h0000_0006 ? array_update_72208 : array_update_72197[6];
  assign array_update_72210[7] = literal_72009 == 32'h0000_0007 ? array_update_72208 : array_update_72197[7];
  assign array_update_72210[8] = literal_72009 == 32'h0000_0008 ? array_update_72208 : array_update_72197[8];
  assign array_update_72210[9] = literal_72009 == 32'h0000_0009 ? array_update_72208 : array_update_72197[9];
  assign array_index_72212 = array_update_72021[add_72209 > 32'h0000_0009 ? 4'h9 : add_72209[3:0]];
  assign array_index_72213 = array_update_72210[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_72217 = smul32b_32b_x_32b(array_index_72024[add_72209 > 32'h0000_0009 ? 4'h9 : add_72209[3:0]], array_index_72212[add_72155 > 32'h0000_0009 ? 4'h9 : add_72155[3:0]]);
  assign add_72219 = array_index_72213[add_72155 > 32'h0000_0009 ? 4'h9 : add_72155[3:0]] + smul_72217;
  assign array_update_72221[0] = add_72155 == 32'h0000_0000 ? add_72219 : array_index_72213[0];
  assign array_update_72221[1] = add_72155 == 32'h0000_0001 ? add_72219 : array_index_72213[1];
  assign array_update_72221[2] = add_72155 == 32'h0000_0002 ? add_72219 : array_index_72213[2];
  assign array_update_72221[3] = add_72155 == 32'h0000_0003 ? add_72219 : array_index_72213[3];
  assign array_update_72221[4] = add_72155 == 32'h0000_0004 ? add_72219 : array_index_72213[4];
  assign array_update_72221[5] = add_72155 == 32'h0000_0005 ? add_72219 : array_index_72213[5];
  assign array_update_72221[6] = add_72155 == 32'h0000_0006 ? add_72219 : array_index_72213[6];
  assign array_update_72221[7] = add_72155 == 32'h0000_0007 ? add_72219 : array_index_72213[7];
  assign array_update_72221[8] = add_72155 == 32'h0000_0008 ? add_72219 : array_index_72213[8];
  assign array_update_72221[9] = add_72155 == 32'h0000_0009 ? add_72219 : array_index_72213[9];
  assign add_72222 = add_72209 + 32'h0000_0001;
  assign array_update_72223[0] = literal_72009 == 32'h0000_0000 ? array_update_72221 : array_update_72210[0];
  assign array_update_72223[1] = literal_72009 == 32'h0000_0001 ? array_update_72221 : array_update_72210[1];
  assign array_update_72223[2] = literal_72009 == 32'h0000_0002 ? array_update_72221 : array_update_72210[2];
  assign array_update_72223[3] = literal_72009 == 32'h0000_0003 ? array_update_72221 : array_update_72210[3];
  assign array_update_72223[4] = literal_72009 == 32'h0000_0004 ? array_update_72221 : array_update_72210[4];
  assign array_update_72223[5] = literal_72009 == 32'h0000_0005 ? array_update_72221 : array_update_72210[5];
  assign array_update_72223[6] = literal_72009 == 32'h0000_0006 ? array_update_72221 : array_update_72210[6];
  assign array_update_72223[7] = literal_72009 == 32'h0000_0007 ? array_update_72221 : array_update_72210[7];
  assign array_update_72223[8] = literal_72009 == 32'h0000_0008 ? array_update_72221 : array_update_72210[8];
  assign array_update_72223[9] = literal_72009 == 32'h0000_0009 ? array_update_72221 : array_update_72210[9];
  assign array_index_72225 = array_update_72021[add_72222 > 32'h0000_0009 ? 4'h9 : add_72222[3:0]];
  assign array_index_72226 = array_update_72223[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_72230 = smul32b_32b_x_32b(array_index_72024[add_72222 > 32'h0000_0009 ? 4'h9 : add_72222[3:0]], array_index_72225[add_72155 > 32'h0000_0009 ? 4'h9 : add_72155[3:0]]);
  assign add_72232 = array_index_72226[add_72155 > 32'h0000_0009 ? 4'h9 : add_72155[3:0]] + smul_72230;
  assign array_update_72234[0] = add_72155 == 32'h0000_0000 ? add_72232 : array_index_72226[0];
  assign array_update_72234[1] = add_72155 == 32'h0000_0001 ? add_72232 : array_index_72226[1];
  assign array_update_72234[2] = add_72155 == 32'h0000_0002 ? add_72232 : array_index_72226[2];
  assign array_update_72234[3] = add_72155 == 32'h0000_0003 ? add_72232 : array_index_72226[3];
  assign array_update_72234[4] = add_72155 == 32'h0000_0004 ? add_72232 : array_index_72226[4];
  assign array_update_72234[5] = add_72155 == 32'h0000_0005 ? add_72232 : array_index_72226[5];
  assign array_update_72234[6] = add_72155 == 32'h0000_0006 ? add_72232 : array_index_72226[6];
  assign array_update_72234[7] = add_72155 == 32'h0000_0007 ? add_72232 : array_index_72226[7];
  assign array_update_72234[8] = add_72155 == 32'h0000_0008 ? add_72232 : array_index_72226[8];
  assign array_update_72234[9] = add_72155 == 32'h0000_0009 ? add_72232 : array_index_72226[9];
  assign add_72235 = add_72222 + 32'h0000_0001;
  assign array_update_72236[0] = literal_72009 == 32'h0000_0000 ? array_update_72234 : array_update_72223[0];
  assign array_update_72236[1] = literal_72009 == 32'h0000_0001 ? array_update_72234 : array_update_72223[1];
  assign array_update_72236[2] = literal_72009 == 32'h0000_0002 ? array_update_72234 : array_update_72223[2];
  assign array_update_72236[3] = literal_72009 == 32'h0000_0003 ? array_update_72234 : array_update_72223[3];
  assign array_update_72236[4] = literal_72009 == 32'h0000_0004 ? array_update_72234 : array_update_72223[4];
  assign array_update_72236[5] = literal_72009 == 32'h0000_0005 ? array_update_72234 : array_update_72223[5];
  assign array_update_72236[6] = literal_72009 == 32'h0000_0006 ? array_update_72234 : array_update_72223[6];
  assign array_update_72236[7] = literal_72009 == 32'h0000_0007 ? array_update_72234 : array_update_72223[7];
  assign array_update_72236[8] = literal_72009 == 32'h0000_0008 ? array_update_72234 : array_update_72223[8];
  assign array_update_72236[9] = literal_72009 == 32'h0000_0009 ? array_update_72234 : array_update_72223[9];
  assign array_index_72238 = array_update_72021[add_72235 > 32'h0000_0009 ? 4'h9 : add_72235[3:0]];
  assign array_index_72239 = array_update_72236[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_72243 = smul32b_32b_x_32b(array_index_72024[add_72235 > 32'h0000_0009 ? 4'h9 : add_72235[3:0]], array_index_72238[add_72155 > 32'h0000_0009 ? 4'h9 : add_72155[3:0]]);
  assign add_72245 = array_index_72239[add_72155 > 32'h0000_0009 ? 4'h9 : add_72155[3:0]] + smul_72243;
  assign array_update_72247[0] = add_72155 == 32'h0000_0000 ? add_72245 : array_index_72239[0];
  assign array_update_72247[1] = add_72155 == 32'h0000_0001 ? add_72245 : array_index_72239[1];
  assign array_update_72247[2] = add_72155 == 32'h0000_0002 ? add_72245 : array_index_72239[2];
  assign array_update_72247[3] = add_72155 == 32'h0000_0003 ? add_72245 : array_index_72239[3];
  assign array_update_72247[4] = add_72155 == 32'h0000_0004 ? add_72245 : array_index_72239[4];
  assign array_update_72247[5] = add_72155 == 32'h0000_0005 ? add_72245 : array_index_72239[5];
  assign array_update_72247[6] = add_72155 == 32'h0000_0006 ? add_72245 : array_index_72239[6];
  assign array_update_72247[7] = add_72155 == 32'h0000_0007 ? add_72245 : array_index_72239[7];
  assign array_update_72247[8] = add_72155 == 32'h0000_0008 ? add_72245 : array_index_72239[8];
  assign array_update_72247[9] = add_72155 == 32'h0000_0009 ? add_72245 : array_index_72239[9];
  assign add_72248 = add_72235 + 32'h0000_0001;
  assign array_update_72249[0] = literal_72009 == 32'h0000_0000 ? array_update_72247 : array_update_72236[0];
  assign array_update_72249[1] = literal_72009 == 32'h0000_0001 ? array_update_72247 : array_update_72236[1];
  assign array_update_72249[2] = literal_72009 == 32'h0000_0002 ? array_update_72247 : array_update_72236[2];
  assign array_update_72249[3] = literal_72009 == 32'h0000_0003 ? array_update_72247 : array_update_72236[3];
  assign array_update_72249[4] = literal_72009 == 32'h0000_0004 ? array_update_72247 : array_update_72236[4];
  assign array_update_72249[5] = literal_72009 == 32'h0000_0005 ? array_update_72247 : array_update_72236[5];
  assign array_update_72249[6] = literal_72009 == 32'h0000_0006 ? array_update_72247 : array_update_72236[6];
  assign array_update_72249[7] = literal_72009 == 32'h0000_0007 ? array_update_72247 : array_update_72236[7];
  assign array_update_72249[8] = literal_72009 == 32'h0000_0008 ? array_update_72247 : array_update_72236[8];
  assign array_update_72249[9] = literal_72009 == 32'h0000_0009 ? array_update_72247 : array_update_72236[9];
  assign array_index_72251 = array_update_72021[add_72248 > 32'h0000_0009 ? 4'h9 : add_72248[3:0]];
  assign array_index_72252 = array_update_72249[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_72256 = smul32b_32b_x_32b(array_index_72024[add_72248 > 32'h0000_0009 ? 4'h9 : add_72248[3:0]], array_index_72251[add_72155 > 32'h0000_0009 ? 4'h9 : add_72155[3:0]]);
  assign add_72258 = array_index_72252[add_72155 > 32'h0000_0009 ? 4'h9 : add_72155[3:0]] + smul_72256;
  assign array_update_72260[0] = add_72155 == 32'h0000_0000 ? add_72258 : array_index_72252[0];
  assign array_update_72260[1] = add_72155 == 32'h0000_0001 ? add_72258 : array_index_72252[1];
  assign array_update_72260[2] = add_72155 == 32'h0000_0002 ? add_72258 : array_index_72252[2];
  assign array_update_72260[3] = add_72155 == 32'h0000_0003 ? add_72258 : array_index_72252[3];
  assign array_update_72260[4] = add_72155 == 32'h0000_0004 ? add_72258 : array_index_72252[4];
  assign array_update_72260[5] = add_72155 == 32'h0000_0005 ? add_72258 : array_index_72252[5];
  assign array_update_72260[6] = add_72155 == 32'h0000_0006 ? add_72258 : array_index_72252[6];
  assign array_update_72260[7] = add_72155 == 32'h0000_0007 ? add_72258 : array_index_72252[7];
  assign array_update_72260[8] = add_72155 == 32'h0000_0008 ? add_72258 : array_index_72252[8];
  assign array_update_72260[9] = add_72155 == 32'h0000_0009 ? add_72258 : array_index_72252[9];
  assign add_72261 = add_72248 + 32'h0000_0001;
  assign array_update_72262[0] = literal_72009 == 32'h0000_0000 ? array_update_72260 : array_update_72249[0];
  assign array_update_72262[1] = literal_72009 == 32'h0000_0001 ? array_update_72260 : array_update_72249[1];
  assign array_update_72262[2] = literal_72009 == 32'h0000_0002 ? array_update_72260 : array_update_72249[2];
  assign array_update_72262[3] = literal_72009 == 32'h0000_0003 ? array_update_72260 : array_update_72249[3];
  assign array_update_72262[4] = literal_72009 == 32'h0000_0004 ? array_update_72260 : array_update_72249[4];
  assign array_update_72262[5] = literal_72009 == 32'h0000_0005 ? array_update_72260 : array_update_72249[5];
  assign array_update_72262[6] = literal_72009 == 32'h0000_0006 ? array_update_72260 : array_update_72249[6];
  assign array_update_72262[7] = literal_72009 == 32'h0000_0007 ? array_update_72260 : array_update_72249[7];
  assign array_update_72262[8] = literal_72009 == 32'h0000_0008 ? array_update_72260 : array_update_72249[8];
  assign array_update_72262[9] = literal_72009 == 32'h0000_0009 ? array_update_72260 : array_update_72249[9];
  assign array_index_72264 = array_update_72021[add_72261 > 32'h0000_0009 ? 4'h9 : add_72261[3:0]];
  assign array_index_72265 = array_update_72262[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_72269 = smul32b_32b_x_32b(array_index_72024[add_72261 > 32'h0000_0009 ? 4'h9 : add_72261[3:0]], array_index_72264[add_72155 > 32'h0000_0009 ? 4'h9 : add_72155[3:0]]);
  assign add_72271 = array_index_72265[add_72155 > 32'h0000_0009 ? 4'h9 : add_72155[3:0]] + smul_72269;
  assign array_update_72273[0] = add_72155 == 32'h0000_0000 ? add_72271 : array_index_72265[0];
  assign array_update_72273[1] = add_72155 == 32'h0000_0001 ? add_72271 : array_index_72265[1];
  assign array_update_72273[2] = add_72155 == 32'h0000_0002 ? add_72271 : array_index_72265[2];
  assign array_update_72273[3] = add_72155 == 32'h0000_0003 ? add_72271 : array_index_72265[3];
  assign array_update_72273[4] = add_72155 == 32'h0000_0004 ? add_72271 : array_index_72265[4];
  assign array_update_72273[5] = add_72155 == 32'h0000_0005 ? add_72271 : array_index_72265[5];
  assign array_update_72273[6] = add_72155 == 32'h0000_0006 ? add_72271 : array_index_72265[6];
  assign array_update_72273[7] = add_72155 == 32'h0000_0007 ? add_72271 : array_index_72265[7];
  assign array_update_72273[8] = add_72155 == 32'h0000_0008 ? add_72271 : array_index_72265[8];
  assign array_update_72273[9] = add_72155 == 32'h0000_0009 ? add_72271 : array_index_72265[9];
  assign add_72274 = add_72261 + 32'h0000_0001;
  assign array_update_72275[0] = literal_72009 == 32'h0000_0000 ? array_update_72273 : array_update_72262[0];
  assign array_update_72275[1] = literal_72009 == 32'h0000_0001 ? array_update_72273 : array_update_72262[1];
  assign array_update_72275[2] = literal_72009 == 32'h0000_0002 ? array_update_72273 : array_update_72262[2];
  assign array_update_72275[3] = literal_72009 == 32'h0000_0003 ? array_update_72273 : array_update_72262[3];
  assign array_update_72275[4] = literal_72009 == 32'h0000_0004 ? array_update_72273 : array_update_72262[4];
  assign array_update_72275[5] = literal_72009 == 32'h0000_0005 ? array_update_72273 : array_update_72262[5];
  assign array_update_72275[6] = literal_72009 == 32'h0000_0006 ? array_update_72273 : array_update_72262[6];
  assign array_update_72275[7] = literal_72009 == 32'h0000_0007 ? array_update_72273 : array_update_72262[7];
  assign array_update_72275[8] = literal_72009 == 32'h0000_0008 ? array_update_72273 : array_update_72262[8];
  assign array_update_72275[9] = literal_72009 == 32'h0000_0009 ? array_update_72273 : array_update_72262[9];
  assign array_index_72277 = array_update_72021[add_72274 > 32'h0000_0009 ? 4'h9 : add_72274[3:0]];
  assign array_index_72278 = array_update_72275[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_72282 = smul32b_32b_x_32b(array_index_72024[add_72274 > 32'h0000_0009 ? 4'h9 : add_72274[3:0]], array_index_72277[add_72155 > 32'h0000_0009 ? 4'h9 : add_72155[3:0]]);
  assign add_72284 = array_index_72278[add_72155 > 32'h0000_0009 ? 4'h9 : add_72155[3:0]] + smul_72282;
  assign array_update_72285[0] = add_72155 == 32'h0000_0000 ? add_72284 : array_index_72278[0];
  assign array_update_72285[1] = add_72155 == 32'h0000_0001 ? add_72284 : array_index_72278[1];
  assign array_update_72285[2] = add_72155 == 32'h0000_0002 ? add_72284 : array_index_72278[2];
  assign array_update_72285[3] = add_72155 == 32'h0000_0003 ? add_72284 : array_index_72278[3];
  assign array_update_72285[4] = add_72155 == 32'h0000_0004 ? add_72284 : array_index_72278[4];
  assign array_update_72285[5] = add_72155 == 32'h0000_0005 ? add_72284 : array_index_72278[5];
  assign array_update_72285[6] = add_72155 == 32'h0000_0006 ? add_72284 : array_index_72278[6];
  assign array_update_72285[7] = add_72155 == 32'h0000_0007 ? add_72284 : array_index_72278[7];
  assign array_update_72285[8] = add_72155 == 32'h0000_0008 ? add_72284 : array_index_72278[8];
  assign array_update_72285[9] = add_72155 == 32'h0000_0009 ? add_72284 : array_index_72278[9];
  assign array_update_72286[0] = literal_72009 == 32'h0000_0000 ? array_update_72285 : array_update_72275[0];
  assign array_update_72286[1] = literal_72009 == 32'h0000_0001 ? array_update_72285 : array_update_72275[1];
  assign array_update_72286[2] = literal_72009 == 32'h0000_0002 ? array_update_72285 : array_update_72275[2];
  assign array_update_72286[3] = literal_72009 == 32'h0000_0003 ? array_update_72285 : array_update_72275[3];
  assign array_update_72286[4] = literal_72009 == 32'h0000_0004 ? array_update_72285 : array_update_72275[4];
  assign array_update_72286[5] = literal_72009 == 32'h0000_0005 ? array_update_72285 : array_update_72275[5];
  assign array_update_72286[6] = literal_72009 == 32'h0000_0006 ? array_update_72285 : array_update_72275[6];
  assign array_update_72286[7] = literal_72009 == 32'h0000_0007 ? array_update_72285 : array_update_72275[7];
  assign array_update_72286[8] = literal_72009 == 32'h0000_0008 ? array_update_72285 : array_update_72275[8];
  assign array_update_72286[9] = literal_72009 == 32'h0000_0009 ? array_update_72285 : array_update_72275[9];
  assign array_index_72288 = array_update_72286[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign add_72290 = add_72155 + 32'h0000_0001;
  assign array_update_72291[0] = add_72290 == 32'h0000_0000 ? 32'h0000_0000 : array_index_72288[0];
  assign array_update_72291[1] = add_72290 == 32'h0000_0001 ? 32'h0000_0000 : array_index_72288[1];
  assign array_update_72291[2] = add_72290 == 32'h0000_0002 ? 32'h0000_0000 : array_index_72288[2];
  assign array_update_72291[3] = add_72290 == 32'h0000_0003 ? 32'h0000_0000 : array_index_72288[3];
  assign array_update_72291[4] = add_72290 == 32'h0000_0004 ? 32'h0000_0000 : array_index_72288[4];
  assign array_update_72291[5] = add_72290 == 32'h0000_0005 ? 32'h0000_0000 : array_index_72288[5];
  assign array_update_72291[6] = add_72290 == 32'h0000_0006 ? 32'h0000_0000 : array_index_72288[6];
  assign array_update_72291[7] = add_72290 == 32'h0000_0007 ? 32'h0000_0000 : array_index_72288[7];
  assign array_update_72291[8] = add_72290 == 32'h0000_0008 ? 32'h0000_0000 : array_index_72288[8];
  assign array_update_72291[9] = add_72290 == 32'h0000_0009 ? 32'h0000_0000 : array_index_72288[9];
  assign literal_72292 = 32'h0000_0000;
  assign array_update_72293[0] = literal_72009 == 32'h0000_0000 ? array_update_72291 : array_update_72286[0];
  assign array_update_72293[1] = literal_72009 == 32'h0000_0001 ? array_update_72291 : array_update_72286[1];
  assign array_update_72293[2] = literal_72009 == 32'h0000_0002 ? array_update_72291 : array_update_72286[2];
  assign array_update_72293[3] = literal_72009 == 32'h0000_0003 ? array_update_72291 : array_update_72286[3];
  assign array_update_72293[4] = literal_72009 == 32'h0000_0004 ? array_update_72291 : array_update_72286[4];
  assign array_update_72293[5] = literal_72009 == 32'h0000_0005 ? array_update_72291 : array_update_72286[5];
  assign array_update_72293[6] = literal_72009 == 32'h0000_0006 ? array_update_72291 : array_update_72286[6];
  assign array_update_72293[7] = literal_72009 == 32'h0000_0007 ? array_update_72291 : array_update_72286[7];
  assign array_update_72293[8] = literal_72009 == 32'h0000_0008 ? array_update_72291 : array_update_72286[8];
  assign array_update_72293[9] = literal_72009 == 32'h0000_0009 ? array_update_72291 : array_update_72286[9];
  assign array_index_72295 = array_update_72021[literal_72292 > 32'h0000_0009 ? 4'h9 : literal_72292[3:0]];
  assign array_index_72296 = array_update_72293[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_72300 = smul32b_32b_x_32b(array_index_72024[literal_72292 > 32'h0000_0009 ? 4'h9 : literal_72292[3:0]], array_index_72295[add_72290 > 32'h0000_0009 ? 4'h9 : add_72290[3:0]]);
  assign add_72302 = array_index_72296[add_72290 > 32'h0000_0009 ? 4'h9 : add_72290[3:0]] + smul_72300;
  assign array_update_72304[0] = add_72290 == 32'h0000_0000 ? add_72302 : array_index_72296[0];
  assign array_update_72304[1] = add_72290 == 32'h0000_0001 ? add_72302 : array_index_72296[1];
  assign array_update_72304[2] = add_72290 == 32'h0000_0002 ? add_72302 : array_index_72296[2];
  assign array_update_72304[3] = add_72290 == 32'h0000_0003 ? add_72302 : array_index_72296[3];
  assign array_update_72304[4] = add_72290 == 32'h0000_0004 ? add_72302 : array_index_72296[4];
  assign array_update_72304[5] = add_72290 == 32'h0000_0005 ? add_72302 : array_index_72296[5];
  assign array_update_72304[6] = add_72290 == 32'h0000_0006 ? add_72302 : array_index_72296[6];
  assign array_update_72304[7] = add_72290 == 32'h0000_0007 ? add_72302 : array_index_72296[7];
  assign array_update_72304[8] = add_72290 == 32'h0000_0008 ? add_72302 : array_index_72296[8];
  assign array_update_72304[9] = add_72290 == 32'h0000_0009 ? add_72302 : array_index_72296[9];
  assign add_72305 = literal_72292 + 32'h0000_0001;
  assign array_update_72306[0] = literal_72009 == 32'h0000_0000 ? array_update_72304 : array_update_72293[0];
  assign array_update_72306[1] = literal_72009 == 32'h0000_0001 ? array_update_72304 : array_update_72293[1];
  assign array_update_72306[2] = literal_72009 == 32'h0000_0002 ? array_update_72304 : array_update_72293[2];
  assign array_update_72306[3] = literal_72009 == 32'h0000_0003 ? array_update_72304 : array_update_72293[3];
  assign array_update_72306[4] = literal_72009 == 32'h0000_0004 ? array_update_72304 : array_update_72293[4];
  assign array_update_72306[5] = literal_72009 == 32'h0000_0005 ? array_update_72304 : array_update_72293[5];
  assign array_update_72306[6] = literal_72009 == 32'h0000_0006 ? array_update_72304 : array_update_72293[6];
  assign array_update_72306[7] = literal_72009 == 32'h0000_0007 ? array_update_72304 : array_update_72293[7];
  assign array_update_72306[8] = literal_72009 == 32'h0000_0008 ? array_update_72304 : array_update_72293[8];
  assign array_update_72306[9] = literal_72009 == 32'h0000_0009 ? array_update_72304 : array_update_72293[9];
  assign array_index_72308 = array_update_72021[add_72305 > 32'h0000_0009 ? 4'h9 : add_72305[3:0]];
  assign array_index_72309 = array_update_72306[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_72313 = smul32b_32b_x_32b(array_index_72024[add_72305 > 32'h0000_0009 ? 4'h9 : add_72305[3:0]], array_index_72308[add_72290 > 32'h0000_0009 ? 4'h9 : add_72290[3:0]]);
  assign add_72315 = array_index_72309[add_72290 > 32'h0000_0009 ? 4'h9 : add_72290[3:0]] + smul_72313;
  assign array_update_72317[0] = add_72290 == 32'h0000_0000 ? add_72315 : array_index_72309[0];
  assign array_update_72317[1] = add_72290 == 32'h0000_0001 ? add_72315 : array_index_72309[1];
  assign array_update_72317[2] = add_72290 == 32'h0000_0002 ? add_72315 : array_index_72309[2];
  assign array_update_72317[3] = add_72290 == 32'h0000_0003 ? add_72315 : array_index_72309[3];
  assign array_update_72317[4] = add_72290 == 32'h0000_0004 ? add_72315 : array_index_72309[4];
  assign array_update_72317[5] = add_72290 == 32'h0000_0005 ? add_72315 : array_index_72309[5];
  assign array_update_72317[6] = add_72290 == 32'h0000_0006 ? add_72315 : array_index_72309[6];
  assign array_update_72317[7] = add_72290 == 32'h0000_0007 ? add_72315 : array_index_72309[7];
  assign array_update_72317[8] = add_72290 == 32'h0000_0008 ? add_72315 : array_index_72309[8];
  assign array_update_72317[9] = add_72290 == 32'h0000_0009 ? add_72315 : array_index_72309[9];
  assign add_72318 = add_72305 + 32'h0000_0001;
  assign array_update_72319[0] = literal_72009 == 32'h0000_0000 ? array_update_72317 : array_update_72306[0];
  assign array_update_72319[1] = literal_72009 == 32'h0000_0001 ? array_update_72317 : array_update_72306[1];
  assign array_update_72319[2] = literal_72009 == 32'h0000_0002 ? array_update_72317 : array_update_72306[2];
  assign array_update_72319[3] = literal_72009 == 32'h0000_0003 ? array_update_72317 : array_update_72306[3];
  assign array_update_72319[4] = literal_72009 == 32'h0000_0004 ? array_update_72317 : array_update_72306[4];
  assign array_update_72319[5] = literal_72009 == 32'h0000_0005 ? array_update_72317 : array_update_72306[5];
  assign array_update_72319[6] = literal_72009 == 32'h0000_0006 ? array_update_72317 : array_update_72306[6];
  assign array_update_72319[7] = literal_72009 == 32'h0000_0007 ? array_update_72317 : array_update_72306[7];
  assign array_update_72319[8] = literal_72009 == 32'h0000_0008 ? array_update_72317 : array_update_72306[8];
  assign array_update_72319[9] = literal_72009 == 32'h0000_0009 ? array_update_72317 : array_update_72306[9];
  assign array_index_72321 = array_update_72021[add_72318 > 32'h0000_0009 ? 4'h9 : add_72318[3:0]];
  assign array_index_72322 = array_update_72319[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_72326 = smul32b_32b_x_32b(array_index_72024[add_72318 > 32'h0000_0009 ? 4'h9 : add_72318[3:0]], array_index_72321[add_72290 > 32'h0000_0009 ? 4'h9 : add_72290[3:0]]);
  assign add_72328 = array_index_72322[add_72290 > 32'h0000_0009 ? 4'h9 : add_72290[3:0]] + smul_72326;
  assign array_update_72330[0] = add_72290 == 32'h0000_0000 ? add_72328 : array_index_72322[0];
  assign array_update_72330[1] = add_72290 == 32'h0000_0001 ? add_72328 : array_index_72322[1];
  assign array_update_72330[2] = add_72290 == 32'h0000_0002 ? add_72328 : array_index_72322[2];
  assign array_update_72330[3] = add_72290 == 32'h0000_0003 ? add_72328 : array_index_72322[3];
  assign array_update_72330[4] = add_72290 == 32'h0000_0004 ? add_72328 : array_index_72322[4];
  assign array_update_72330[5] = add_72290 == 32'h0000_0005 ? add_72328 : array_index_72322[5];
  assign array_update_72330[6] = add_72290 == 32'h0000_0006 ? add_72328 : array_index_72322[6];
  assign array_update_72330[7] = add_72290 == 32'h0000_0007 ? add_72328 : array_index_72322[7];
  assign array_update_72330[8] = add_72290 == 32'h0000_0008 ? add_72328 : array_index_72322[8];
  assign array_update_72330[9] = add_72290 == 32'h0000_0009 ? add_72328 : array_index_72322[9];
  assign add_72331 = add_72318 + 32'h0000_0001;
  assign array_update_72332[0] = literal_72009 == 32'h0000_0000 ? array_update_72330 : array_update_72319[0];
  assign array_update_72332[1] = literal_72009 == 32'h0000_0001 ? array_update_72330 : array_update_72319[1];
  assign array_update_72332[2] = literal_72009 == 32'h0000_0002 ? array_update_72330 : array_update_72319[2];
  assign array_update_72332[3] = literal_72009 == 32'h0000_0003 ? array_update_72330 : array_update_72319[3];
  assign array_update_72332[4] = literal_72009 == 32'h0000_0004 ? array_update_72330 : array_update_72319[4];
  assign array_update_72332[5] = literal_72009 == 32'h0000_0005 ? array_update_72330 : array_update_72319[5];
  assign array_update_72332[6] = literal_72009 == 32'h0000_0006 ? array_update_72330 : array_update_72319[6];
  assign array_update_72332[7] = literal_72009 == 32'h0000_0007 ? array_update_72330 : array_update_72319[7];
  assign array_update_72332[8] = literal_72009 == 32'h0000_0008 ? array_update_72330 : array_update_72319[8];
  assign array_update_72332[9] = literal_72009 == 32'h0000_0009 ? array_update_72330 : array_update_72319[9];
  assign array_index_72334 = array_update_72021[add_72331 > 32'h0000_0009 ? 4'h9 : add_72331[3:0]];
  assign array_index_72335 = array_update_72332[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_72339 = smul32b_32b_x_32b(array_index_72024[add_72331 > 32'h0000_0009 ? 4'h9 : add_72331[3:0]], array_index_72334[add_72290 > 32'h0000_0009 ? 4'h9 : add_72290[3:0]]);
  assign add_72341 = array_index_72335[add_72290 > 32'h0000_0009 ? 4'h9 : add_72290[3:0]] + smul_72339;
  assign array_update_72343[0] = add_72290 == 32'h0000_0000 ? add_72341 : array_index_72335[0];
  assign array_update_72343[1] = add_72290 == 32'h0000_0001 ? add_72341 : array_index_72335[1];
  assign array_update_72343[2] = add_72290 == 32'h0000_0002 ? add_72341 : array_index_72335[2];
  assign array_update_72343[3] = add_72290 == 32'h0000_0003 ? add_72341 : array_index_72335[3];
  assign array_update_72343[4] = add_72290 == 32'h0000_0004 ? add_72341 : array_index_72335[4];
  assign array_update_72343[5] = add_72290 == 32'h0000_0005 ? add_72341 : array_index_72335[5];
  assign array_update_72343[6] = add_72290 == 32'h0000_0006 ? add_72341 : array_index_72335[6];
  assign array_update_72343[7] = add_72290 == 32'h0000_0007 ? add_72341 : array_index_72335[7];
  assign array_update_72343[8] = add_72290 == 32'h0000_0008 ? add_72341 : array_index_72335[8];
  assign array_update_72343[9] = add_72290 == 32'h0000_0009 ? add_72341 : array_index_72335[9];
  assign add_72344 = add_72331 + 32'h0000_0001;
  assign array_update_72345[0] = literal_72009 == 32'h0000_0000 ? array_update_72343 : array_update_72332[0];
  assign array_update_72345[1] = literal_72009 == 32'h0000_0001 ? array_update_72343 : array_update_72332[1];
  assign array_update_72345[2] = literal_72009 == 32'h0000_0002 ? array_update_72343 : array_update_72332[2];
  assign array_update_72345[3] = literal_72009 == 32'h0000_0003 ? array_update_72343 : array_update_72332[3];
  assign array_update_72345[4] = literal_72009 == 32'h0000_0004 ? array_update_72343 : array_update_72332[4];
  assign array_update_72345[5] = literal_72009 == 32'h0000_0005 ? array_update_72343 : array_update_72332[5];
  assign array_update_72345[6] = literal_72009 == 32'h0000_0006 ? array_update_72343 : array_update_72332[6];
  assign array_update_72345[7] = literal_72009 == 32'h0000_0007 ? array_update_72343 : array_update_72332[7];
  assign array_update_72345[8] = literal_72009 == 32'h0000_0008 ? array_update_72343 : array_update_72332[8];
  assign array_update_72345[9] = literal_72009 == 32'h0000_0009 ? array_update_72343 : array_update_72332[9];
  assign array_index_72347 = array_update_72021[add_72344 > 32'h0000_0009 ? 4'h9 : add_72344[3:0]];
  assign array_index_72348 = array_update_72345[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_72352 = smul32b_32b_x_32b(array_index_72024[add_72344 > 32'h0000_0009 ? 4'h9 : add_72344[3:0]], array_index_72347[add_72290 > 32'h0000_0009 ? 4'h9 : add_72290[3:0]]);
  assign add_72354 = array_index_72348[add_72290 > 32'h0000_0009 ? 4'h9 : add_72290[3:0]] + smul_72352;
  assign array_update_72356[0] = add_72290 == 32'h0000_0000 ? add_72354 : array_index_72348[0];
  assign array_update_72356[1] = add_72290 == 32'h0000_0001 ? add_72354 : array_index_72348[1];
  assign array_update_72356[2] = add_72290 == 32'h0000_0002 ? add_72354 : array_index_72348[2];
  assign array_update_72356[3] = add_72290 == 32'h0000_0003 ? add_72354 : array_index_72348[3];
  assign array_update_72356[4] = add_72290 == 32'h0000_0004 ? add_72354 : array_index_72348[4];
  assign array_update_72356[5] = add_72290 == 32'h0000_0005 ? add_72354 : array_index_72348[5];
  assign array_update_72356[6] = add_72290 == 32'h0000_0006 ? add_72354 : array_index_72348[6];
  assign array_update_72356[7] = add_72290 == 32'h0000_0007 ? add_72354 : array_index_72348[7];
  assign array_update_72356[8] = add_72290 == 32'h0000_0008 ? add_72354 : array_index_72348[8];
  assign array_update_72356[9] = add_72290 == 32'h0000_0009 ? add_72354 : array_index_72348[9];
  assign add_72357 = add_72344 + 32'h0000_0001;
  assign array_update_72358[0] = literal_72009 == 32'h0000_0000 ? array_update_72356 : array_update_72345[0];
  assign array_update_72358[1] = literal_72009 == 32'h0000_0001 ? array_update_72356 : array_update_72345[1];
  assign array_update_72358[2] = literal_72009 == 32'h0000_0002 ? array_update_72356 : array_update_72345[2];
  assign array_update_72358[3] = literal_72009 == 32'h0000_0003 ? array_update_72356 : array_update_72345[3];
  assign array_update_72358[4] = literal_72009 == 32'h0000_0004 ? array_update_72356 : array_update_72345[4];
  assign array_update_72358[5] = literal_72009 == 32'h0000_0005 ? array_update_72356 : array_update_72345[5];
  assign array_update_72358[6] = literal_72009 == 32'h0000_0006 ? array_update_72356 : array_update_72345[6];
  assign array_update_72358[7] = literal_72009 == 32'h0000_0007 ? array_update_72356 : array_update_72345[7];
  assign array_update_72358[8] = literal_72009 == 32'h0000_0008 ? array_update_72356 : array_update_72345[8];
  assign array_update_72358[9] = literal_72009 == 32'h0000_0009 ? array_update_72356 : array_update_72345[9];
  assign array_index_72360 = array_update_72021[add_72357 > 32'h0000_0009 ? 4'h9 : add_72357[3:0]];
  assign array_index_72361 = array_update_72358[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_72365 = smul32b_32b_x_32b(array_index_72024[add_72357 > 32'h0000_0009 ? 4'h9 : add_72357[3:0]], array_index_72360[add_72290 > 32'h0000_0009 ? 4'h9 : add_72290[3:0]]);
  assign add_72367 = array_index_72361[add_72290 > 32'h0000_0009 ? 4'h9 : add_72290[3:0]] + smul_72365;
  assign array_update_72369[0] = add_72290 == 32'h0000_0000 ? add_72367 : array_index_72361[0];
  assign array_update_72369[1] = add_72290 == 32'h0000_0001 ? add_72367 : array_index_72361[1];
  assign array_update_72369[2] = add_72290 == 32'h0000_0002 ? add_72367 : array_index_72361[2];
  assign array_update_72369[3] = add_72290 == 32'h0000_0003 ? add_72367 : array_index_72361[3];
  assign array_update_72369[4] = add_72290 == 32'h0000_0004 ? add_72367 : array_index_72361[4];
  assign array_update_72369[5] = add_72290 == 32'h0000_0005 ? add_72367 : array_index_72361[5];
  assign array_update_72369[6] = add_72290 == 32'h0000_0006 ? add_72367 : array_index_72361[6];
  assign array_update_72369[7] = add_72290 == 32'h0000_0007 ? add_72367 : array_index_72361[7];
  assign array_update_72369[8] = add_72290 == 32'h0000_0008 ? add_72367 : array_index_72361[8];
  assign array_update_72369[9] = add_72290 == 32'h0000_0009 ? add_72367 : array_index_72361[9];
  assign add_72370 = add_72357 + 32'h0000_0001;
  assign array_update_72371[0] = literal_72009 == 32'h0000_0000 ? array_update_72369 : array_update_72358[0];
  assign array_update_72371[1] = literal_72009 == 32'h0000_0001 ? array_update_72369 : array_update_72358[1];
  assign array_update_72371[2] = literal_72009 == 32'h0000_0002 ? array_update_72369 : array_update_72358[2];
  assign array_update_72371[3] = literal_72009 == 32'h0000_0003 ? array_update_72369 : array_update_72358[3];
  assign array_update_72371[4] = literal_72009 == 32'h0000_0004 ? array_update_72369 : array_update_72358[4];
  assign array_update_72371[5] = literal_72009 == 32'h0000_0005 ? array_update_72369 : array_update_72358[5];
  assign array_update_72371[6] = literal_72009 == 32'h0000_0006 ? array_update_72369 : array_update_72358[6];
  assign array_update_72371[7] = literal_72009 == 32'h0000_0007 ? array_update_72369 : array_update_72358[7];
  assign array_update_72371[8] = literal_72009 == 32'h0000_0008 ? array_update_72369 : array_update_72358[8];
  assign array_update_72371[9] = literal_72009 == 32'h0000_0009 ? array_update_72369 : array_update_72358[9];
  assign array_index_72373 = array_update_72021[add_72370 > 32'h0000_0009 ? 4'h9 : add_72370[3:0]];
  assign array_index_72374 = array_update_72371[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_72378 = smul32b_32b_x_32b(array_index_72024[add_72370 > 32'h0000_0009 ? 4'h9 : add_72370[3:0]], array_index_72373[add_72290 > 32'h0000_0009 ? 4'h9 : add_72290[3:0]]);
  assign add_72380 = array_index_72374[add_72290 > 32'h0000_0009 ? 4'h9 : add_72290[3:0]] + smul_72378;
  assign array_update_72382[0] = add_72290 == 32'h0000_0000 ? add_72380 : array_index_72374[0];
  assign array_update_72382[1] = add_72290 == 32'h0000_0001 ? add_72380 : array_index_72374[1];
  assign array_update_72382[2] = add_72290 == 32'h0000_0002 ? add_72380 : array_index_72374[2];
  assign array_update_72382[3] = add_72290 == 32'h0000_0003 ? add_72380 : array_index_72374[3];
  assign array_update_72382[4] = add_72290 == 32'h0000_0004 ? add_72380 : array_index_72374[4];
  assign array_update_72382[5] = add_72290 == 32'h0000_0005 ? add_72380 : array_index_72374[5];
  assign array_update_72382[6] = add_72290 == 32'h0000_0006 ? add_72380 : array_index_72374[6];
  assign array_update_72382[7] = add_72290 == 32'h0000_0007 ? add_72380 : array_index_72374[7];
  assign array_update_72382[8] = add_72290 == 32'h0000_0008 ? add_72380 : array_index_72374[8];
  assign array_update_72382[9] = add_72290 == 32'h0000_0009 ? add_72380 : array_index_72374[9];
  assign add_72383 = add_72370 + 32'h0000_0001;
  assign array_update_72384[0] = literal_72009 == 32'h0000_0000 ? array_update_72382 : array_update_72371[0];
  assign array_update_72384[1] = literal_72009 == 32'h0000_0001 ? array_update_72382 : array_update_72371[1];
  assign array_update_72384[2] = literal_72009 == 32'h0000_0002 ? array_update_72382 : array_update_72371[2];
  assign array_update_72384[3] = literal_72009 == 32'h0000_0003 ? array_update_72382 : array_update_72371[3];
  assign array_update_72384[4] = literal_72009 == 32'h0000_0004 ? array_update_72382 : array_update_72371[4];
  assign array_update_72384[5] = literal_72009 == 32'h0000_0005 ? array_update_72382 : array_update_72371[5];
  assign array_update_72384[6] = literal_72009 == 32'h0000_0006 ? array_update_72382 : array_update_72371[6];
  assign array_update_72384[7] = literal_72009 == 32'h0000_0007 ? array_update_72382 : array_update_72371[7];
  assign array_update_72384[8] = literal_72009 == 32'h0000_0008 ? array_update_72382 : array_update_72371[8];
  assign array_update_72384[9] = literal_72009 == 32'h0000_0009 ? array_update_72382 : array_update_72371[9];
  assign array_index_72386 = array_update_72021[add_72383 > 32'h0000_0009 ? 4'h9 : add_72383[3:0]];
  assign array_index_72387 = array_update_72384[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_72391 = smul32b_32b_x_32b(array_index_72024[add_72383 > 32'h0000_0009 ? 4'h9 : add_72383[3:0]], array_index_72386[add_72290 > 32'h0000_0009 ? 4'h9 : add_72290[3:0]]);
  assign add_72393 = array_index_72387[add_72290 > 32'h0000_0009 ? 4'h9 : add_72290[3:0]] + smul_72391;
  assign array_update_72395[0] = add_72290 == 32'h0000_0000 ? add_72393 : array_index_72387[0];
  assign array_update_72395[1] = add_72290 == 32'h0000_0001 ? add_72393 : array_index_72387[1];
  assign array_update_72395[2] = add_72290 == 32'h0000_0002 ? add_72393 : array_index_72387[2];
  assign array_update_72395[3] = add_72290 == 32'h0000_0003 ? add_72393 : array_index_72387[3];
  assign array_update_72395[4] = add_72290 == 32'h0000_0004 ? add_72393 : array_index_72387[4];
  assign array_update_72395[5] = add_72290 == 32'h0000_0005 ? add_72393 : array_index_72387[5];
  assign array_update_72395[6] = add_72290 == 32'h0000_0006 ? add_72393 : array_index_72387[6];
  assign array_update_72395[7] = add_72290 == 32'h0000_0007 ? add_72393 : array_index_72387[7];
  assign array_update_72395[8] = add_72290 == 32'h0000_0008 ? add_72393 : array_index_72387[8];
  assign array_update_72395[9] = add_72290 == 32'h0000_0009 ? add_72393 : array_index_72387[9];
  assign add_72396 = add_72383 + 32'h0000_0001;
  assign array_update_72397[0] = literal_72009 == 32'h0000_0000 ? array_update_72395 : array_update_72384[0];
  assign array_update_72397[1] = literal_72009 == 32'h0000_0001 ? array_update_72395 : array_update_72384[1];
  assign array_update_72397[2] = literal_72009 == 32'h0000_0002 ? array_update_72395 : array_update_72384[2];
  assign array_update_72397[3] = literal_72009 == 32'h0000_0003 ? array_update_72395 : array_update_72384[3];
  assign array_update_72397[4] = literal_72009 == 32'h0000_0004 ? array_update_72395 : array_update_72384[4];
  assign array_update_72397[5] = literal_72009 == 32'h0000_0005 ? array_update_72395 : array_update_72384[5];
  assign array_update_72397[6] = literal_72009 == 32'h0000_0006 ? array_update_72395 : array_update_72384[6];
  assign array_update_72397[7] = literal_72009 == 32'h0000_0007 ? array_update_72395 : array_update_72384[7];
  assign array_update_72397[8] = literal_72009 == 32'h0000_0008 ? array_update_72395 : array_update_72384[8];
  assign array_update_72397[9] = literal_72009 == 32'h0000_0009 ? array_update_72395 : array_update_72384[9];
  assign array_index_72399 = array_update_72021[add_72396 > 32'h0000_0009 ? 4'h9 : add_72396[3:0]];
  assign array_index_72400 = array_update_72397[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_72404 = smul32b_32b_x_32b(array_index_72024[add_72396 > 32'h0000_0009 ? 4'h9 : add_72396[3:0]], array_index_72399[add_72290 > 32'h0000_0009 ? 4'h9 : add_72290[3:0]]);
  assign add_72406 = array_index_72400[add_72290 > 32'h0000_0009 ? 4'h9 : add_72290[3:0]] + smul_72404;
  assign array_update_72408[0] = add_72290 == 32'h0000_0000 ? add_72406 : array_index_72400[0];
  assign array_update_72408[1] = add_72290 == 32'h0000_0001 ? add_72406 : array_index_72400[1];
  assign array_update_72408[2] = add_72290 == 32'h0000_0002 ? add_72406 : array_index_72400[2];
  assign array_update_72408[3] = add_72290 == 32'h0000_0003 ? add_72406 : array_index_72400[3];
  assign array_update_72408[4] = add_72290 == 32'h0000_0004 ? add_72406 : array_index_72400[4];
  assign array_update_72408[5] = add_72290 == 32'h0000_0005 ? add_72406 : array_index_72400[5];
  assign array_update_72408[6] = add_72290 == 32'h0000_0006 ? add_72406 : array_index_72400[6];
  assign array_update_72408[7] = add_72290 == 32'h0000_0007 ? add_72406 : array_index_72400[7];
  assign array_update_72408[8] = add_72290 == 32'h0000_0008 ? add_72406 : array_index_72400[8];
  assign array_update_72408[9] = add_72290 == 32'h0000_0009 ? add_72406 : array_index_72400[9];
  assign add_72409 = add_72396 + 32'h0000_0001;
  assign array_update_72410[0] = literal_72009 == 32'h0000_0000 ? array_update_72408 : array_update_72397[0];
  assign array_update_72410[1] = literal_72009 == 32'h0000_0001 ? array_update_72408 : array_update_72397[1];
  assign array_update_72410[2] = literal_72009 == 32'h0000_0002 ? array_update_72408 : array_update_72397[2];
  assign array_update_72410[3] = literal_72009 == 32'h0000_0003 ? array_update_72408 : array_update_72397[3];
  assign array_update_72410[4] = literal_72009 == 32'h0000_0004 ? array_update_72408 : array_update_72397[4];
  assign array_update_72410[5] = literal_72009 == 32'h0000_0005 ? array_update_72408 : array_update_72397[5];
  assign array_update_72410[6] = literal_72009 == 32'h0000_0006 ? array_update_72408 : array_update_72397[6];
  assign array_update_72410[7] = literal_72009 == 32'h0000_0007 ? array_update_72408 : array_update_72397[7];
  assign array_update_72410[8] = literal_72009 == 32'h0000_0008 ? array_update_72408 : array_update_72397[8];
  assign array_update_72410[9] = literal_72009 == 32'h0000_0009 ? array_update_72408 : array_update_72397[9];
  assign array_index_72412 = array_update_72021[add_72409 > 32'h0000_0009 ? 4'h9 : add_72409[3:0]];
  assign array_index_72413 = array_update_72410[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_72417 = smul32b_32b_x_32b(array_index_72024[add_72409 > 32'h0000_0009 ? 4'h9 : add_72409[3:0]], array_index_72412[add_72290 > 32'h0000_0009 ? 4'h9 : add_72290[3:0]]);
  assign add_72419 = array_index_72413[add_72290 > 32'h0000_0009 ? 4'h9 : add_72290[3:0]] + smul_72417;
  assign array_update_72420[0] = add_72290 == 32'h0000_0000 ? add_72419 : array_index_72413[0];
  assign array_update_72420[1] = add_72290 == 32'h0000_0001 ? add_72419 : array_index_72413[1];
  assign array_update_72420[2] = add_72290 == 32'h0000_0002 ? add_72419 : array_index_72413[2];
  assign array_update_72420[3] = add_72290 == 32'h0000_0003 ? add_72419 : array_index_72413[3];
  assign array_update_72420[4] = add_72290 == 32'h0000_0004 ? add_72419 : array_index_72413[4];
  assign array_update_72420[5] = add_72290 == 32'h0000_0005 ? add_72419 : array_index_72413[5];
  assign array_update_72420[6] = add_72290 == 32'h0000_0006 ? add_72419 : array_index_72413[6];
  assign array_update_72420[7] = add_72290 == 32'h0000_0007 ? add_72419 : array_index_72413[7];
  assign array_update_72420[8] = add_72290 == 32'h0000_0008 ? add_72419 : array_index_72413[8];
  assign array_update_72420[9] = add_72290 == 32'h0000_0009 ? add_72419 : array_index_72413[9];
  assign array_update_72421[0] = literal_72009 == 32'h0000_0000 ? array_update_72420 : array_update_72410[0];
  assign array_update_72421[1] = literal_72009 == 32'h0000_0001 ? array_update_72420 : array_update_72410[1];
  assign array_update_72421[2] = literal_72009 == 32'h0000_0002 ? array_update_72420 : array_update_72410[2];
  assign array_update_72421[3] = literal_72009 == 32'h0000_0003 ? array_update_72420 : array_update_72410[3];
  assign array_update_72421[4] = literal_72009 == 32'h0000_0004 ? array_update_72420 : array_update_72410[4];
  assign array_update_72421[5] = literal_72009 == 32'h0000_0005 ? array_update_72420 : array_update_72410[5];
  assign array_update_72421[6] = literal_72009 == 32'h0000_0006 ? array_update_72420 : array_update_72410[6];
  assign array_update_72421[7] = literal_72009 == 32'h0000_0007 ? array_update_72420 : array_update_72410[7];
  assign array_update_72421[8] = literal_72009 == 32'h0000_0008 ? array_update_72420 : array_update_72410[8];
  assign array_update_72421[9] = literal_72009 == 32'h0000_0009 ? array_update_72420 : array_update_72410[9];
  assign array_index_72423 = array_update_72421[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign add_72425 = add_72290 + 32'h0000_0001;
  assign array_update_72426[0] = add_72425 == 32'h0000_0000 ? 32'h0000_0000 : array_index_72423[0];
  assign array_update_72426[1] = add_72425 == 32'h0000_0001 ? 32'h0000_0000 : array_index_72423[1];
  assign array_update_72426[2] = add_72425 == 32'h0000_0002 ? 32'h0000_0000 : array_index_72423[2];
  assign array_update_72426[3] = add_72425 == 32'h0000_0003 ? 32'h0000_0000 : array_index_72423[3];
  assign array_update_72426[4] = add_72425 == 32'h0000_0004 ? 32'h0000_0000 : array_index_72423[4];
  assign array_update_72426[5] = add_72425 == 32'h0000_0005 ? 32'h0000_0000 : array_index_72423[5];
  assign array_update_72426[6] = add_72425 == 32'h0000_0006 ? 32'h0000_0000 : array_index_72423[6];
  assign array_update_72426[7] = add_72425 == 32'h0000_0007 ? 32'h0000_0000 : array_index_72423[7];
  assign array_update_72426[8] = add_72425 == 32'h0000_0008 ? 32'h0000_0000 : array_index_72423[8];
  assign array_update_72426[9] = add_72425 == 32'h0000_0009 ? 32'h0000_0000 : array_index_72423[9];
  assign literal_72427 = 32'h0000_0000;
  assign array_update_72428[0] = literal_72009 == 32'h0000_0000 ? array_update_72426 : array_update_72421[0];
  assign array_update_72428[1] = literal_72009 == 32'h0000_0001 ? array_update_72426 : array_update_72421[1];
  assign array_update_72428[2] = literal_72009 == 32'h0000_0002 ? array_update_72426 : array_update_72421[2];
  assign array_update_72428[3] = literal_72009 == 32'h0000_0003 ? array_update_72426 : array_update_72421[3];
  assign array_update_72428[4] = literal_72009 == 32'h0000_0004 ? array_update_72426 : array_update_72421[4];
  assign array_update_72428[5] = literal_72009 == 32'h0000_0005 ? array_update_72426 : array_update_72421[5];
  assign array_update_72428[6] = literal_72009 == 32'h0000_0006 ? array_update_72426 : array_update_72421[6];
  assign array_update_72428[7] = literal_72009 == 32'h0000_0007 ? array_update_72426 : array_update_72421[7];
  assign array_update_72428[8] = literal_72009 == 32'h0000_0008 ? array_update_72426 : array_update_72421[8];
  assign array_update_72428[9] = literal_72009 == 32'h0000_0009 ? array_update_72426 : array_update_72421[9];
  assign array_index_72430 = array_update_72021[literal_72427 > 32'h0000_0009 ? 4'h9 : literal_72427[3:0]];
  assign array_index_72431 = array_update_72428[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_72435 = smul32b_32b_x_32b(array_index_72024[literal_72427 > 32'h0000_0009 ? 4'h9 : literal_72427[3:0]], array_index_72430[add_72425 > 32'h0000_0009 ? 4'h9 : add_72425[3:0]]);
  assign add_72437 = array_index_72431[add_72425 > 32'h0000_0009 ? 4'h9 : add_72425[3:0]] + smul_72435;
  assign array_update_72439[0] = add_72425 == 32'h0000_0000 ? add_72437 : array_index_72431[0];
  assign array_update_72439[1] = add_72425 == 32'h0000_0001 ? add_72437 : array_index_72431[1];
  assign array_update_72439[2] = add_72425 == 32'h0000_0002 ? add_72437 : array_index_72431[2];
  assign array_update_72439[3] = add_72425 == 32'h0000_0003 ? add_72437 : array_index_72431[3];
  assign array_update_72439[4] = add_72425 == 32'h0000_0004 ? add_72437 : array_index_72431[4];
  assign array_update_72439[5] = add_72425 == 32'h0000_0005 ? add_72437 : array_index_72431[5];
  assign array_update_72439[6] = add_72425 == 32'h0000_0006 ? add_72437 : array_index_72431[6];
  assign array_update_72439[7] = add_72425 == 32'h0000_0007 ? add_72437 : array_index_72431[7];
  assign array_update_72439[8] = add_72425 == 32'h0000_0008 ? add_72437 : array_index_72431[8];
  assign array_update_72439[9] = add_72425 == 32'h0000_0009 ? add_72437 : array_index_72431[9];
  assign add_72440 = literal_72427 + 32'h0000_0001;
  assign array_update_72441[0] = literal_72009 == 32'h0000_0000 ? array_update_72439 : array_update_72428[0];
  assign array_update_72441[1] = literal_72009 == 32'h0000_0001 ? array_update_72439 : array_update_72428[1];
  assign array_update_72441[2] = literal_72009 == 32'h0000_0002 ? array_update_72439 : array_update_72428[2];
  assign array_update_72441[3] = literal_72009 == 32'h0000_0003 ? array_update_72439 : array_update_72428[3];
  assign array_update_72441[4] = literal_72009 == 32'h0000_0004 ? array_update_72439 : array_update_72428[4];
  assign array_update_72441[5] = literal_72009 == 32'h0000_0005 ? array_update_72439 : array_update_72428[5];
  assign array_update_72441[6] = literal_72009 == 32'h0000_0006 ? array_update_72439 : array_update_72428[6];
  assign array_update_72441[7] = literal_72009 == 32'h0000_0007 ? array_update_72439 : array_update_72428[7];
  assign array_update_72441[8] = literal_72009 == 32'h0000_0008 ? array_update_72439 : array_update_72428[8];
  assign array_update_72441[9] = literal_72009 == 32'h0000_0009 ? array_update_72439 : array_update_72428[9];
  assign array_index_72443 = array_update_72021[add_72440 > 32'h0000_0009 ? 4'h9 : add_72440[3:0]];
  assign array_index_72444 = array_update_72441[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_72448 = smul32b_32b_x_32b(array_index_72024[add_72440 > 32'h0000_0009 ? 4'h9 : add_72440[3:0]], array_index_72443[add_72425 > 32'h0000_0009 ? 4'h9 : add_72425[3:0]]);
  assign add_72450 = array_index_72444[add_72425 > 32'h0000_0009 ? 4'h9 : add_72425[3:0]] + smul_72448;
  assign array_update_72452[0] = add_72425 == 32'h0000_0000 ? add_72450 : array_index_72444[0];
  assign array_update_72452[1] = add_72425 == 32'h0000_0001 ? add_72450 : array_index_72444[1];
  assign array_update_72452[2] = add_72425 == 32'h0000_0002 ? add_72450 : array_index_72444[2];
  assign array_update_72452[3] = add_72425 == 32'h0000_0003 ? add_72450 : array_index_72444[3];
  assign array_update_72452[4] = add_72425 == 32'h0000_0004 ? add_72450 : array_index_72444[4];
  assign array_update_72452[5] = add_72425 == 32'h0000_0005 ? add_72450 : array_index_72444[5];
  assign array_update_72452[6] = add_72425 == 32'h0000_0006 ? add_72450 : array_index_72444[6];
  assign array_update_72452[7] = add_72425 == 32'h0000_0007 ? add_72450 : array_index_72444[7];
  assign array_update_72452[8] = add_72425 == 32'h0000_0008 ? add_72450 : array_index_72444[8];
  assign array_update_72452[9] = add_72425 == 32'h0000_0009 ? add_72450 : array_index_72444[9];
  assign add_72453 = add_72440 + 32'h0000_0001;
  assign array_update_72454[0] = literal_72009 == 32'h0000_0000 ? array_update_72452 : array_update_72441[0];
  assign array_update_72454[1] = literal_72009 == 32'h0000_0001 ? array_update_72452 : array_update_72441[1];
  assign array_update_72454[2] = literal_72009 == 32'h0000_0002 ? array_update_72452 : array_update_72441[2];
  assign array_update_72454[3] = literal_72009 == 32'h0000_0003 ? array_update_72452 : array_update_72441[3];
  assign array_update_72454[4] = literal_72009 == 32'h0000_0004 ? array_update_72452 : array_update_72441[4];
  assign array_update_72454[5] = literal_72009 == 32'h0000_0005 ? array_update_72452 : array_update_72441[5];
  assign array_update_72454[6] = literal_72009 == 32'h0000_0006 ? array_update_72452 : array_update_72441[6];
  assign array_update_72454[7] = literal_72009 == 32'h0000_0007 ? array_update_72452 : array_update_72441[7];
  assign array_update_72454[8] = literal_72009 == 32'h0000_0008 ? array_update_72452 : array_update_72441[8];
  assign array_update_72454[9] = literal_72009 == 32'h0000_0009 ? array_update_72452 : array_update_72441[9];
  assign array_index_72456 = array_update_72021[add_72453 > 32'h0000_0009 ? 4'h9 : add_72453[3:0]];
  assign array_index_72457 = array_update_72454[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_72461 = smul32b_32b_x_32b(array_index_72024[add_72453 > 32'h0000_0009 ? 4'h9 : add_72453[3:0]], array_index_72456[add_72425 > 32'h0000_0009 ? 4'h9 : add_72425[3:0]]);
  assign add_72463 = array_index_72457[add_72425 > 32'h0000_0009 ? 4'h9 : add_72425[3:0]] + smul_72461;
  assign array_update_72465[0] = add_72425 == 32'h0000_0000 ? add_72463 : array_index_72457[0];
  assign array_update_72465[1] = add_72425 == 32'h0000_0001 ? add_72463 : array_index_72457[1];
  assign array_update_72465[2] = add_72425 == 32'h0000_0002 ? add_72463 : array_index_72457[2];
  assign array_update_72465[3] = add_72425 == 32'h0000_0003 ? add_72463 : array_index_72457[3];
  assign array_update_72465[4] = add_72425 == 32'h0000_0004 ? add_72463 : array_index_72457[4];
  assign array_update_72465[5] = add_72425 == 32'h0000_0005 ? add_72463 : array_index_72457[5];
  assign array_update_72465[6] = add_72425 == 32'h0000_0006 ? add_72463 : array_index_72457[6];
  assign array_update_72465[7] = add_72425 == 32'h0000_0007 ? add_72463 : array_index_72457[7];
  assign array_update_72465[8] = add_72425 == 32'h0000_0008 ? add_72463 : array_index_72457[8];
  assign array_update_72465[9] = add_72425 == 32'h0000_0009 ? add_72463 : array_index_72457[9];
  assign add_72466 = add_72453 + 32'h0000_0001;
  assign array_update_72467[0] = literal_72009 == 32'h0000_0000 ? array_update_72465 : array_update_72454[0];
  assign array_update_72467[1] = literal_72009 == 32'h0000_0001 ? array_update_72465 : array_update_72454[1];
  assign array_update_72467[2] = literal_72009 == 32'h0000_0002 ? array_update_72465 : array_update_72454[2];
  assign array_update_72467[3] = literal_72009 == 32'h0000_0003 ? array_update_72465 : array_update_72454[3];
  assign array_update_72467[4] = literal_72009 == 32'h0000_0004 ? array_update_72465 : array_update_72454[4];
  assign array_update_72467[5] = literal_72009 == 32'h0000_0005 ? array_update_72465 : array_update_72454[5];
  assign array_update_72467[6] = literal_72009 == 32'h0000_0006 ? array_update_72465 : array_update_72454[6];
  assign array_update_72467[7] = literal_72009 == 32'h0000_0007 ? array_update_72465 : array_update_72454[7];
  assign array_update_72467[8] = literal_72009 == 32'h0000_0008 ? array_update_72465 : array_update_72454[8];
  assign array_update_72467[9] = literal_72009 == 32'h0000_0009 ? array_update_72465 : array_update_72454[9];
  assign array_index_72469 = array_update_72021[add_72466 > 32'h0000_0009 ? 4'h9 : add_72466[3:0]];
  assign array_index_72470 = array_update_72467[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_72474 = smul32b_32b_x_32b(array_index_72024[add_72466 > 32'h0000_0009 ? 4'h9 : add_72466[3:0]], array_index_72469[add_72425 > 32'h0000_0009 ? 4'h9 : add_72425[3:0]]);
  assign add_72476 = array_index_72470[add_72425 > 32'h0000_0009 ? 4'h9 : add_72425[3:0]] + smul_72474;
  assign array_update_72478[0] = add_72425 == 32'h0000_0000 ? add_72476 : array_index_72470[0];
  assign array_update_72478[1] = add_72425 == 32'h0000_0001 ? add_72476 : array_index_72470[1];
  assign array_update_72478[2] = add_72425 == 32'h0000_0002 ? add_72476 : array_index_72470[2];
  assign array_update_72478[3] = add_72425 == 32'h0000_0003 ? add_72476 : array_index_72470[3];
  assign array_update_72478[4] = add_72425 == 32'h0000_0004 ? add_72476 : array_index_72470[4];
  assign array_update_72478[5] = add_72425 == 32'h0000_0005 ? add_72476 : array_index_72470[5];
  assign array_update_72478[6] = add_72425 == 32'h0000_0006 ? add_72476 : array_index_72470[6];
  assign array_update_72478[7] = add_72425 == 32'h0000_0007 ? add_72476 : array_index_72470[7];
  assign array_update_72478[8] = add_72425 == 32'h0000_0008 ? add_72476 : array_index_72470[8];
  assign array_update_72478[9] = add_72425 == 32'h0000_0009 ? add_72476 : array_index_72470[9];
  assign add_72479 = add_72466 + 32'h0000_0001;
  assign array_update_72480[0] = literal_72009 == 32'h0000_0000 ? array_update_72478 : array_update_72467[0];
  assign array_update_72480[1] = literal_72009 == 32'h0000_0001 ? array_update_72478 : array_update_72467[1];
  assign array_update_72480[2] = literal_72009 == 32'h0000_0002 ? array_update_72478 : array_update_72467[2];
  assign array_update_72480[3] = literal_72009 == 32'h0000_0003 ? array_update_72478 : array_update_72467[3];
  assign array_update_72480[4] = literal_72009 == 32'h0000_0004 ? array_update_72478 : array_update_72467[4];
  assign array_update_72480[5] = literal_72009 == 32'h0000_0005 ? array_update_72478 : array_update_72467[5];
  assign array_update_72480[6] = literal_72009 == 32'h0000_0006 ? array_update_72478 : array_update_72467[6];
  assign array_update_72480[7] = literal_72009 == 32'h0000_0007 ? array_update_72478 : array_update_72467[7];
  assign array_update_72480[8] = literal_72009 == 32'h0000_0008 ? array_update_72478 : array_update_72467[8];
  assign array_update_72480[9] = literal_72009 == 32'h0000_0009 ? array_update_72478 : array_update_72467[9];
  assign array_index_72482 = array_update_72021[add_72479 > 32'h0000_0009 ? 4'h9 : add_72479[3:0]];
  assign array_index_72483 = array_update_72480[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_72487 = smul32b_32b_x_32b(array_index_72024[add_72479 > 32'h0000_0009 ? 4'h9 : add_72479[3:0]], array_index_72482[add_72425 > 32'h0000_0009 ? 4'h9 : add_72425[3:0]]);
  assign add_72489 = array_index_72483[add_72425 > 32'h0000_0009 ? 4'h9 : add_72425[3:0]] + smul_72487;
  assign array_update_72491[0] = add_72425 == 32'h0000_0000 ? add_72489 : array_index_72483[0];
  assign array_update_72491[1] = add_72425 == 32'h0000_0001 ? add_72489 : array_index_72483[1];
  assign array_update_72491[2] = add_72425 == 32'h0000_0002 ? add_72489 : array_index_72483[2];
  assign array_update_72491[3] = add_72425 == 32'h0000_0003 ? add_72489 : array_index_72483[3];
  assign array_update_72491[4] = add_72425 == 32'h0000_0004 ? add_72489 : array_index_72483[4];
  assign array_update_72491[5] = add_72425 == 32'h0000_0005 ? add_72489 : array_index_72483[5];
  assign array_update_72491[6] = add_72425 == 32'h0000_0006 ? add_72489 : array_index_72483[6];
  assign array_update_72491[7] = add_72425 == 32'h0000_0007 ? add_72489 : array_index_72483[7];
  assign array_update_72491[8] = add_72425 == 32'h0000_0008 ? add_72489 : array_index_72483[8];
  assign array_update_72491[9] = add_72425 == 32'h0000_0009 ? add_72489 : array_index_72483[9];
  assign add_72492 = add_72479 + 32'h0000_0001;
  assign array_update_72493[0] = literal_72009 == 32'h0000_0000 ? array_update_72491 : array_update_72480[0];
  assign array_update_72493[1] = literal_72009 == 32'h0000_0001 ? array_update_72491 : array_update_72480[1];
  assign array_update_72493[2] = literal_72009 == 32'h0000_0002 ? array_update_72491 : array_update_72480[2];
  assign array_update_72493[3] = literal_72009 == 32'h0000_0003 ? array_update_72491 : array_update_72480[3];
  assign array_update_72493[4] = literal_72009 == 32'h0000_0004 ? array_update_72491 : array_update_72480[4];
  assign array_update_72493[5] = literal_72009 == 32'h0000_0005 ? array_update_72491 : array_update_72480[5];
  assign array_update_72493[6] = literal_72009 == 32'h0000_0006 ? array_update_72491 : array_update_72480[6];
  assign array_update_72493[7] = literal_72009 == 32'h0000_0007 ? array_update_72491 : array_update_72480[7];
  assign array_update_72493[8] = literal_72009 == 32'h0000_0008 ? array_update_72491 : array_update_72480[8];
  assign array_update_72493[9] = literal_72009 == 32'h0000_0009 ? array_update_72491 : array_update_72480[9];
  assign array_index_72495 = array_update_72021[add_72492 > 32'h0000_0009 ? 4'h9 : add_72492[3:0]];
  assign array_index_72496 = array_update_72493[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_72500 = smul32b_32b_x_32b(array_index_72024[add_72492 > 32'h0000_0009 ? 4'h9 : add_72492[3:0]], array_index_72495[add_72425 > 32'h0000_0009 ? 4'h9 : add_72425[3:0]]);
  assign add_72502 = array_index_72496[add_72425 > 32'h0000_0009 ? 4'h9 : add_72425[3:0]] + smul_72500;
  assign array_update_72504[0] = add_72425 == 32'h0000_0000 ? add_72502 : array_index_72496[0];
  assign array_update_72504[1] = add_72425 == 32'h0000_0001 ? add_72502 : array_index_72496[1];
  assign array_update_72504[2] = add_72425 == 32'h0000_0002 ? add_72502 : array_index_72496[2];
  assign array_update_72504[3] = add_72425 == 32'h0000_0003 ? add_72502 : array_index_72496[3];
  assign array_update_72504[4] = add_72425 == 32'h0000_0004 ? add_72502 : array_index_72496[4];
  assign array_update_72504[5] = add_72425 == 32'h0000_0005 ? add_72502 : array_index_72496[5];
  assign array_update_72504[6] = add_72425 == 32'h0000_0006 ? add_72502 : array_index_72496[6];
  assign array_update_72504[7] = add_72425 == 32'h0000_0007 ? add_72502 : array_index_72496[7];
  assign array_update_72504[8] = add_72425 == 32'h0000_0008 ? add_72502 : array_index_72496[8];
  assign array_update_72504[9] = add_72425 == 32'h0000_0009 ? add_72502 : array_index_72496[9];
  assign add_72505 = add_72492 + 32'h0000_0001;
  assign array_update_72506[0] = literal_72009 == 32'h0000_0000 ? array_update_72504 : array_update_72493[0];
  assign array_update_72506[1] = literal_72009 == 32'h0000_0001 ? array_update_72504 : array_update_72493[1];
  assign array_update_72506[2] = literal_72009 == 32'h0000_0002 ? array_update_72504 : array_update_72493[2];
  assign array_update_72506[3] = literal_72009 == 32'h0000_0003 ? array_update_72504 : array_update_72493[3];
  assign array_update_72506[4] = literal_72009 == 32'h0000_0004 ? array_update_72504 : array_update_72493[4];
  assign array_update_72506[5] = literal_72009 == 32'h0000_0005 ? array_update_72504 : array_update_72493[5];
  assign array_update_72506[6] = literal_72009 == 32'h0000_0006 ? array_update_72504 : array_update_72493[6];
  assign array_update_72506[7] = literal_72009 == 32'h0000_0007 ? array_update_72504 : array_update_72493[7];
  assign array_update_72506[8] = literal_72009 == 32'h0000_0008 ? array_update_72504 : array_update_72493[8];
  assign array_update_72506[9] = literal_72009 == 32'h0000_0009 ? array_update_72504 : array_update_72493[9];
  assign array_index_72508 = array_update_72021[add_72505 > 32'h0000_0009 ? 4'h9 : add_72505[3:0]];
  assign array_index_72509 = array_update_72506[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_72513 = smul32b_32b_x_32b(array_index_72024[add_72505 > 32'h0000_0009 ? 4'h9 : add_72505[3:0]], array_index_72508[add_72425 > 32'h0000_0009 ? 4'h9 : add_72425[3:0]]);
  assign add_72515 = array_index_72509[add_72425 > 32'h0000_0009 ? 4'h9 : add_72425[3:0]] + smul_72513;
  assign array_update_72517[0] = add_72425 == 32'h0000_0000 ? add_72515 : array_index_72509[0];
  assign array_update_72517[1] = add_72425 == 32'h0000_0001 ? add_72515 : array_index_72509[1];
  assign array_update_72517[2] = add_72425 == 32'h0000_0002 ? add_72515 : array_index_72509[2];
  assign array_update_72517[3] = add_72425 == 32'h0000_0003 ? add_72515 : array_index_72509[3];
  assign array_update_72517[4] = add_72425 == 32'h0000_0004 ? add_72515 : array_index_72509[4];
  assign array_update_72517[5] = add_72425 == 32'h0000_0005 ? add_72515 : array_index_72509[5];
  assign array_update_72517[6] = add_72425 == 32'h0000_0006 ? add_72515 : array_index_72509[6];
  assign array_update_72517[7] = add_72425 == 32'h0000_0007 ? add_72515 : array_index_72509[7];
  assign array_update_72517[8] = add_72425 == 32'h0000_0008 ? add_72515 : array_index_72509[8];
  assign array_update_72517[9] = add_72425 == 32'h0000_0009 ? add_72515 : array_index_72509[9];
  assign add_72518 = add_72505 + 32'h0000_0001;
  assign array_update_72519[0] = literal_72009 == 32'h0000_0000 ? array_update_72517 : array_update_72506[0];
  assign array_update_72519[1] = literal_72009 == 32'h0000_0001 ? array_update_72517 : array_update_72506[1];
  assign array_update_72519[2] = literal_72009 == 32'h0000_0002 ? array_update_72517 : array_update_72506[2];
  assign array_update_72519[3] = literal_72009 == 32'h0000_0003 ? array_update_72517 : array_update_72506[3];
  assign array_update_72519[4] = literal_72009 == 32'h0000_0004 ? array_update_72517 : array_update_72506[4];
  assign array_update_72519[5] = literal_72009 == 32'h0000_0005 ? array_update_72517 : array_update_72506[5];
  assign array_update_72519[6] = literal_72009 == 32'h0000_0006 ? array_update_72517 : array_update_72506[6];
  assign array_update_72519[7] = literal_72009 == 32'h0000_0007 ? array_update_72517 : array_update_72506[7];
  assign array_update_72519[8] = literal_72009 == 32'h0000_0008 ? array_update_72517 : array_update_72506[8];
  assign array_update_72519[9] = literal_72009 == 32'h0000_0009 ? array_update_72517 : array_update_72506[9];
  assign array_index_72521 = array_update_72021[add_72518 > 32'h0000_0009 ? 4'h9 : add_72518[3:0]];
  assign array_index_72522 = array_update_72519[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_72526 = smul32b_32b_x_32b(array_index_72024[add_72518 > 32'h0000_0009 ? 4'h9 : add_72518[3:0]], array_index_72521[add_72425 > 32'h0000_0009 ? 4'h9 : add_72425[3:0]]);
  assign add_72528 = array_index_72522[add_72425 > 32'h0000_0009 ? 4'h9 : add_72425[3:0]] + smul_72526;
  assign array_update_72530[0] = add_72425 == 32'h0000_0000 ? add_72528 : array_index_72522[0];
  assign array_update_72530[1] = add_72425 == 32'h0000_0001 ? add_72528 : array_index_72522[1];
  assign array_update_72530[2] = add_72425 == 32'h0000_0002 ? add_72528 : array_index_72522[2];
  assign array_update_72530[3] = add_72425 == 32'h0000_0003 ? add_72528 : array_index_72522[3];
  assign array_update_72530[4] = add_72425 == 32'h0000_0004 ? add_72528 : array_index_72522[4];
  assign array_update_72530[5] = add_72425 == 32'h0000_0005 ? add_72528 : array_index_72522[5];
  assign array_update_72530[6] = add_72425 == 32'h0000_0006 ? add_72528 : array_index_72522[6];
  assign array_update_72530[7] = add_72425 == 32'h0000_0007 ? add_72528 : array_index_72522[7];
  assign array_update_72530[8] = add_72425 == 32'h0000_0008 ? add_72528 : array_index_72522[8];
  assign array_update_72530[9] = add_72425 == 32'h0000_0009 ? add_72528 : array_index_72522[9];
  assign add_72531 = add_72518 + 32'h0000_0001;
  assign array_update_72532[0] = literal_72009 == 32'h0000_0000 ? array_update_72530 : array_update_72519[0];
  assign array_update_72532[1] = literal_72009 == 32'h0000_0001 ? array_update_72530 : array_update_72519[1];
  assign array_update_72532[2] = literal_72009 == 32'h0000_0002 ? array_update_72530 : array_update_72519[2];
  assign array_update_72532[3] = literal_72009 == 32'h0000_0003 ? array_update_72530 : array_update_72519[3];
  assign array_update_72532[4] = literal_72009 == 32'h0000_0004 ? array_update_72530 : array_update_72519[4];
  assign array_update_72532[5] = literal_72009 == 32'h0000_0005 ? array_update_72530 : array_update_72519[5];
  assign array_update_72532[6] = literal_72009 == 32'h0000_0006 ? array_update_72530 : array_update_72519[6];
  assign array_update_72532[7] = literal_72009 == 32'h0000_0007 ? array_update_72530 : array_update_72519[7];
  assign array_update_72532[8] = literal_72009 == 32'h0000_0008 ? array_update_72530 : array_update_72519[8];
  assign array_update_72532[9] = literal_72009 == 32'h0000_0009 ? array_update_72530 : array_update_72519[9];
  assign array_index_72534 = array_update_72021[add_72531 > 32'h0000_0009 ? 4'h9 : add_72531[3:0]];
  assign array_index_72535 = array_update_72532[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_72539 = smul32b_32b_x_32b(array_index_72024[add_72531 > 32'h0000_0009 ? 4'h9 : add_72531[3:0]], array_index_72534[add_72425 > 32'h0000_0009 ? 4'h9 : add_72425[3:0]]);
  assign add_72541 = array_index_72535[add_72425 > 32'h0000_0009 ? 4'h9 : add_72425[3:0]] + smul_72539;
  assign array_update_72543[0] = add_72425 == 32'h0000_0000 ? add_72541 : array_index_72535[0];
  assign array_update_72543[1] = add_72425 == 32'h0000_0001 ? add_72541 : array_index_72535[1];
  assign array_update_72543[2] = add_72425 == 32'h0000_0002 ? add_72541 : array_index_72535[2];
  assign array_update_72543[3] = add_72425 == 32'h0000_0003 ? add_72541 : array_index_72535[3];
  assign array_update_72543[4] = add_72425 == 32'h0000_0004 ? add_72541 : array_index_72535[4];
  assign array_update_72543[5] = add_72425 == 32'h0000_0005 ? add_72541 : array_index_72535[5];
  assign array_update_72543[6] = add_72425 == 32'h0000_0006 ? add_72541 : array_index_72535[6];
  assign array_update_72543[7] = add_72425 == 32'h0000_0007 ? add_72541 : array_index_72535[7];
  assign array_update_72543[8] = add_72425 == 32'h0000_0008 ? add_72541 : array_index_72535[8];
  assign array_update_72543[9] = add_72425 == 32'h0000_0009 ? add_72541 : array_index_72535[9];
  assign add_72544 = add_72531 + 32'h0000_0001;
  assign array_update_72545[0] = literal_72009 == 32'h0000_0000 ? array_update_72543 : array_update_72532[0];
  assign array_update_72545[1] = literal_72009 == 32'h0000_0001 ? array_update_72543 : array_update_72532[1];
  assign array_update_72545[2] = literal_72009 == 32'h0000_0002 ? array_update_72543 : array_update_72532[2];
  assign array_update_72545[3] = literal_72009 == 32'h0000_0003 ? array_update_72543 : array_update_72532[3];
  assign array_update_72545[4] = literal_72009 == 32'h0000_0004 ? array_update_72543 : array_update_72532[4];
  assign array_update_72545[5] = literal_72009 == 32'h0000_0005 ? array_update_72543 : array_update_72532[5];
  assign array_update_72545[6] = literal_72009 == 32'h0000_0006 ? array_update_72543 : array_update_72532[6];
  assign array_update_72545[7] = literal_72009 == 32'h0000_0007 ? array_update_72543 : array_update_72532[7];
  assign array_update_72545[8] = literal_72009 == 32'h0000_0008 ? array_update_72543 : array_update_72532[8];
  assign array_update_72545[9] = literal_72009 == 32'h0000_0009 ? array_update_72543 : array_update_72532[9];
  assign array_index_72547 = array_update_72021[add_72544 > 32'h0000_0009 ? 4'h9 : add_72544[3:0]];
  assign array_index_72548 = array_update_72545[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_72552 = smul32b_32b_x_32b(array_index_72024[add_72544 > 32'h0000_0009 ? 4'h9 : add_72544[3:0]], array_index_72547[add_72425 > 32'h0000_0009 ? 4'h9 : add_72425[3:0]]);
  assign add_72554 = array_index_72548[add_72425 > 32'h0000_0009 ? 4'h9 : add_72425[3:0]] + smul_72552;
  assign array_update_72555[0] = add_72425 == 32'h0000_0000 ? add_72554 : array_index_72548[0];
  assign array_update_72555[1] = add_72425 == 32'h0000_0001 ? add_72554 : array_index_72548[1];
  assign array_update_72555[2] = add_72425 == 32'h0000_0002 ? add_72554 : array_index_72548[2];
  assign array_update_72555[3] = add_72425 == 32'h0000_0003 ? add_72554 : array_index_72548[3];
  assign array_update_72555[4] = add_72425 == 32'h0000_0004 ? add_72554 : array_index_72548[4];
  assign array_update_72555[5] = add_72425 == 32'h0000_0005 ? add_72554 : array_index_72548[5];
  assign array_update_72555[6] = add_72425 == 32'h0000_0006 ? add_72554 : array_index_72548[6];
  assign array_update_72555[7] = add_72425 == 32'h0000_0007 ? add_72554 : array_index_72548[7];
  assign array_update_72555[8] = add_72425 == 32'h0000_0008 ? add_72554 : array_index_72548[8];
  assign array_update_72555[9] = add_72425 == 32'h0000_0009 ? add_72554 : array_index_72548[9];
  assign array_update_72556[0] = literal_72009 == 32'h0000_0000 ? array_update_72555 : array_update_72545[0];
  assign array_update_72556[1] = literal_72009 == 32'h0000_0001 ? array_update_72555 : array_update_72545[1];
  assign array_update_72556[2] = literal_72009 == 32'h0000_0002 ? array_update_72555 : array_update_72545[2];
  assign array_update_72556[3] = literal_72009 == 32'h0000_0003 ? array_update_72555 : array_update_72545[3];
  assign array_update_72556[4] = literal_72009 == 32'h0000_0004 ? array_update_72555 : array_update_72545[4];
  assign array_update_72556[5] = literal_72009 == 32'h0000_0005 ? array_update_72555 : array_update_72545[5];
  assign array_update_72556[6] = literal_72009 == 32'h0000_0006 ? array_update_72555 : array_update_72545[6];
  assign array_update_72556[7] = literal_72009 == 32'h0000_0007 ? array_update_72555 : array_update_72545[7];
  assign array_update_72556[8] = literal_72009 == 32'h0000_0008 ? array_update_72555 : array_update_72545[8];
  assign array_update_72556[9] = literal_72009 == 32'h0000_0009 ? array_update_72555 : array_update_72545[9];
  assign array_index_72558 = array_update_72556[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign add_72560 = add_72425 + 32'h0000_0001;
  assign array_update_72561[0] = add_72560 == 32'h0000_0000 ? 32'h0000_0000 : array_index_72558[0];
  assign array_update_72561[1] = add_72560 == 32'h0000_0001 ? 32'h0000_0000 : array_index_72558[1];
  assign array_update_72561[2] = add_72560 == 32'h0000_0002 ? 32'h0000_0000 : array_index_72558[2];
  assign array_update_72561[3] = add_72560 == 32'h0000_0003 ? 32'h0000_0000 : array_index_72558[3];
  assign array_update_72561[4] = add_72560 == 32'h0000_0004 ? 32'h0000_0000 : array_index_72558[4];
  assign array_update_72561[5] = add_72560 == 32'h0000_0005 ? 32'h0000_0000 : array_index_72558[5];
  assign array_update_72561[6] = add_72560 == 32'h0000_0006 ? 32'h0000_0000 : array_index_72558[6];
  assign array_update_72561[7] = add_72560 == 32'h0000_0007 ? 32'h0000_0000 : array_index_72558[7];
  assign array_update_72561[8] = add_72560 == 32'h0000_0008 ? 32'h0000_0000 : array_index_72558[8];
  assign array_update_72561[9] = add_72560 == 32'h0000_0009 ? 32'h0000_0000 : array_index_72558[9];
  assign literal_72562 = 32'h0000_0000;
  assign array_update_72563[0] = literal_72009 == 32'h0000_0000 ? array_update_72561 : array_update_72556[0];
  assign array_update_72563[1] = literal_72009 == 32'h0000_0001 ? array_update_72561 : array_update_72556[1];
  assign array_update_72563[2] = literal_72009 == 32'h0000_0002 ? array_update_72561 : array_update_72556[2];
  assign array_update_72563[3] = literal_72009 == 32'h0000_0003 ? array_update_72561 : array_update_72556[3];
  assign array_update_72563[4] = literal_72009 == 32'h0000_0004 ? array_update_72561 : array_update_72556[4];
  assign array_update_72563[5] = literal_72009 == 32'h0000_0005 ? array_update_72561 : array_update_72556[5];
  assign array_update_72563[6] = literal_72009 == 32'h0000_0006 ? array_update_72561 : array_update_72556[6];
  assign array_update_72563[7] = literal_72009 == 32'h0000_0007 ? array_update_72561 : array_update_72556[7];
  assign array_update_72563[8] = literal_72009 == 32'h0000_0008 ? array_update_72561 : array_update_72556[8];
  assign array_update_72563[9] = literal_72009 == 32'h0000_0009 ? array_update_72561 : array_update_72556[9];
  assign array_index_72565 = array_update_72021[literal_72562 > 32'h0000_0009 ? 4'h9 : literal_72562[3:0]];
  assign array_index_72566 = array_update_72563[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_72570 = smul32b_32b_x_32b(array_index_72024[literal_72562 > 32'h0000_0009 ? 4'h9 : literal_72562[3:0]], array_index_72565[add_72560 > 32'h0000_0009 ? 4'h9 : add_72560[3:0]]);
  assign add_72572 = array_index_72566[add_72560 > 32'h0000_0009 ? 4'h9 : add_72560[3:0]] + smul_72570;
  assign array_update_72574[0] = add_72560 == 32'h0000_0000 ? add_72572 : array_index_72566[0];
  assign array_update_72574[1] = add_72560 == 32'h0000_0001 ? add_72572 : array_index_72566[1];
  assign array_update_72574[2] = add_72560 == 32'h0000_0002 ? add_72572 : array_index_72566[2];
  assign array_update_72574[3] = add_72560 == 32'h0000_0003 ? add_72572 : array_index_72566[3];
  assign array_update_72574[4] = add_72560 == 32'h0000_0004 ? add_72572 : array_index_72566[4];
  assign array_update_72574[5] = add_72560 == 32'h0000_0005 ? add_72572 : array_index_72566[5];
  assign array_update_72574[6] = add_72560 == 32'h0000_0006 ? add_72572 : array_index_72566[6];
  assign array_update_72574[7] = add_72560 == 32'h0000_0007 ? add_72572 : array_index_72566[7];
  assign array_update_72574[8] = add_72560 == 32'h0000_0008 ? add_72572 : array_index_72566[8];
  assign array_update_72574[9] = add_72560 == 32'h0000_0009 ? add_72572 : array_index_72566[9];
  assign add_72575 = literal_72562 + 32'h0000_0001;
  assign array_update_72576[0] = literal_72009 == 32'h0000_0000 ? array_update_72574 : array_update_72563[0];
  assign array_update_72576[1] = literal_72009 == 32'h0000_0001 ? array_update_72574 : array_update_72563[1];
  assign array_update_72576[2] = literal_72009 == 32'h0000_0002 ? array_update_72574 : array_update_72563[2];
  assign array_update_72576[3] = literal_72009 == 32'h0000_0003 ? array_update_72574 : array_update_72563[3];
  assign array_update_72576[4] = literal_72009 == 32'h0000_0004 ? array_update_72574 : array_update_72563[4];
  assign array_update_72576[5] = literal_72009 == 32'h0000_0005 ? array_update_72574 : array_update_72563[5];
  assign array_update_72576[6] = literal_72009 == 32'h0000_0006 ? array_update_72574 : array_update_72563[6];
  assign array_update_72576[7] = literal_72009 == 32'h0000_0007 ? array_update_72574 : array_update_72563[7];
  assign array_update_72576[8] = literal_72009 == 32'h0000_0008 ? array_update_72574 : array_update_72563[8];
  assign array_update_72576[9] = literal_72009 == 32'h0000_0009 ? array_update_72574 : array_update_72563[9];
  assign array_index_72578 = array_update_72021[add_72575 > 32'h0000_0009 ? 4'h9 : add_72575[3:0]];
  assign array_index_72579 = array_update_72576[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_72583 = smul32b_32b_x_32b(array_index_72024[add_72575 > 32'h0000_0009 ? 4'h9 : add_72575[3:0]], array_index_72578[add_72560 > 32'h0000_0009 ? 4'h9 : add_72560[3:0]]);
  assign add_72585 = array_index_72579[add_72560 > 32'h0000_0009 ? 4'h9 : add_72560[3:0]] + smul_72583;
  assign array_update_72587[0] = add_72560 == 32'h0000_0000 ? add_72585 : array_index_72579[0];
  assign array_update_72587[1] = add_72560 == 32'h0000_0001 ? add_72585 : array_index_72579[1];
  assign array_update_72587[2] = add_72560 == 32'h0000_0002 ? add_72585 : array_index_72579[2];
  assign array_update_72587[3] = add_72560 == 32'h0000_0003 ? add_72585 : array_index_72579[3];
  assign array_update_72587[4] = add_72560 == 32'h0000_0004 ? add_72585 : array_index_72579[4];
  assign array_update_72587[5] = add_72560 == 32'h0000_0005 ? add_72585 : array_index_72579[5];
  assign array_update_72587[6] = add_72560 == 32'h0000_0006 ? add_72585 : array_index_72579[6];
  assign array_update_72587[7] = add_72560 == 32'h0000_0007 ? add_72585 : array_index_72579[7];
  assign array_update_72587[8] = add_72560 == 32'h0000_0008 ? add_72585 : array_index_72579[8];
  assign array_update_72587[9] = add_72560 == 32'h0000_0009 ? add_72585 : array_index_72579[9];
  assign add_72588 = add_72575 + 32'h0000_0001;
  assign array_update_72589[0] = literal_72009 == 32'h0000_0000 ? array_update_72587 : array_update_72576[0];
  assign array_update_72589[1] = literal_72009 == 32'h0000_0001 ? array_update_72587 : array_update_72576[1];
  assign array_update_72589[2] = literal_72009 == 32'h0000_0002 ? array_update_72587 : array_update_72576[2];
  assign array_update_72589[3] = literal_72009 == 32'h0000_0003 ? array_update_72587 : array_update_72576[3];
  assign array_update_72589[4] = literal_72009 == 32'h0000_0004 ? array_update_72587 : array_update_72576[4];
  assign array_update_72589[5] = literal_72009 == 32'h0000_0005 ? array_update_72587 : array_update_72576[5];
  assign array_update_72589[6] = literal_72009 == 32'h0000_0006 ? array_update_72587 : array_update_72576[6];
  assign array_update_72589[7] = literal_72009 == 32'h0000_0007 ? array_update_72587 : array_update_72576[7];
  assign array_update_72589[8] = literal_72009 == 32'h0000_0008 ? array_update_72587 : array_update_72576[8];
  assign array_update_72589[9] = literal_72009 == 32'h0000_0009 ? array_update_72587 : array_update_72576[9];
  assign array_index_72591 = array_update_72021[add_72588 > 32'h0000_0009 ? 4'h9 : add_72588[3:0]];
  assign array_index_72592 = array_update_72589[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_72596 = smul32b_32b_x_32b(array_index_72024[add_72588 > 32'h0000_0009 ? 4'h9 : add_72588[3:0]], array_index_72591[add_72560 > 32'h0000_0009 ? 4'h9 : add_72560[3:0]]);
  assign add_72598 = array_index_72592[add_72560 > 32'h0000_0009 ? 4'h9 : add_72560[3:0]] + smul_72596;
  assign array_update_72600[0] = add_72560 == 32'h0000_0000 ? add_72598 : array_index_72592[0];
  assign array_update_72600[1] = add_72560 == 32'h0000_0001 ? add_72598 : array_index_72592[1];
  assign array_update_72600[2] = add_72560 == 32'h0000_0002 ? add_72598 : array_index_72592[2];
  assign array_update_72600[3] = add_72560 == 32'h0000_0003 ? add_72598 : array_index_72592[3];
  assign array_update_72600[4] = add_72560 == 32'h0000_0004 ? add_72598 : array_index_72592[4];
  assign array_update_72600[5] = add_72560 == 32'h0000_0005 ? add_72598 : array_index_72592[5];
  assign array_update_72600[6] = add_72560 == 32'h0000_0006 ? add_72598 : array_index_72592[6];
  assign array_update_72600[7] = add_72560 == 32'h0000_0007 ? add_72598 : array_index_72592[7];
  assign array_update_72600[8] = add_72560 == 32'h0000_0008 ? add_72598 : array_index_72592[8];
  assign array_update_72600[9] = add_72560 == 32'h0000_0009 ? add_72598 : array_index_72592[9];
  assign add_72601 = add_72588 + 32'h0000_0001;
  assign array_update_72602[0] = literal_72009 == 32'h0000_0000 ? array_update_72600 : array_update_72589[0];
  assign array_update_72602[1] = literal_72009 == 32'h0000_0001 ? array_update_72600 : array_update_72589[1];
  assign array_update_72602[2] = literal_72009 == 32'h0000_0002 ? array_update_72600 : array_update_72589[2];
  assign array_update_72602[3] = literal_72009 == 32'h0000_0003 ? array_update_72600 : array_update_72589[3];
  assign array_update_72602[4] = literal_72009 == 32'h0000_0004 ? array_update_72600 : array_update_72589[4];
  assign array_update_72602[5] = literal_72009 == 32'h0000_0005 ? array_update_72600 : array_update_72589[5];
  assign array_update_72602[6] = literal_72009 == 32'h0000_0006 ? array_update_72600 : array_update_72589[6];
  assign array_update_72602[7] = literal_72009 == 32'h0000_0007 ? array_update_72600 : array_update_72589[7];
  assign array_update_72602[8] = literal_72009 == 32'h0000_0008 ? array_update_72600 : array_update_72589[8];
  assign array_update_72602[9] = literal_72009 == 32'h0000_0009 ? array_update_72600 : array_update_72589[9];
  assign array_index_72604 = array_update_72021[add_72601 > 32'h0000_0009 ? 4'h9 : add_72601[3:0]];
  assign array_index_72605 = array_update_72602[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_72609 = smul32b_32b_x_32b(array_index_72024[add_72601 > 32'h0000_0009 ? 4'h9 : add_72601[3:0]], array_index_72604[add_72560 > 32'h0000_0009 ? 4'h9 : add_72560[3:0]]);
  assign add_72611 = array_index_72605[add_72560 > 32'h0000_0009 ? 4'h9 : add_72560[3:0]] + smul_72609;
  assign array_update_72613[0] = add_72560 == 32'h0000_0000 ? add_72611 : array_index_72605[0];
  assign array_update_72613[1] = add_72560 == 32'h0000_0001 ? add_72611 : array_index_72605[1];
  assign array_update_72613[2] = add_72560 == 32'h0000_0002 ? add_72611 : array_index_72605[2];
  assign array_update_72613[3] = add_72560 == 32'h0000_0003 ? add_72611 : array_index_72605[3];
  assign array_update_72613[4] = add_72560 == 32'h0000_0004 ? add_72611 : array_index_72605[4];
  assign array_update_72613[5] = add_72560 == 32'h0000_0005 ? add_72611 : array_index_72605[5];
  assign array_update_72613[6] = add_72560 == 32'h0000_0006 ? add_72611 : array_index_72605[6];
  assign array_update_72613[7] = add_72560 == 32'h0000_0007 ? add_72611 : array_index_72605[7];
  assign array_update_72613[8] = add_72560 == 32'h0000_0008 ? add_72611 : array_index_72605[8];
  assign array_update_72613[9] = add_72560 == 32'h0000_0009 ? add_72611 : array_index_72605[9];
  assign add_72614 = add_72601 + 32'h0000_0001;
  assign array_update_72615[0] = literal_72009 == 32'h0000_0000 ? array_update_72613 : array_update_72602[0];
  assign array_update_72615[1] = literal_72009 == 32'h0000_0001 ? array_update_72613 : array_update_72602[1];
  assign array_update_72615[2] = literal_72009 == 32'h0000_0002 ? array_update_72613 : array_update_72602[2];
  assign array_update_72615[3] = literal_72009 == 32'h0000_0003 ? array_update_72613 : array_update_72602[3];
  assign array_update_72615[4] = literal_72009 == 32'h0000_0004 ? array_update_72613 : array_update_72602[4];
  assign array_update_72615[5] = literal_72009 == 32'h0000_0005 ? array_update_72613 : array_update_72602[5];
  assign array_update_72615[6] = literal_72009 == 32'h0000_0006 ? array_update_72613 : array_update_72602[6];
  assign array_update_72615[7] = literal_72009 == 32'h0000_0007 ? array_update_72613 : array_update_72602[7];
  assign array_update_72615[8] = literal_72009 == 32'h0000_0008 ? array_update_72613 : array_update_72602[8];
  assign array_update_72615[9] = literal_72009 == 32'h0000_0009 ? array_update_72613 : array_update_72602[9];
  assign array_index_72617 = array_update_72021[add_72614 > 32'h0000_0009 ? 4'h9 : add_72614[3:0]];
  assign array_index_72618 = array_update_72615[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_72622 = smul32b_32b_x_32b(array_index_72024[add_72614 > 32'h0000_0009 ? 4'h9 : add_72614[3:0]], array_index_72617[add_72560 > 32'h0000_0009 ? 4'h9 : add_72560[3:0]]);
  assign add_72624 = array_index_72618[add_72560 > 32'h0000_0009 ? 4'h9 : add_72560[3:0]] + smul_72622;
  assign array_update_72626[0] = add_72560 == 32'h0000_0000 ? add_72624 : array_index_72618[0];
  assign array_update_72626[1] = add_72560 == 32'h0000_0001 ? add_72624 : array_index_72618[1];
  assign array_update_72626[2] = add_72560 == 32'h0000_0002 ? add_72624 : array_index_72618[2];
  assign array_update_72626[3] = add_72560 == 32'h0000_0003 ? add_72624 : array_index_72618[3];
  assign array_update_72626[4] = add_72560 == 32'h0000_0004 ? add_72624 : array_index_72618[4];
  assign array_update_72626[5] = add_72560 == 32'h0000_0005 ? add_72624 : array_index_72618[5];
  assign array_update_72626[6] = add_72560 == 32'h0000_0006 ? add_72624 : array_index_72618[6];
  assign array_update_72626[7] = add_72560 == 32'h0000_0007 ? add_72624 : array_index_72618[7];
  assign array_update_72626[8] = add_72560 == 32'h0000_0008 ? add_72624 : array_index_72618[8];
  assign array_update_72626[9] = add_72560 == 32'h0000_0009 ? add_72624 : array_index_72618[9];
  assign add_72627 = add_72614 + 32'h0000_0001;
  assign array_update_72628[0] = literal_72009 == 32'h0000_0000 ? array_update_72626 : array_update_72615[0];
  assign array_update_72628[1] = literal_72009 == 32'h0000_0001 ? array_update_72626 : array_update_72615[1];
  assign array_update_72628[2] = literal_72009 == 32'h0000_0002 ? array_update_72626 : array_update_72615[2];
  assign array_update_72628[3] = literal_72009 == 32'h0000_0003 ? array_update_72626 : array_update_72615[3];
  assign array_update_72628[4] = literal_72009 == 32'h0000_0004 ? array_update_72626 : array_update_72615[4];
  assign array_update_72628[5] = literal_72009 == 32'h0000_0005 ? array_update_72626 : array_update_72615[5];
  assign array_update_72628[6] = literal_72009 == 32'h0000_0006 ? array_update_72626 : array_update_72615[6];
  assign array_update_72628[7] = literal_72009 == 32'h0000_0007 ? array_update_72626 : array_update_72615[7];
  assign array_update_72628[8] = literal_72009 == 32'h0000_0008 ? array_update_72626 : array_update_72615[8];
  assign array_update_72628[9] = literal_72009 == 32'h0000_0009 ? array_update_72626 : array_update_72615[9];
  assign array_index_72630 = array_update_72021[add_72627 > 32'h0000_0009 ? 4'h9 : add_72627[3:0]];
  assign array_index_72631 = array_update_72628[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_72635 = smul32b_32b_x_32b(array_index_72024[add_72627 > 32'h0000_0009 ? 4'h9 : add_72627[3:0]], array_index_72630[add_72560 > 32'h0000_0009 ? 4'h9 : add_72560[3:0]]);
  assign add_72637 = array_index_72631[add_72560 > 32'h0000_0009 ? 4'h9 : add_72560[3:0]] + smul_72635;
  assign array_update_72639[0] = add_72560 == 32'h0000_0000 ? add_72637 : array_index_72631[0];
  assign array_update_72639[1] = add_72560 == 32'h0000_0001 ? add_72637 : array_index_72631[1];
  assign array_update_72639[2] = add_72560 == 32'h0000_0002 ? add_72637 : array_index_72631[2];
  assign array_update_72639[3] = add_72560 == 32'h0000_0003 ? add_72637 : array_index_72631[3];
  assign array_update_72639[4] = add_72560 == 32'h0000_0004 ? add_72637 : array_index_72631[4];
  assign array_update_72639[5] = add_72560 == 32'h0000_0005 ? add_72637 : array_index_72631[5];
  assign array_update_72639[6] = add_72560 == 32'h0000_0006 ? add_72637 : array_index_72631[6];
  assign array_update_72639[7] = add_72560 == 32'h0000_0007 ? add_72637 : array_index_72631[7];
  assign array_update_72639[8] = add_72560 == 32'h0000_0008 ? add_72637 : array_index_72631[8];
  assign array_update_72639[9] = add_72560 == 32'h0000_0009 ? add_72637 : array_index_72631[9];
  assign add_72640 = add_72627 + 32'h0000_0001;
  assign array_update_72641[0] = literal_72009 == 32'h0000_0000 ? array_update_72639 : array_update_72628[0];
  assign array_update_72641[1] = literal_72009 == 32'h0000_0001 ? array_update_72639 : array_update_72628[1];
  assign array_update_72641[2] = literal_72009 == 32'h0000_0002 ? array_update_72639 : array_update_72628[2];
  assign array_update_72641[3] = literal_72009 == 32'h0000_0003 ? array_update_72639 : array_update_72628[3];
  assign array_update_72641[4] = literal_72009 == 32'h0000_0004 ? array_update_72639 : array_update_72628[4];
  assign array_update_72641[5] = literal_72009 == 32'h0000_0005 ? array_update_72639 : array_update_72628[5];
  assign array_update_72641[6] = literal_72009 == 32'h0000_0006 ? array_update_72639 : array_update_72628[6];
  assign array_update_72641[7] = literal_72009 == 32'h0000_0007 ? array_update_72639 : array_update_72628[7];
  assign array_update_72641[8] = literal_72009 == 32'h0000_0008 ? array_update_72639 : array_update_72628[8];
  assign array_update_72641[9] = literal_72009 == 32'h0000_0009 ? array_update_72639 : array_update_72628[9];
  assign array_index_72643 = array_update_72021[add_72640 > 32'h0000_0009 ? 4'h9 : add_72640[3:0]];
  assign array_index_72644 = array_update_72641[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_72648 = smul32b_32b_x_32b(array_index_72024[add_72640 > 32'h0000_0009 ? 4'h9 : add_72640[3:0]], array_index_72643[add_72560 > 32'h0000_0009 ? 4'h9 : add_72560[3:0]]);
  assign add_72650 = array_index_72644[add_72560 > 32'h0000_0009 ? 4'h9 : add_72560[3:0]] + smul_72648;
  assign array_update_72652[0] = add_72560 == 32'h0000_0000 ? add_72650 : array_index_72644[0];
  assign array_update_72652[1] = add_72560 == 32'h0000_0001 ? add_72650 : array_index_72644[1];
  assign array_update_72652[2] = add_72560 == 32'h0000_0002 ? add_72650 : array_index_72644[2];
  assign array_update_72652[3] = add_72560 == 32'h0000_0003 ? add_72650 : array_index_72644[3];
  assign array_update_72652[4] = add_72560 == 32'h0000_0004 ? add_72650 : array_index_72644[4];
  assign array_update_72652[5] = add_72560 == 32'h0000_0005 ? add_72650 : array_index_72644[5];
  assign array_update_72652[6] = add_72560 == 32'h0000_0006 ? add_72650 : array_index_72644[6];
  assign array_update_72652[7] = add_72560 == 32'h0000_0007 ? add_72650 : array_index_72644[7];
  assign array_update_72652[8] = add_72560 == 32'h0000_0008 ? add_72650 : array_index_72644[8];
  assign array_update_72652[9] = add_72560 == 32'h0000_0009 ? add_72650 : array_index_72644[9];
  assign add_72653 = add_72640 + 32'h0000_0001;
  assign array_update_72654[0] = literal_72009 == 32'h0000_0000 ? array_update_72652 : array_update_72641[0];
  assign array_update_72654[1] = literal_72009 == 32'h0000_0001 ? array_update_72652 : array_update_72641[1];
  assign array_update_72654[2] = literal_72009 == 32'h0000_0002 ? array_update_72652 : array_update_72641[2];
  assign array_update_72654[3] = literal_72009 == 32'h0000_0003 ? array_update_72652 : array_update_72641[3];
  assign array_update_72654[4] = literal_72009 == 32'h0000_0004 ? array_update_72652 : array_update_72641[4];
  assign array_update_72654[5] = literal_72009 == 32'h0000_0005 ? array_update_72652 : array_update_72641[5];
  assign array_update_72654[6] = literal_72009 == 32'h0000_0006 ? array_update_72652 : array_update_72641[6];
  assign array_update_72654[7] = literal_72009 == 32'h0000_0007 ? array_update_72652 : array_update_72641[7];
  assign array_update_72654[8] = literal_72009 == 32'h0000_0008 ? array_update_72652 : array_update_72641[8];
  assign array_update_72654[9] = literal_72009 == 32'h0000_0009 ? array_update_72652 : array_update_72641[9];
  assign array_index_72656 = array_update_72021[add_72653 > 32'h0000_0009 ? 4'h9 : add_72653[3:0]];
  assign array_index_72657 = array_update_72654[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_72661 = smul32b_32b_x_32b(array_index_72024[add_72653 > 32'h0000_0009 ? 4'h9 : add_72653[3:0]], array_index_72656[add_72560 > 32'h0000_0009 ? 4'h9 : add_72560[3:0]]);
  assign add_72663 = array_index_72657[add_72560 > 32'h0000_0009 ? 4'h9 : add_72560[3:0]] + smul_72661;
  assign array_update_72665[0] = add_72560 == 32'h0000_0000 ? add_72663 : array_index_72657[0];
  assign array_update_72665[1] = add_72560 == 32'h0000_0001 ? add_72663 : array_index_72657[1];
  assign array_update_72665[2] = add_72560 == 32'h0000_0002 ? add_72663 : array_index_72657[2];
  assign array_update_72665[3] = add_72560 == 32'h0000_0003 ? add_72663 : array_index_72657[3];
  assign array_update_72665[4] = add_72560 == 32'h0000_0004 ? add_72663 : array_index_72657[4];
  assign array_update_72665[5] = add_72560 == 32'h0000_0005 ? add_72663 : array_index_72657[5];
  assign array_update_72665[6] = add_72560 == 32'h0000_0006 ? add_72663 : array_index_72657[6];
  assign array_update_72665[7] = add_72560 == 32'h0000_0007 ? add_72663 : array_index_72657[7];
  assign array_update_72665[8] = add_72560 == 32'h0000_0008 ? add_72663 : array_index_72657[8];
  assign array_update_72665[9] = add_72560 == 32'h0000_0009 ? add_72663 : array_index_72657[9];
  assign add_72666 = add_72653 + 32'h0000_0001;
  assign array_update_72667[0] = literal_72009 == 32'h0000_0000 ? array_update_72665 : array_update_72654[0];
  assign array_update_72667[1] = literal_72009 == 32'h0000_0001 ? array_update_72665 : array_update_72654[1];
  assign array_update_72667[2] = literal_72009 == 32'h0000_0002 ? array_update_72665 : array_update_72654[2];
  assign array_update_72667[3] = literal_72009 == 32'h0000_0003 ? array_update_72665 : array_update_72654[3];
  assign array_update_72667[4] = literal_72009 == 32'h0000_0004 ? array_update_72665 : array_update_72654[4];
  assign array_update_72667[5] = literal_72009 == 32'h0000_0005 ? array_update_72665 : array_update_72654[5];
  assign array_update_72667[6] = literal_72009 == 32'h0000_0006 ? array_update_72665 : array_update_72654[6];
  assign array_update_72667[7] = literal_72009 == 32'h0000_0007 ? array_update_72665 : array_update_72654[7];
  assign array_update_72667[8] = literal_72009 == 32'h0000_0008 ? array_update_72665 : array_update_72654[8];
  assign array_update_72667[9] = literal_72009 == 32'h0000_0009 ? array_update_72665 : array_update_72654[9];
  assign array_index_72669 = array_update_72021[add_72666 > 32'h0000_0009 ? 4'h9 : add_72666[3:0]];
  assign array_index_72670 = array_update_72667[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_72674 = smul32b_32b_x_32b(array_index_72024[add_72666 > 32'h0000_0009 ? 4'h9 : add_72666[3:0]], array_index_72669[add_72560 > 32'h0000_0009 ? 4'h9 : add_72560[3:0]]);
  assign add_72676 = array_index_72670[add_72560 > 32'h0000_0009 ? 4'h9 : add_72560[3:0]] + smul_72674;
  assign array_update_72678[0] = add_72560 == 32'h0000_0000 ? add_72676 : array_index_72670[0];
  assign array_update_72678[1] = add_72560 == 32'h0000_0001 ? add_72676 : array_index_72670[1];
  assign array_update_72678[2] = add_72560 == 32'h0000_0002 ? add_72676 : array_index_72670[2];
  assign array_update_72678[3] = add_72560 == 32'h0000_0003 ? add_72676 : array_index_72670[3];
  assign array_update_72678[4] = add_72560 == 32'h0000_0004 ? add_72676 : array_index_72670[4];
  assign array_update_72678[5] = add_72560 == 32'h0000_0005 ? add_72676 : array_index_72670[5];
  assign array_update_72678[6] = add_72560 == 32'h0000_0006 ? add_72676 : array_index_72670[6];
  assign array_update_72678[7] = add_72560 == 32'h0000_0007 ? add_72676 : array_index_72670[7];
  assign array_update_72678[8] = add_72560 == 32'h0000_0008 ? add_72676 : array_index_72670[8];
  assign array_update_72678[9] = add_72560 == 32'h0000_0009 ? add_72676 : array_index_72670[9];
  assign add_72679 = add_72666 + 32'h0000_0001;
  assign array_update_72680[0] = literal_72009 == 32'h0000_0000 ? array_update_72678 : array_update_72667[0];
  assign array_update_72680[1] = literal_72009 == 32'h0000_0001 ? array_update_72678 : array_update_72667[1];
  assign array_update_72680[2] = literal_72009 == 32'h0000_0002 ? array_update_72678 : array_update_72667[2];
  assign array_update_72680[3] = literal_72009 == 32'h0000_0003 ? array_update_72678 : array_update_72667[3];
  assign array_update_72680[4] = literal_72009 == 32'h0000_0004 ? array_update_72678 : array_update_72667[4];
  assign array_update_72680[5] = literal_72009 == 32'h0000_0005 ? array_update_72678 : array_update_72667[5];
  assign array_update_72680[6] = literal_72009 == 32'h0000_0006 ? array_update_72678 : array_update_72667[6];
  assign array_update_72680[7] = literal_72009 == 32'h0000_0007 ? array_update_72678 : array_update_72667[7];
  assign array_update_72680[8] = literal_72009 == 32'h0000_0008 ? array_update_72678 : array_update_72667[8];
  assign array_update_72680[9] = literal_72009 == 32'h0000_0009 ? array_update_72678 : array_update_72667[9];
  assign array_index_72682 = array_update_72021[add_72679 > 32'h0000_0009 ? 4'h9 : add_72679[3:0]];
  assign array_index_72683 = array_update_72680[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_72687 = smul32b_32b_x_32b(array_index_72024[add_72679 > 32'h0000_0009 ? 4'h9 : add_72679[3:0]], array_index_72682[add_72560 > 32'h0000_0009 ? 4'h9 : add_72560[3:0]]);
  assign add_72689 = array_index_72683[add_72560 > 32'h0000_0009 ? 4'h9 : add_72560[3:0]] + smul_72687;
  assign array_update_72690[0] = add_72560 == 32'h0000_0000 ? add_72689 : array_index_72683[0];
  assign array_update_72690[1] = add_72560 == 32'h0000_0001 ? add_72689 : array_index_72683[1];
  assign array_update_72690[2] = add_72560 == 32'h0000_0002 ? add_72689 : array_index_72683[2];
  assign array_update_72690[3] = add_72560 == 32'h0000_0003 ? add_72689 : array_index_72683[3];
  assign array_update_72690[4] = add_72560 == 32'h0000_0004 ? add_72689 : array_index_72683[4];
  assign array_update_72690[5] = add_72560 == 32'h0000_0005 ? add_72689 : array_index_72683[5];
  assign array_update_72690[6] = add_72560 == 32'h0000_0006 ? add_72689 : array_index_72683[6];
  assign array_update_72690[7] = add_72560 == 32'h0000_0007 ? add_72689 : array_index_72683[7];
  assign array_update_72690[8] = add_72560 == 32'h0000_0008 ? add_72689 : array_index_72683[8];
  assign array_update_72690[9] = add_72560 == 32'h0000_0009 ? add_72689 : array_index_72683[9];
  assign array_update_72691[0] = literal_72009 == 32'h0000_0000 ? array_update_72690 : array_update_72680[0];
  assign array_update_72691[1] = literal_72009 == 32'h0000_0001 ? array_update_72690 : array_update_72680[1];
  assign array_update_72691[2] = literal_72009 == 32'h0000_0002 ? array_update_72690 : array_update_72680[2];
  assign array_update_72691[3] = literal_72009 == 32'h0000_0003 ? array_update_72690 : array_update_72680[3];
  assign array_update_72691[4] = literal_72009 == 32'h0000_0004 ? array_update_72690 : array_update_72680[4];
  assign array_update_72691[5] = literal_72009 == 32'h0000_0005 ? array_update_72690 : array_update_72680[5];
  assign array_update_72691[6] = literal_72009 == 32'h0000_0006 ? array_update_72690 : array_update_72680[6];
  assign array_update_72691[7] = literal_72009 == 32'h0000_0007 ? array_update_72690 : array_update_72680[7];
  assign array_update_72691[8] = literal_72009 == 32'h0000_0008 ? array_update_72690 : array_update_72680[8];
  assign array_update_72691[9] = literal_72009 == 32'h0000_0009 ? array_update_72690 : array_update_72680[9];
  assign array_index_72693 = array_update_72691[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign add_72695 = add_72560 + 32'h0000_0001;
  assign array_update_72696[0] = add_72695 == 32'h0000_0000 ? 32'h0000_0000 : array_index_72693[0];
  assign array_update_72696[1] = add_72695 == 32'h0000_0001 ? 32'h0000_0000 : array_index_72693[1];
  assign array_update_72696[2] = add_72695 == 32'h0000_0002 ? 32'h0000_0000 : array_index_72693[2];
  assign array_update_72696[3] = add_72695 == 32'h0000_0003 ? 32'h0000_0000 : array_index_72693[3];
  assign array_update_72696[4] = add_72695 == 32'h0000_0004 ? 32'h0000_0000 : array_index_72693[4];
  assign array_update_72696[5] = add_72695 == 32'h0000_0005 ? 32'h0000_0000 : array_index_72693[5];
  assign array_update_72696[6] = add_72695 == 32'h0000_0006 ? 32'h0000_0000 : array_index_72693[6];
  assign array_update_72696[7] = add_72695 == 32'h0000_0007 ? 32'h0000_0000 : array_index_72693[7];
  assign array_update_72696[8] = add_72695 == 32'h0000_0008 ? 32'h0000_0000 : array_index_72693[8];
  assign array_update_72696[9] = add_72695 == 32'h0000_0009 ? 32'h0000_0000 : array_index_72693[9];
  assign literal_72697 = 32'h0000_0000;
  assign array_update_72698[0] = literal_72009 == 32'h0000_0000 ? array_update_72696 : array_update_72691[0];
  assign array_update_72698[1] = literal_72009 == 32'h0000_0001 ? array_update_72696 : array_update_72691[1];
  assign array_update_72698[2] = literal_72009 == 32'h0000_0002 ? array_update_72696 : array_update_72691[2];
  assign array_update_72698[3] = literal_72009 == 32'h0000_0003 ? array_update_72696 : array_update_72691[3];
  assign array_update_72698[4] = literal_72009 == 32'h0000_0004 ? array_update_72696 : array_update_72691[4];
  assign array_update_72698[5] = literal_72009 == 32'h0000_0005 ? array_update_72696 : array_update_72691[5];
  assign array_update_72698[6] = literal_72009 == 32'h0000_0006 ? array_update_72696 : array_update_72691[6];
  assign array_update_72698[7] = literal_72009 == 32'h0000_0007 ? array_update_72696 : array_update_72691[7];
  assign array_update_72698[8] = literal_72009 == 32'h0000_0008 ? array_update_72696 : array_update_72691[8];
  assign array_update_72698[9] = literal_72009 == 32'h0000_0009 ? array_update_72696 : array_update_72691[9];
  assign array_index_72700 = array_update_72021[literal_72697 > 32'h0000_0009 ? 4'h9 : literal_72697[3:0]];
  assign array_index_72701 = array_update_72698[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_72705 = smul32b_32b_x_32b(array_index_72024[literal_72697 > 32'h0000_0009 ? 4'h9 : literal_72697[3:0]], array_index_72700[add_72695 > 32'h0000_0009 ? 4'h9 : add_72695[3:0]]);
  assign add_72707 = array_index_72701[add_72695 > 32'h0000_0009 ? 4'h9 : add_72695[3:0]] + smul_72705;
  assign array_update_72709[0] = add_72695 == 32'h0000_0000 ? add_72707 : array_index_72701[0];
  assign array_update_72709[1] = add_72695 == 32'h0000_0001 ? add_72707 : array_index_72701[1];
  assign array_update_72709[2] = add_72695 == 32'h0000_0002 ? add_72707 : array_index_72701[2];
  assign array_update_72709[3] = add_72695 == 32'h0000_0003 ? add_72707 : array_index_72701[3];
  assign array_update_72709[4] = add_72695 == 32'h0000_0004 ? add_72707 : array_index_72701[4];
  assign array_update_72709[5] = add_72695 == 32'h0000_0005 ? add_72707 : array_index_72701[5];
  assign array_update_72709[6] = add_72695 == 32'h0000_0006 ? add_72707 : array_index_72701[6];
  assign array_update_72709[7] = add_72695 == 32'h0000_0007 ? add_72707 : array_index_72701[7];
  assign array_update_72709[8] = add_72695 == 32'h0000_0008 ? add_72707 : array_index_72701[8];
  assign array_update_72709[9] = add_72695 == 32'h0000_0009 ? add_72707 : array_index_72701[9];
  assign add_72710 = literal_72697 + 32'h0000_0001;
  assign array_update_72711[0] = literal_72009 == 32'h0000_0000 ? array_update_72709 : array_update_72698[0];
  assign array_update_72711[1] = literal_72009 == 32'h0000_0001 ? array_update_72709 : array_update_72698[1];
  assign array_update_72711[2] = literal_72009 == 32'h0000_0002 ? array_update_72709 : array_update_72698[2];
  assign array_update_72711[3] = literal_72009 == 32'h0000_0003 ? array_update_72709 : array_update_72698[3];
  assign array_update_72711[4] = literal_72009 == 32'h0000_0004 ? array_update_72709 : array_update_72698[4];
  assign array_update_72711[5] = literal_72009 == 32'h0000_0005 ? array_update_72709 : array_update_72698[5];
  assign array_update_72711[6] = literal_72009 == 32'h0000_0006 ? array_update_72709 : array_update_72698[6];
  assign array_update_72711[7] = literal_72009 == 32'h0000_0007 ? array_update_72709 : array_update_72698[7];
  assign array_update_72711[8] = literal_72009 == 32'h0000_0008 ? array_update_72709 : array_update_72698[8];
  assign array_update_72711[9] = literal_72009 == 32'h0000_0009 ? array_update_72709 : array_update_72698[9];
  assign array_index_72713 = array_update_72021[add_72710 > 32'h0000_0009 ? 4'h9 : add_72710[3:0]];
  assign array_index_72714 = array_update_72711[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_72718 = smul32b_32b_x_32b(array_index_72024[add_72710 > 32'h0000_0009 ? 4'h9 : add_72710[3:0]], array_index_72713[add_72695 > 32'h0000_0009 ? 4'h9 : add_72695[3:0]]);
  assign add_72720 = array_index_72714[add_72695 > 32'h0000_0009 ? 4'h9 : add_72695[3:0]] + smul_72718;
  assign array_update_72722[0] = add_72695 == 32'h0000_0000 ? add_72720 : array_index_72714[0];
  assign array_update_72722[1] = add_72695 == 32'h0000_0001 ? add_72720 : array_index_72714[1];
  assign array_update_72722[2] = add_72695 == 32'h0000_0002 ? add_72720 : array_index_72714[2];
  assign array_update_72722[3] = add_72695 == 32'h0000_0003 ? add_72720 : array_index_72714[3];
  assign array_update_72722[4] = add_72695 == 32'h0000_0004 ? add_72720 : array_index_72714[4];
  assign array_update_72722[5] = add_72695 == 32'h0000_0005 ? add_72720 : array_index_72714[5];
  assign array_update_72722[6] = add_72695 == 32'h0000_0006 ? add_72720 : array_index_72714[6];
  assign array_update_72722[7] = add_72695 == 32'h0000_0007 ? add_72720 : array_index_72714[7];
  assign array_update_72722[8] = add_72695 == 32'h0000_0008 ? add_72720 : array_index_72714[8];
  assign array_update_72722[9] = add_72695 == 32'h0000_0009 ? add_72720 : array_index_72714[9];
  assign add_72723 = add_72710 + 32'h0000_0001;
  assign array_update_72724[0] = literal_72009 == 32'h0000_0000 ? array_update_72722 : array_update_72711[0];
  assign array_update_72724[1] = literal_72009 == 32'h0000_0001 ? array_update_72722 : array_update_72711[1];
  assign array_update_72724[2] = literal_72009 == 32'h0000_0002 ? array_update_72722 : array_update_72711[2];
  assign array_update_72724[3] = literal_72009 == 32'h0000_0003 ? array_update_72722 : array_update_72711[3];
  assign array_update_72724[4] = literal_72009 == 32'h0000_0004 ? array_update_72722 : array_update_72711[4];
  assign array_update_72724[5] = literal_72009 == 32'h0000_0005 ? array_update_72722 : array_update_72711[5];
  assign array_update_72724[6] = literal_72009 == 32'h0000_0006 ? array_update_72722 : array_update_72711[6];
  assign array_update_72724[7] = literal_72009 == 32'h0000_0007 ? array_update_72722 : array_update_72711[7];
  assign array_update_72724[8] = literal_72009 == 32'h0000_0008 ? array_update_72722 : array_update_72711[8];
  assign array_update_72724[9] = literal_72009 == 32'h0000_0009 ? array_update_72722 : array_update_72711[9];
  assign array_index_72726 = array_update_72021[add_72723 > 32'h0000_0009 ? 4'h9 : add_72723[3:0]];
  assign array_index_72727 = array_update_72724[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_72731 = smul32b_32b_x_32b(array_index_72024[add_72723 > 32'h0000_0009 ? 4'h9 : add_72723[3:0]], array_index_72726[add_72695 > 32'h0000_0009 ? 4'h9 : add_72695[3:0]]);
  assign add_72733 = array_index_72727[add_72695 > 32'h0000_0009 ? 4'h9 : add_72695[3:0]] + smul_72731;
  assign array_update_72735[0] = add_72695 == 32'h0000_0000 ? add_72733 : array_index_72727[0];
  assign array_update_72735[1] = add_72695 == 32'h0000_0001 ? add_72733 : array_index_72727[1];
  assign array_update_72735[2] = add_72695 == 32'h0000_0002 ? add_72733 : array_index_72727[2];
  assign array_update_72735[3] = add_72695 == 32'h0000_0003 ? add_72733 : array_index_72727[3];
  assign array_update_72735[4] = add_72695 == 32'h0000_0004 ? add_72733 : array_index_72727[4];
  assign array_update_72735[5] = add_72695 == 32'h0000_0005 ? add_72733 : array_index_72727[5];
  assign array_update_72735[6] = add_72695 == 32'h0000_0006 ? add_72733 : array_index_72727[6];
  assign array_update_72735[7] = add_72695 == 32'h0000_0007 ? add_72733 : array_index_72727[7];
  assign array_update_72735[8] = add_72695 == 32'h0000_0008 ? add_72733 : array_index_72727[8];
  assign array_update_72735[9] = add_72695 == 32'h0000_0009 ? add_72733 : array_index_72727[9];
  assign add_72736 = add_72723 + 32'h0000_0001;
  assign array_update_72737[0] = literal_72009 == 32'h0000_0000 ? array_update_72735 : array_update_72724[0];
  assign array_update_72737[1] = literal_72009 == 32'h0000_0001 ? array_update_72735 : array_update_72724[1];
  assign array_update_72737[2] = literal_72009 == 32'h0000_0002 ? array_update_72735 : array_update_72724[2];
  assign array_update_72737[3] = literal_72009 == 32'h0000_0003 ? array_update_72735 : array_update_72724[3];
  assign array_update_72737[4] = literal_72009 == 32'h0000_0004 ? array_update_72735 : array_update_72724[4];
  assign array_update_72737[5] = literal_72009 == 32'h0000_0005 ? array_update_72735 : array_update_72724[5];
  assign array_update_72737[6] = literal_72009 == 32'h0000_0006 ? array_update_72735 : array_update_72724[6];
  assign array_update_72737[7] = literal_72009 == 32'h0000_0007 ? array_update_72735 : array_update_72724[7];
  assign array_update_72737[8] = literal_72009 == 32'h0000_0008 ? array_update_72735 : array_update_72724[8];
  assign array_update_72737[9] = literal_72009 == 32'h0000_0009 ? array_update_72735 : array_update_72724[9];
  assign array_index_72739 = array_update_72021[add_72736 > 32'h0000_0009 ? 4'h9 : add_72736[3:0]];
  assign array_index_72740 = array_update_72737[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_72744 = smul32b_32b_x_32b(array_index_72024[add_72736 > 32'h0000_0009 ? 4'h9 : add_72736[3:0]], array_index_72739[add_72695 > 32'h0000_0009 ? 4'h9 : add_72695[3:0]]);
  assign add_72746 = array_index_72740[add_72695 > 32'h0000_0009 ? 4'h9 : add_72695[3:0]] + smul_72744;
  assign array_update_72748[0] = add_72695 == 32'h0000_0000 ? add_72746 : array_index_72740[0];
  assign array_update_72748[1] = add_72695 == 32'h0000_0001 ? add_72746 : array_index_72740[1];
  assign array_update_72748[2] = add_72695 == 32'h0000_0002 ? add_72746 : array_index_72740[2];
  assign array_update_72748[3] = add_72695 == 32'h0000_0003 ? add_72746 : array_index_72740[3];
  assign array_update_72748[4] = add_72695 == 32'h0000_0004 ? add_72746 : array_index_72740[4];
  assign array_update_72748[5] = add_72695 == 32'h0000_0005 ? add_72746 : array_index_72740[5];
  assign array_update_72748[6] = add_72695 == 32'h0000_0006 ? add_72746 : array_index_72740[6];
  assign array_update_72748[7] = add_72695 == 32'h0000_0007 ? add_72746 : array_index_72740[7];
  assign array_update_72748[8] = add_72695 == 32'h0000_0008 ? add_72746 : array_index_72740[8];
  assign array_update_72748[9] = add_72695 == 32'h0000_0009 ? add_72746 : array_index_72740[9];
  assign add_72749 = add_72736 + 32'h0000_0001;
  assign array_update_72750[0] = literal_72009 == 32'h0000_0000 ? array_update_72748 : array_update_72737[0];
  assign array_update_72750[1] = literal_72009 == 32'h0000_0001 ? array_update_72748 : array_update_72737[1];
  assign array_update_72750[2] = literal_72009 == 32'h0000_0002 ? array_update_72748 : array_update_72737[2];
  assign array_update_72750[3] = literal_72009 == 32'h0000_0003 ? array_update_72748 : array_update_72737[3];
  assign array_update_72750[4] = literal_72009 == 32'h0000_0004 ? array_update_72748 : array_update_72737[4];
  assign array_update_72750[5] = literal_72009 == 32'h0000_0005 ? array_update_72748 : array_update_72737[5];
  assign array_update_72750[6] = literal_72009 == 32'h0000_0006 ? array_update_72748 : array_update_72737[6];
  assign array_update_72750[7] = literal_72009 == 32'h0000_0007 ? array_update_72748 : array_update_72737[7];
  assign array_update_72750[8] = literal_72009 == 32'h0000_0008 ? array_update_72748 : array_update_72737[8];
  assign array_update_72750[9] = literal_72009 == 32'h0000_0009 ? array_update_72748 : array_update_72737[9];
  assign array_index_72752 = array_update_72021[add_72749 > 32'h0000_0009 ? 4'h9 : add_72749[3:0]];
  assign array_index_72753 = array_update_72750[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_72757 = smul32b_32b_x_32b(array_index_72024[add_72749 > 32'h0000_0009 ? 4'h9 : add_72749[3:0]], array_index_72752[add_72695 > 32'h0000_0009 ? 4'h9 : add_72695[3:0]]);
  assign add_72759 = array_index_72753[add_72695 > 32'h0000_0009 ? 4'h9 : add_72695[3:0]] + smul_72757;
  assign array_update_72761[0] = add_72695 == 32'h0000_0000 ? add_72759 : array_index_72753[0];
  assign array_update_72761[1] = add_72695 == 32'h0000_0001 ? add_72759 : array_index_72753[1];
  assign array_update_72761[2] = add_72695 == 32'h0000_0002 ? add_72759 : array_index_72753[2];
  assign array_update_72761[3] = add_72695 == 32'h0000_0003 ? add_72759 : array_index_72753[3];
  assign array_update_72761[4] = add_72695 == 32'h0000_0004 ? add_72759 : array_index_72753[4];
  assign array_update_72761[5] = add_72695 == 32'h0000_0005 ? add_72759 : array_index_72753[5];
  assign array_update_72761[6] = add_72695 == 32'h0000_0006 ? add_72759 : array_index_72753[6];
  assign array_update_72761[7] = add_72695 == 32'h0000_0007 ? add_72759 : array_index_72753[7];
  assign array_update_72761[8] = add_72695 == 32'h0000_0008 ? add_72759 : array_index_72753[8];
  assign array_update_72761[9] = add_72695 == 32'h0000_0009 ? add_72759 : array_index_72753[9];
  assign add_72762 = add_72749 + 32'h0000_0001;
  assign array_update_72763[0] = literal_72009 == 32'h0000_0000 ? array_update_72761 : array_update_72750[0];
  assign array_update_72763[1] = literal_72009 == 32'h0000_0001 ? array_update_72761 : array_update_72750[1];
  assign array_update_72763[2] = literal_72009 == 32'h0000_0002 ? array_update_72761 : array_update_72750[2];
  assign array_update_72763[3] = literal_72009 == 32'h0000_0003 ? array_update_72761 : array_update_72750[3];
  assign array_update_72763[4] = literal_72009 == 32'h0000_0004 ? array_update_72761 : array_update_72750[4];
  assign array_update_72763[5] = literal_72009 == 32'h0000_0005 ? array_update_72761 : array_update_72750[5];
  assign array_update_72763[6] = literal_72009 == 32'h0000_0006 ? array_update_72761 : array_update_72750[6];
  assign array_update_72763[7] = literal_72009 == 32'h0000_0007 ? array_update_72761 : array_update_72750[7];
  assign array_update_72763[8] = literal_72009 == 32'h0000_0008 ? array_update_72761 : array_update_72750[8];
  assign array_update_72763[9] = literal_72009 == 32'h0000_0009 ? array_update_72761 : array_update_72750[9];
  assign array_index_72765 = array_update_72021[add_72762 > 32'h0000_0009 ? 4'h9 : add_72762[3:0]];
  assign array_index_72766 = array_update_72763[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_72770 = smul32b_32b_x_32b(array_index_72024[add_72762 > 32'h0000_0009 ? 4'h9 : add_72762[3:0]], array_index_72765[add_72695 > 32'h0000_0009 ? 4'h9 : add_72695[3:0]]);
  assign add_72772 = array_index_72766[add_72695 > 32'h0000_0009 ? 4'h9 : add_72695[3:0]] + smul_72770;
  assign array_update_72774[0] = add_72695 == 32'h0000_0000 ? add_72772 : array_index_72766[0];
  assign array_update_72774[1] = add_72695 == 32'h0000_0001 ? add_72772 : array_index_72766[1];
  assign array_update_72774[2] = add_72695 == 32'h0000_0002 ? add_72772 : array_index_72766[2];
  assign array_update_72774[3] = add_72695 == 32'h0000_0003 ? add_72772 : array_index_72766[3];
  assign array_update_72774[4] = add_72695 == 32'h0000_0004 ? add_72772 : array_index_72766[4];
  assign array_update_72774[5] = add_72695 == 32'h0000_0005 ? add_72772 : array_index_72766[5];
  assign array_update_72774[6] = add_72695 == 32'h0000_0006 ? add_72772 : array_index_72766[6];
  assign array_update_72774[7] = add_72695 == 32'h0000_0007 ? add_72772 : array_index_72766[7];
  assign array_update_72774[8] = add_72695 == 32'h0000_0008 ? add_72772 : array_index_72766[8];
  assign array_update_72774[9] = add_72695 == 32'h0000_0009 ? add_72772 : array_index_72766[9];
  assign add_72775 = add_72762 + 32'h0000_0001;
  assign array_update_72776[0] = literal_72009 == 32'h0000_0000 ? array_update_72774 : array_update_72763[0];
  assign array_update_72776[1] = literal_72009 == 32'h0000_0001 ? array_update_72774 : array_update_72763[1];
  assign array_update_72776[2] = literal_72009 == 32'h0000_0002 ? array_update_72774 : array_update_72763[2];
  assign array_update_72776[3] = literal_72009 == 32'h0000_0003 ? array_update_72774 : array_update_72763[3];
  assign array_update_72776[4] = literal_72009 == 32'h0000_0004 ? array_update_72774 : array_update_72763[4];
  assign array_update_72776[5] = literal_72009 == 32'h0000_0005 ? array_update_72774 : array_update_72763[5];
  assign array_update_72776[6] = literal_72009 == 32'h0000_0006 ? array_update_72774 : array_update_72763[6];
  assign array_update_72776[7] = literal_72009 == 32'h0000_0007 ? array_update_72774 : array_update_72763[7];
  assign array_update_72776[8] = literal_72009 == 32'h0000_0008 ? array_update_72774 : array_update_72763[8];
  assign array_update_72776[9] = literal_72009 == 32'h0000_0009 ? array_update_72774 : array_update_72763[9];
  assign array_index_72778 = array_update_72021[add_72775 > 32'h0000_0009 ? 4'h9 : add_72775[3:0]];
  assign array_index_72779 = array_update_72776[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_72783 = smul32b_32b_x_32b(array_index_72024[add_72775 > 32'h0000_0009 ? 4'h9 : add_72775[3:0]], array_index_72778[add_72695 > 32'h0000_0009 ? 4'h9 : add_72695[3:0]]);
  assign add_72785 = array_index_72779[add_72695 > 32'h0000_0009 ? 4'h9 : add_72695[3:0]] + smul_72783;
  assign array_update_72787[0] = add_72695 == 32'h0000_0000 ? add_72785 : array_index_72779[0];
  assign array_update_72787[1] = add_72695 == 32'h0000_0001 ? add_72785 : array_index_72779[1];
  assign array_update_72787[2] = add_72695 == 32'h0000_0002 ? add_72785 : array_index_72779[2];
  assign array_update_72787[3] = add_72695 == 32'h0000_0003 ? add_72785 : array_index_72779[3];
  assign array_update_72787[4] = add_72695 == 32'h0000_0004 ? add_72785 : array_index_72779[4];
  assign array_update_72787[5] = add_72695 == 32'h0000_0005 ? add_72785 : array_index_72779[5];
  assign array_update_72787[6] = add_72695 == 32'h0000_0006 ? add_72785 : array_index_72779[6];
  assign array_update_72787[7] = add_72695 == 32'h0000_0007 ? add_72785 : array_index_72779[7];
  assign array_update_72787[8] = add_72695 == 32'h0000_0008 ? add_72785 : array_index_72779[8];
  assign array_update_72787[9] = add_72695 == 32'h0000_0009 ? add_72785 : array_index_72779[9];
  assign add_72788 = add_72775 + 32'h0000_0001;
  assign array_update_72789[0] = literal_72009 == 32'h0000_0000 ? array_update_72787 : array_update_72776[0];
  assign array_update_72789[1] = literal_72009 == 32'h0000_0001 ? array_update_72787 : array_update_72776[1];
  assign array_update_72789[2] = literal_72009 == 32'h0000_0002 ? array_update_72787 : array_update_72776[2];
  assign array_update_72789[3] = literal_72009 == 32'h0000_0003 ? array_update_72787 : array_update_72776[3];
  assign array_update_72789[4] = literal_72009 == 32'h0000_0004 ? array_update_72787 : array_update_72776[4];
  assign array_update_72789[5] = literal_72009 == 32'h0000_0005 ? array_update_72787 : array_update_72776[5];
  assign array_update_72789[6] = literal_72009 == 32'h0000_0006 ? array_update_72787 : array_update_72776[6];
  assign array_update_72789[7] = literal_72009 == 32'h0000_0007 ? array_update_72787 : array_update_72776[7];
  assign array_update_72789[8] = literal_72009 == 32'h0000_0008 ? array_update_72787 : array_update_72776[8];
  assign array_update_72789[9] = literal_72009 == 32'h0000_0009 ? array_update_72787 : array_update_72776[9];
  assign array_index_72791 = array_update_72021[add_72788 > 32'h0000_0009 ? 4'h9 : add_72788[3:0]];
  assign array_index_72792 = array_update_72789[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_72796 = smul32b_32b_x_32b(array_index_72024[add_72788 > 32'h0000_0009 ? 4'h9 : add_72788[3:0]], array_index_72791[add_72695 > 32'h0000_0009 ? 4'h9 : add_72695[3:0]]);
  assign add_72798 = array_index_72792[add_72695 > 32'h0000_0009 ? 4'h9 : add_72695[3:0]] + smul_72796;
  assign array_update_72800[0] = add_72695 == 32'h0000_0000 ? add_72798 : array_index_72792[0];
  assign array_update_72800[1] = add_72695 == 32'h0000_0001 ? add_72798 : array_index_72792[1];
  assign array_update_72800[2] = add_72695 == 32'h0000_0002 ? add_72798 : array_index_72792[2];
  assign array_update_72800[3] = add_72695 == 32'h0000_0003 ? add_72798 : array_index_72792[3];
  assign array_update_72800[4] = add_72695 == 32'h0000_0004 ? add_72798 : array_index_72792[4];
  assign array_update_72800[5] = add_72695 == 32'h0000_0005 ? add_72798 : array_index_72792[5];
  assign array_update_72800[6] = add_72695 == 32'h0000_0006 ? add_72798 : array_index_72792[6];
  assign array_update_72800[7] = add_72695 == 32'h0000_0007 ? add_72798 : array_index_72792[7];
  assign array_update_72800[8] = add_72695 == 32'h0000_0008 ? add_72798 : array_index_72792[8];
  assign array_update_72800[9] = add_72695 == 32'h0000_0009 ? add_72798 : array_index_72792[9];
  assign add_72801 = add_72788 + 32'h0000_0001;
  assign array_update_72802[0] = literal_72009 == 32'h0000_0000 ? array_update_72800 : array_update_72789[0];
  assign array_update_72802[1] = literal_72009 == 32'h0000_0001 ? array_update_72800 : array_update_72789[1];
  assign array_update_72802[2] = literal_72009 == 32'h0000_0002 ? array_update_72800 : array_update_72789[2];
  assign array_update_72802[3] = literal_72009 == 32'h0000_0003 ? array_update_72800 : array_update_72789[3];
  assign array_update_72802[4] = literal_72009 == 32'h0000_0004 ? array_update_72800 : array_update_72789[4];
  assign array_update_72802[5] = literal_72009 == 32'h0000_0005 ? array_update_72800 : array_update_72789[5];
  assign array_update_72802[6] = literal_72009 == 32'h0000_0006 ? array_update_72800 : array_update_72789[6];
  assign array_update_72802[7] = literal_72009 == 32'h0000_0007 ? array_update_72800 : array_update_72789[7];
  assign array_update_72802[8] = literal_72009 == 32'h0000_0008 ? array_update_72800 : array_update_72789[8];
  assign array_update_72802[9] = literal_72009 == 32'h0000_0009 ? array_update_72800 : array_update_72789[9];
  assign array_index_72804 = array_update_72021[add_72801 > 32'h0000_0009 ? 4'h9 : add_72801[3:0]];
  assign array_index_72805 = array_update_72802[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_72809 = smul32b_32b_x_32b(array_index_72024[add_72801 > 32'h0000_0009 ? 4'h9 : add_72801[3:0]], array_index_72804[add_72695 > 32'h0000_0009 ? 4'h9 : add_72695[3:0]]);
  assign add_72811 = array_index_72805[add_72695 > 32'h0000_0009 ? 4'h9 : add_72695[3:0]] + smul_72809;
  assign array_update_72813[0] = add_72695 == 32'h0000_0000 ? add_72811 : array_index_72805[0];
  assign array_update_72813[1] = add_72695 == 32'h0000_0001 ? add_72811 : array_index_72805[1];
  assign array_update_72813[2] = add_72695 == 32'h0000_0002 ? add_72811 : array_index_72805[2];
  assign array_update_72813[3] = add_72695 == 32'h0000_0003 ? add_72811 : array_index_72805[3];
  assign array_update_72813[4] = add_72695 == 32'h0000_0004 ? add_72811 : array_index_72805[4];
  assign array_update_72813[5] = add_72695 == 32'h0000_0005 ? add_72811 : array_index_72805[5];
  assign array_update_72813[6] = add_72695 == 32'h0000_0006 ? add_72811 : array_index_72805[6];
  assign array_update_72813[7] = add_72695 == 32'h0000_0007 ? add_72811 : array_index_72805[7];
  assign array_update_72813[8] = add_72695 == 32'h0000_0008 ? add_72811 : array_index_72805[8];
  assign array_update_72813[9] = add_72695 == 32'h0000_0009 ? add_72811 : array_index_72805[9];
  assign add_72814 = add_72801 + 32'h0000_0001;
  assign array_update_72815[0] = literal_72009 == 32'h0000_0000 ? array_update_72813 : array_update_72802[0];
  assign array_update_72815[1] = literal_72009 == 32'h0000_0001 ? array_update_72813 : array_update_72802[1];
  assign array_update_72815[2] = literal_72009 == 32'h0000_0002 ? array_update_72813 : array_update_72802[2];
  assign array_update_72815[3] = literal_72009 == 32'h0000_0003 ? array_update_72813 : array_update_72802[3];
  assign array_update_72815[4] = literal_72009 == 32'h0000_0004 ? array_update_72813 : array_update_72802[4];
  assign array_update_72815[5] = literal_72009 == 32'h0000_0005 ? array_update_72813 : array_update_72802[5];
  assign array_update_72815[6] = literal_72009 == 32'h0000_0006 ? array_update_72813 : array_update_72802[6];
  assign array_update_72815[7] = literal_72009 == 32'h0000_0007 ? array_update_72813 : array_update_72802[7];
  assign array_update_72815[8] = literal_72009 == 32'h0000_0008 ? array_update_72813 : array_update_72802[8];
  assign array_update_72815[9] = literal_72009 == 32'h0000_0009 ? array_update_72813 : array_update_72802[9];
  assign array_index_72817 = array_update_72021[add_72814 > 32'h0000_0009 ? 4'h9 : add_72814[3:0]];
  assign array_index_72818 = array_update_72815[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_72822 = smul32b_32b_x_32b(array_index_72024[add_72814 > 32'h0000_0009 ? 4'h9 : add_72814[3:0]], array_index_72817[add_72695 > 32'h0000_0009 ? 4'h9 : add_72695[3:0]]);
  assign add_72824 = array_index_72818[add_72695 > 32'h0000_0009 ? 4'h9 : add_72695[3:0]] + smul_72822;
  assign array_update_72825[0] = add_72695 == 32'h0000_0000 ? add_72824 : array_index_72818[0];
  assign array_update_72825[1] = add_72695 == 32'h0000_0001 ? add_72824 : array_index_72818[1];
  assign array_update_72825[2] = add_72695 == 32'h0000_0002 ? add_72824 : array_index_72818[2];
  assign array_update_72825[3] = add_72695 == 32'h0000_0003 ? add_72824 : array_index_72818[3];
  assign array_update_72825[4] = add_72695 == 32'h0000_0004 ? add_72824 : array_index_72818[4];
  assign array_update_72825[5] = add_72695 == 32'h0000_0005 ? add_72824 : array_index_72818[5];
  assign array_update_72825[6] = add_72695 == 32'h0000_0006 ? add_72824 : array_index_72818[6];
  assign array_update_72825[7] = add_72695 == 32'h0000_0007 ? add_72824 : array_index_72818[7];
  assign array_update_72825[8] = add_72695 == 32'h0000_0008 ? add_72824 : array_index_72818[8];
  assign array_update_72825[9] = add_72695 == 32'h0000_0009 ? add_72824 : array_index_72818[9];
  assign array_update_72826[0] = literal_72009 == 32'h0000_0000 ? array_update_72825 : array_update_72815[0];
  assign array_update_72826[1] = literal_72009 == 32'h0000_0001 ? array_update_72825 : array_update_72815[1];
  assign array_update_72826[2] = literal_72009 == 32'h0000_0002 ? array_update_72825 : array_update_72815[2];
  assign array_update_72826[3] = literal_72009 == 32'h0000_0003 ? array_update_72825 : array_update_72815[3];
  assign array_update_72826[4] = literal_72009 == 32'h0000_0004 ? array_update_72825 : array_update_72815[4];
  assign array_update_72826[5] = literal_72009 == 32'h0000_0005 ? array_update_72825 : array_update_72815[5];
  assign array_update_72826[6] = literal_72009 == 32'h0000_0006 ? array_update_72825 : array_update_72815[6];
  assign array_update_72826[7] = literal_72009 == 32'h0000_0007 ? array_update_72825 : array_update_72815[7];
  assign array_update_72826[8] = literal_72009 == 32'h0000_0008 ? array_update_72825 : array_update_72815[8];
  assign array_update_72826[9] = literal_72009 == 32'h0000_0009 ? array_update_72825 : array_update_72815[9];
  assign array_index_72828 = array_update_72826[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign add_72830 = add_72695 + 32'h0000_0001;
  assign array_update_72831[0] = add_72830 == 32'h0000_0000 ? 32'h0000_0000 : array_index_72828[0];
  assign array_update_72831[1] = add_72830 == 32'h0000_0001 ? 32'h0000_0000 : array_index_72828[1];
  assign array_update_72831[2] = add_72830 == 32'h0000_0002 ? 32'h0000_0000 : array_index_72828[2];
  assign array_update_72831[3] = add_72830 == 32'h0000_0003 ? 32'h0000_0000 : array_index_72828[3];
  assign array_update_72831[4] = add_72830 == 32'h0000_0004 ? 32'h0000_0000 : array_index_72828[4];
  assign array_update_72831[5] = add_72830 == 32'h0000_0005 ? 32'h0000_0000 : array_index_72828[5];
  assign array_update_72831[6] = add_72830 == 32'h0000_0006 ? 32'h0000_0000 : array_index_72828[6];
  assign array_update_72831[7] = add_72830 == 32'h0000_0007 ? 32'h0000_0000 : array_index_72828[7];
  assign array_update_72831[8] = add_72830 == 32'h0000_0008 ? 32'h0000_0000 : array_index_72828[8];
  assign array_update_72831[9] = add_72830 == 32'h0000_0009 ? 32'h0000_0000 : array_index_72828[9];
  assign literal_72832 = 32'h0000_0000;
  assign array_update_72833[0] = literal_72009 == 32'h0000_0000 ? array_update_72831 : array_update_72826[0];
  assign array_update_72833[1] = literal_72009 == 32'h0000_0001 ? array_update_72831 : array_update_72826[1];
  assign array_update_72833[2] = literal_72009 == 32'h0000_0002 ? array_update_72831 : array_update_72826[2];
  assign array_update_72833[3] = literal_72009 == 32'h0000_0003 ? array_update_72831 : array_update_72826[3];
  assign array_update_72833[4] = literal_72009 == 32'h0000_0004 ? array_update_72831 : array_update_72826[4];
  assign array_update_72833[5] = literal_72009 == 32'h0000_0005 ? array_update_72831 : array_update_72826[5];
  assign array_update_72833[6] = literal_72009 == 32'h0000_0006 ? array_update_72831 : array_update_72826[6];
  assign array_update_72833[7] = literal_72009 == 32'h0000_0007 ? array_update_72831 : array_update_72826[7];
  assign array_update_72833[8] = literal_72009 == 32'h0000_0008 ? array_update_72831 : array_update_72826[8];
  assign array_update_72833[9] = literal_72009 == 32'h0000_0009 ? array_update_72831 : array_update_72826[9];
  assign array_index_72835 = array_update_72021[literal_72832 > 32'h0000_0009 ? 4'h9 : literal_72832[3:0]];
  assign array_index_72836 = array_update_72833[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_72840 = smul32b_32b_x_32b(array_index_72024[literal_72832 > 32'h0000_0009 ? 4'h9 : literal_72832[3:0]], array_index_72835[add_72830 > 32'h0000_0009 ? 4'h9 : add_72830[3:0]]);
  assign add_72842 = array_index_72836[add_72830 > 32'h0000_0009 ? 4'h9 : add_72830[3:0]] + smul_72840;
  assign array_update_72844[0] = add_72830 == 32'h0000_0000 ? add_72842 : array_index_72836[0];
  assign array_update_72844[1] = add_72830 == 32'h0000_0001 ? add_72842 : array_index_72836[1];
  assign array_update_72844[2] = add_72830 == 32'h0000_0002 ? add_72842 : array_index_72836[2];
  assign array_update_72844[3] = add_72830 == 32'h0000_0003 ? add_72842 : array_index_72836[3];
  assign array_update_72844[4] = add_72830 == 32'h0000_0004 ? add_72842 : array_index_72836[4];
  assign array_update_72844[5] = add_72830 == 32'h0000_0005 ? add_72842 : array_index_72836[5];
  assign array_update_72844[6] = add_72830 == 32'h0000_0006 ? add_72842 : array_index_72836[6];
  assign array_update_72844[7] = add_72830 == 32'h0000_0007 ? add_72842 : array_index_72836[7];
  assign array_update_72844[8] = add_72830 == 32'h0000_0008 ? add_72842 : array_index_72836[8];
  assign array_update_72844[9] = add_72830 == 32'h0000_0009 ? add_72842 : array_index_72836[9];
  assign add_72845 = literal_72832 + 32'h0000_0001;
  assign array_update_72846[0] = literal_72009 == 32'h0000_0000 ? array_update_72844 : array_update_72833[0];
  assign array_update_72846[1] = literal_72009 == 32'h0000_0001 ? array_update_72844 : array_update_72833[1];
  assign array_update_72846[2] = literal_72009 == 32'h0000_0002 ? array_update_72844 : array_update_72833[2];
  assign array_update_72846[3] = literal_72009 == 32'h0000_0003 ? array_update_72844 : array_update_72833[3];
  assign array_update_72846[4] = literal_72009 == 32'h0000_0004 ? array_update_72844 : array_update_72833[4];
  assign array_update_72846[5] = literal_72009 == 32'h0000_0005 ? array_update_72844 : array_update_72833[5];
  assign array_update_72846[6] = literal_72009 == 32'h0000_0006 ? array_update_72844 : array_update_72833[6];
  assign array_update_72846[7] = literal_72009 == 32'h0000_0007 ? array_update_72844 : array_update_72833[7];
  assign array_update_72846[8] = literal_72009 == 32'h0000_0008 ? array_update_72844 : array_update_72833[8];
  assign array_update_72846[9] = literal_72009 == 32'h0000_0009 ? array_update_72844 : array_update_72833[9];
  assign array_index_72848 = array_update_72021[add_72845 > 32'h0000_0009 ? 4'h9 : add_72845[3:0]];
  assign array_index_72849 = array_update_72846[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_72853 = smul32b_32b_x_32b(array_index_72024[add_72845 > 32'h0000_0009 ? 4'h9 : add_72845[3:0]], array_index_72848[add_72830 > 32'h0000_0009 ? 4'h9 : add_72830[3:0]]);
  assign add_72855 = array_index_72849[add_72830 > 32'h0000_0009 ? 4'h9 : add_72830[3:0]] + smul_72853;
  assign array_update_72857[0] = add_72830 == 32'h0000_0000 ? add_72855 : array_index_72849[0];
  assign array_update_72857[1] = add_72830 == 32'h0000_0001 ? add_72855 : array_index_72849[1];
  assign array_update_72857[2] = add_72830 == 32'h0000_0002 ? add_72855 : array_index_72849[2];
  assign array_update_72857[3] = add_72830 == 32'h0000_0003 ? add_72855 : array_index_72849[3];
  assign array_update_72857[4] = add_72830 == 32'h0000_0004 ? add_72855 : array_index_72849[4];
  assign array_update_72857[5] = add_72830 == 32'h0000_0005 ? add_72855 : array_index_72849[5];
  assign array_update_72857[6] = add_72830 == 32'h0000_0006 ? add_72855 : array_index_72849[6];
  assign array_update_72857[7] = add_72830 == 32'h0000_0007 ? add_72855 : array_index_72849[7];
  assign array_update_72857[8] = add_72830 == 32'h0000_0008 ? add_72855 : array_index_72849[8];
  assign array_update_72857[9] = add_72830 == 32'h0000_0009 ? add_72855 : array_index_72849[9];
  assign add_72858 = add_72845 + 32'h0000_0001;
  assign array_update_72859[0] = literal_72009 == 32'h0000_0000 ? array_update_72857 : array_update_72846[0];
  assign array_update_72859[1] = literal_72009 == 32'h0000_0001 ? array_update_72857 : array_update_72846[1];
  assign array_update_72859[2] = literal_72009 == 32'h0000_0002 ? array_update_72857 : array_update_72846[2];
  assign array_update_72859[3] = literal_72009 == 32'h0000_0003 ? array_update_72857 : array_update_72846[3];
  assign array_update_72859[4] = literal_72009 == 32'h0000_0004 ? array_update_72857 : array_update_72846[4];
  assign array_update_72859[5] = literal_72009 == 32'h0000_0005 ? array_update_72857 : array_update_72846[5];
  assign array_update_72859[6] = literal_72009 == 32'h0000_0006 ? array_update_72857 : array_update_72846[6];
  assign array_update_72859[7] = literal_72009 == 32'h0000_0007 ? array_update_72857 : array_update_72846[7];
  assign array_update_72859[8] = literal_72009 == 32'h0000_0008 ? array_update_72857 : array_update_72846[8];
  assign array_update_72859[9] = literal_72009 == 32'h0000_0009 ? array_update_72857 : array_update_72846[9];
  assign array_index_72861 = array_update_72021[add_72858 > 32'h0000_0009 ? 4'h9 : add_72858[3:0]];
  assign array_index_72862 = array_update_72859[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_72866 = smul32b_32b_x_32b(array_index_72024[add_72858 > 32'h0000_0009 ? 4'h9 : add_72858[3:0]], array_index_72861[add_72830 > 32'h0000_0009 ? 4'h9 : add_72830[3:0]]);
  assign add_72868 = array_index_72862[add_72830 > 32'h0000_0009 ? 4'h9 : add_72830[3:0]] + smul_72866;
  assign array_update_72870[0] = add_72830 == 32'h0000_0000 ? add_72868 : array_index_72862[0];
  assign array_update_72870[1] = add_72830 == 32'h0000_0001 ? add_72868 : array_index_72862[1];
  assign array_update_72870[2] = add_72830 == 32'h0000_0002 ? add_72868 : array_index_72862[2];
  assign array_update_72870[3] = add_72830 == 32'h0000_0003 ? add_72868 : array_index_72862[3];
  assign array_update_72870[4] = add_72830 == 32'h0000_0004 ? add_72868 : array_index_72862[4];
  assign array_update_72870[5] = add_72830 == 32'h0000_0005 ? add_72868 : array_index_72862[5];
  assign array_update_72870[6] = add_72830 == 32'h0000_0006 ? add_72868 : array_index_72862[6];
  assign array_update_72870[7] = add_72830 == 32'h0000_0007 ? add_72868 : array_index_72862[7];
  assign array_update_72870[8] = add_72830 == 32'h0000_0008 ? add_72868 : array_index_72862[8];
  assign array_update_72870[9] = add_72830 == 32'h0000_0009 ? add_72868 : array_index_72862[9];
  assign add_72871 = add_72858 + 32'h0000_0001;
  assign array_update_72872[0] = literal_72009 == 32'h0000_0000 ? array_update_72870 : array_update_72859[0];
  assign array_update_72872[1] = literal_72009 == 32'h0000_0001 ? array_update_72870 : array_update_72859[1];
  assign array_update_72872[2] = literal_72009 == 32'h0000_0002 ? array_update_72870 : array_update_72859[2];
  assign array_update_72872[3] = literal_72009 == 32'h0000_0003 ? array_update_72870 : array_update_72859[3];
  assign array_update_72872[4] = literal_72009 == 32'h0000_0004 ? array_update_72870 : array_update_72859[4];
  assign array_update_72872[5] = literal_72009 == 32'h0000_0005 ? array_update_72870 : array_update_72859[5];
  assign array_update_72872[6] = literal_72009 == 32'h0000_0006 ? array_update_72870 : array_update_72859[6];
  assign array_update_72872[7] = literal_72009 == 32'h0000_0007 ? array_update_72870 : array_update_72859[7];
  assign array_update_72872[8] = literal_72009 == 32'h0000_0008 ? array_update_72870 : array_update_72859[8];
  assign array_update_72872[9] = literal_72009 == 32'h0000_0009 ? array_update_72870 : array_update_72859[9];
  assign array_index_72874 = array_update_72021[add_72871 > 32'h0000_0009 ? 4'h9 : add_72871[3:0]];
  assign array_index_72875 = array_update_72872[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_72879 = smul32b_32b_x_32b(array_index_72024[add_72871 > 32'h0000_0009 ? 4'h9 : add_72871[3:0]], array_index_72874[add_72830 > 32'h0000_0009 ? 4'h9 : add_72830[3:0]]);
  assign add_72881 = array_index_72875[add_72830 > 32'h0000_0009 ? 4'h9 : add_72830[3:0]] + smul_72879;
  assign array_update_72883[0] = add_72830 == 32'h0000_0000 ? add_72881 : array_index_72875[0];
  assign array_update_72883[1] = add_72830 == 32'h0000_0001 ? add_72881 : array_index_72875[1];
  assign array_update_72883[2] = add_72830 == 32'h0000_0002 ? add_72881 : array_index_72875[2];
  assign array_update_72883[3] = add_72830 == 32'h0000_0003 ? add_72881 : array_index_72875[3];
  assign array_update_72883[4] = add_72830 == 32'h0000_0004 ? add_72881 : array_index_72875[4];
  assign array_update_72883[5] = add_72830 == 32'h0000_0005 ? add_72881 : array_index_72875[5];
  assign array_update_72883[6] = add_72830 == 32'h0000_0006 ? add_72881 : array_index_72875[6];
  assign array_update_72883[7] = add_72830 == 32'h0000_0007 ? add_72881 : array_index_72875[7];
  assign array_update_72883[8] = add_72830 == 32'h0000_0008 ? add_72881 : array_index_72875[8];
  assign array_update_72883[9] = add_72830 == 32'h0000_0009 ? add_72881 : array_index_72875[9];
  assign add_72884 = add_72871 + 32'h0000_0001;
  assign array_update_72885[0] = literal_72009 == 32'h0000_0000 ? array_update_72883 : array_update_72872[0];
  assign array_update_72885[1] = literal_72009 == 32'h0000_0001 ? array_update_72883 : array_update_72872[1];
  assign array_update_72885[2] = literal_72009 == 32'h0000_0002 ? array_update_72883 : array_update_72872[2];
  assign array_update_72885[3] = literal_72009 == 32'h0000_0003 ? array_update_72883 : array_update_72872[3];
  assign array_update_72885[4] = literal_72009 == 32'h0000_0004 ? array_update_72883 : array_update_72872[4];
  assign array_update_72885[5] = literal_72009 == 32'h0000_0005 ? array_update_72883 : array_update_72872[5];
  assign array_update_72885[6] = literal_72009 == 32'h0000_0006 ? array_update_72883 : array_update_72872[6];
  assign array_update_72885[7] = literal_72009 == 32'h0000_0007 ? array_update_72883 : array_update_72872[7];
  assign array_update_72885[8] = literal_72009 == 32'h0000_0008 ? array_update_72883 : array_update_72872[8];
  assign array_update_72885[9] = literal_72009 == 32'h0000_0009 ? array_update_72883 : array_update_72872[9];
  assign array_index_72887 = array_update_72021[add_72884 > 32'h0000_0009 ? 4'h9 : add_72884[3:0]];
  assign array_index_72888 = array_update_72885[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_72892 = smul32b_32b_x_32b(array_index_72024[add_72884 > 32'h0000_0009 ? 4'h9 : add_72884[3:0]], array_index_72887[add_72830 > 32'h0000_0009 ? 4'h9 : add_72830[3:0]]);
  assign add_72894 = array_index_72888[add_72830 > 32'h0000_0009 ? 4'h9 : add_72830[3:0]] + smul_72892;
  assign array_update_72896[0] = add_72830 == 32'h0000_0000 ? add_72894 : array_index_72888[0];
  assign array_update_72896[1] = add_72830 == 32'h0000_0001 ? add_72894 : array_index_72888[1];
  assign array_update_72896[2] = add_72830 == 32'h0000_0002 ? add_72894 : array_index_72888[2];
  assign array_update_72896[3] = add_72830 == 32'h0000_0003 ? add_72894 : array_index_72888[3];
  assign array_update_72896[4] = add_72830 == 32'h0000_0004 ? add_72894 : array_index_72888[4];
  assign array_update_72896[5] = add_72830 == 32'h0000_0005 ? add_72894 : array_index_72888[5];
  assign array_update_72896[6] = add_72830 == 32'h0000_0006 ? add_72894 : array_index_72888[6];
  assign array_update_72896[7] = add_72830 == 32'h0000_0007 ? add_72894 : array_index_72888[7];
  assign array_update_72896[8] = add_72830 == 32'h0000_0008 ? add_72894 : array_index_72888[8];
  assign array_update_72896[9] = add_72830 == 32'h0000_0009 ? add_72894 : array_index_72888[9];
  assign add_72897 = add_72884 + 32'h0000_0001;
  assign array_update_72898[0] = literal_72009 == 32'h0000_0000 ? array_update_72896 : array_update_72885[0];
  assign array_update_72898[1] = literal_72009 == 32'h0000_0001 ? array_update_72896 : array_update_72885[1];
  assign array_update_72898[2] = literal_72009 == 32'h0000_0002 ? array_update_72896 : array_update_72885[2];
  assign array_update_72898[3] = literal_72009 == 32'h0000_0003 ? array_update_72896 : array_update_72885[3];
  assign array_update_72898[4] = literal_72009 == 32'h0000_0004 ? array_update_72896 : array_update_72885[4];
  assign array_update_72898[5] = literal_72009 == 32'h0000_0005 ? array_update_72896 : array_update_72885[5];
  assign array_update_72898[6] = literal_72009 == 32'h0000_0006 ? array_update_72896 : array_update_72885[6];
  assign array_update_72898[7] = literal_72009 == 32'h0000_0007 ? array_update_72896 : array_update_72885[7];
  assign array_update_72898[8] = literal_72009 == 32'h0000_0008 ? array_update_72896 : array_update_72885[8];
  assign array_update_72898[9] = literal_72009 == 32'h0000_0009 ? array_update_72896 : array_update_72885[9];
  assign array_index_72900 = array_update_72021[add_72897 > 32'h0000_0009 ? 4'h9 : add_72897[3:0]];
  assign array_index_72901 = array_update_72898[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_72905 = smul32b_32b_x_32b(array_index_72024[add_72897 > 32'h0000_0009 ? 4'h9 : add_72897[3:0]], array_index_72900[add_72830 > 32'h0000_0009 ? 4'h9 : add_72830[3:0]]);
  assign add_72907 = array_index_72901[add_72830 > 32'h0000_0009 ? 4'h9 : add_72830[3:0]] + smul_72905;
  assign array_update_72909[0] = add_72830 == 32'h0000_0000 ? add_72907 : array_index_72901[0];
  assign array_update_72909[1] = add_72830 == 32'h0000_0001 ? add_72907 : array_index_72901[1];
  assign array_update_72909[2] = add_72830 == 32'h0000_0002 ? add_72907 : array_index_72901[2];
  assign array_update_72909[3] = add_72830 == 32'h0000_0003 ? add_72907 : array_index_72901[3];
  assign array_update_72909[4] = add_72830 == 32'h0000_0004 ? add_72907 : array_index_72901[4];
  assign array_update_72909[5] = add_72830 == 32'h0000_0005 ? add_72907 : array_index_72901[5];
  assign array_update_72909[6] = add_72830 == 32'h0000_0006 ? add_72907 : array_index_72901[6];
  assign array_update_72909[7] = add_72830 == 32'h0000_0007 ? add_72907 : array_index_72901[7];
  assign array_update_72909[8] = add_72830 == 32'h0000_0008 ? add_72907 : array_index_72901[8];
  assign array_update_72909[9] = add_72830 == 32'h0000_0009 ? add_72907 : array_index_72901[9];
  assign add_72910 = add_72897 + 32'h0000_0001;
  assign array_update_72911[0] = literal_72009 == 32'h0000_0000 ? array_update_72909 : array_update_72898[0];
  assign array_update_72911[1] = literal_72009 == 32'h0000_0001 ? array_update_72909 : array_update_72898[1];
  assign array_update_72911[2] = literal_72009 == 32'h0000_0002 ? array_update_72909 : array_update_72898[2];
  assign array_update_72911[3] = literal_72009 == 32'h0000_0003 ? array_update_72909 : array_update_72898[3];
  assign array_update_72911[4] = literal_72009 == 32'h0000_0004 ? array_update_72909 : array_update_72898[4];
  assign array_update_72911[5] = literal_72009 == 32'h0000_0005 ? array_update_72909 : array_update_72898[5];
  assign array_update_72911[6] = literal_72009 == 32'h0000_0006 ? array_update_72909 : array_update_72898[6];
  assign array_update_72911[7] = literal_72009 == 32'h0000_0007 ? array_update_72909 : array_update_72898[7];
  assign array_update_72911[8] = literal_72009 == 32'h0000_0008 ? array_update_72909 : array_update_72898[8];
  assign array_update_72911[9] = literal_72009 == 32'h0000_0009 ? array_update_72909 : array_update_72898[9];
  assign array_index_72913 = array_update_72021[add_72910 > 32'h0000_0009 ? 4'h9 : add_72910[3:0]];
  assign array_index_72914 = array_update_72911[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_72918 = smul32b_32b_x_32b(array_index_72024[add_72910 > 32'h0000_0009 ? 4'h9 : add_72910[3:0]], array_index_72913[add_72830 > 32'h0000_0009 ? 4'h9 : add_72830[3:0]]);
  assign add_72920 = array_index_72914[add_72830 > 32'h0000_0009 ? 4'h9 : add_72830[3:0]] + smul_72918;
  assign array_update_72922[0] = add_72830 == 32'h0000_0000 ? add_72920 : array_index_72914[0];
  assign array_update_72922[1] = add_72830 == 32'h0000_0001 ? add_72920 : array_index_72914[1];
  assign array_update_72922[2] = add_72830 == 32'h0000_0002 ? add_72920 : array_index_72914[2];
  assign array_update_72922[3] = add_72830 == 32'h0000_0003 ? add_72920 : array_index_72914[3];
  assign array_update_72922[4] = add_72830 == 32'h0000_0004 ? add_72920 : array_index_72914[4];
  assign array_update_72922[5] = add_72830 == 32'h0000_0005 ? add_72920 : array_index_72914[5];
  assign array_update_72922[6] = add_72830 == 32'h0000_0006 ? add_72920 : array_index_72914[6];
  assign array_update_72922[7] = add_72830 == 32'h0000_0007 ? add_72920 : array_index_72914[7];
  assign array_update_72922[8] = add_72830 == 32'h0000_0008 ? add_72920 : array_index_72914[8];
  assign array_update_72922[9] = add_72830 == 32'h0000_0009 ? add_72920 : array_index_72914[9];
  assign add_72923 = add_72910 + 32'h0000_0001;
  assign array_update_72924[0] = literal_72009 == 32'h0000_0000 ? array_update_72922 : array_update_72911[0];
  assign array_update_72924[1] = literal_72009 == 32'h0000_0001 ? array_update_72922 : array_update_72911[1];
  assign array_update_72924[2] = literal_72009 == 32'h0000_0002 ? array_update_72922 : array_update_72911[2];
  assign array_update_72924[3] = literal_72009 == 32'h0000_0003 ? array_update_72922 : array_update_72911[3];
  assign array_update_72924[4] = literal_72009 == 32'h0000_0004 ? array_update_72922 : array_update_72911[4];
  assign array_update_72924[5] = literal_72009 == 32'h0000_0005 ? array_update_72922 : array_update_72911[5];
  assign array_update_72924[6] = literal_72009 == 32'h0000_0006 ? array_update_72922 : array_update_72911[6];
  assign array_update_72924[7] = literal_72009 == 32'h0000_0007 ? array_update_72922 : array_update_72911[7];
  assign array_update_72924[8] = literal_72009 == 32'h0000_0008 ? array_update_72922 : array_update_72911[8];
  assign array_update_72924[9] = literal_72009 == 32'h0000_0009 ? array_update_72922 : array_update_72911[9];
  assign array_index_72926 = array_update_72021[add_72923 > 32'h0000_0009 ? 4'h9 : add_72923[3:0]];
  assign array_index_72927 = array_update_72924[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_72931 = smul32b_32b_x_32b(array_index_72024[add_72923 > 32'h0000_0009 ? 4'h9 : add_72923[3:0]], array_index_72926[add_72830 > 32'h0000_0009 ? 4'h9 : add_72830[3:0]]);
  assign add_72933 = array_index_72927[add_72830 > 32'h0000_0009 ? 4'h9 : add_72830[3:0]] + smul_72931;
  assign array_update_72935[0] = add_72830 == 32'h0000_0000 ? add_72933 : array_index_72927[0];
  assign array_update_72935[1] = add_72830 == 32'h0000_0001 ? add_72933 : array_index_72927[1];
  assign array_update_72935[2] = add_72830 == 32'h0000_0002 ? add_72933 : array_index_72927[2];
  assign array_update_72935[3] = add_72830 == 32'h0000_0003 ? add_72933 : array_index_72927[3];
  assign array_update_72935[4] = add_72830 == 32'h0000_0004 ? add_72933 : array_index_72927[4];
  assign array_update_72935[5] = add_72830 == 32'h0000_0005 ? add_72933 : array_index_72927[5];
  assign array_update_72935[6] = add_72830 == 32'h0000_0006 ? add_72933 : array_index_72927[6];
  assign array_update_72935[7] = add_72830 == 32'h0000_0007 ? add_72933 : array_index_72927[7];
  assign array_update_72935[8] = add_72830 == 32'h0000_0008 ? add_72933 : array_index_72927[8];
  assign array_update_72935[9] = add_72830 == 32'h0000_0009 ? add_72933 : array_index_72927[9];
  assign add_72936 = add_72923 + 32'h0000_0001;
  assign array_update_72937[0] = literal_72009 == 32'h0000_0000 ? array_update_72935 : array_update_72924[0];
  assign array_update_72937[1] = literal_72009 == 32'h0000_0001 ? array_update_72935 : array_update_72924[1];
  assign array_update_72937[2] = literal_72009 == 32'h0000_0002 ? array_update_72935 : array_update_72924[2];
  assign array_update_72937[3] = literal_72009 == 32'h0000_0003 ? array_update_72935 : array_update_72924[3];
  assign array_update_72937[4] = literal_72009 == 32'h0000_0004 ? array_update_72935 : array_update_72924[4];
  assign array_update_72937[5] = literal_72009 == 32'h0000_0005 ? array_update_72935 : array_update_72924[5];
  assign array_update_72937[6] = literal_72009 == 32'h0000_0006 ? array_update_72935 : array_update_72924[6];
  assign array_update_72937[7] = literal_72009 == 32'h0000_0007 ? array_update_72935 : array_update_72924[7];
  assign array_update_72937[8] = literal_72009 == 32'h0000_0008 ? array_update_72935 : array_update_72924[8];
  assign array_update_72937[9] = literal_72009 == 32'h0000_0009 ? array_update_72935 : array_update_72924[9];
  assign array_index_72939 = array_update_72021[add_72936 > 32'h0000_0009 ? 4'h9 : add_72936[3:0]];
  assign array_index_72940 = array_update_72937[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_72944 = smul32b_32b_x_32b(array_index_72024[add_72936 > 32'h0000_0009 ? 4'h9 : add_72936[3:0]], array_index_72939[add_72830 > 32'h0000_0009 ? 4'h9 : add_72830[3:0]]);
  assign add_72946 = array_index_72940[add_72830 > 32'h0000_0009 ? 4'h9 : add_72830[3:0]] + smul_72944;
  assign array_update_72948[0] = add_72830 == 32'h0000_0000 ? add_72946 : array_index_72940[0];
  assign array_update_72948[1] = add_72830 == 32'h0000_0001 ? add_72946 : array_index_72940[1];
  assign array_update_72948[2] = add_72830 == 32'h0000_0002 ? add_72946 : array_index_72940[2];
  assign array_update_72948[3] = add_72830 == 32'h0000_0003 ? add_72946 : array_index_72940[3];
  assign array_update_72948[4] = add_72830 == 32'h0000_0004 ? add_72946 : array_index_72940[4];
  assign array_update_72948[5] = add_72830 == 32'h0000_0005 ? add_72946 : array_index_72940[5];
  assign array_update_72948[6] = add_72830 == 32'h0000_0006 ? add_72946 : array_index_72940[6];
  assign array_update_72948[7] = add_72830 == 32'h0000_0007 ? add_72946 : array_index_72940[7];
  assign array_update_72948[8] = add_72830 == 32'h0000_0008 ? add_72946 : array_index_72940[8];
  assign array_update_72948[9] = add_72830 == 32'h0000_0009 ? add_72946 : array_index_72940[9];
  assign add_72949 = add_72936 + 32'h0000_0001;
  assign array_update_72950[0] = literal_72009 == 32'h0000_0000 ? array_update_72948 : array_update_72937[0];
  assign array_update_72950[1] = literal_72009 == 32'h0000_0001 ? array_update_72948 : array_update_72937[1];
  assign array_update_72950[2] = literal_72009 == 32'h0000_0002 ? array_update_72948 : array_update_72937[2];
  assign array_update_72950[3] = literal_72009 == 32'h0000_0003 ? array_update_72948 : array_update_72937[3];
  assign array_update_72950[4] = literal_72009 == 32'h0000_0004 ? array_update_72948 : array_update_72937[4];
  assign array_update_72950[5] = literal_72009 == 32'h0000_0005 ? array_update_72948 : array_update_72937[5];
  assign array_update_72950[6] = literal_72009 == 32'h0000_0006 ? array_update_72948 : array_update_72937[6];
  assign array_update_72950[7] = literal_72009 == 32'h0000_0007 ? array_update_72948 : array_update_72937[7];
  assign array_update_72950[8] = literal_72009 == 32'h0000_0008 ? array_update_72948 : array_update_72937[8];
  assign array_update_72950[9] = literal_72009 == 32'h0000_0009 ? array_update_72948 : array_update_72937[9];
  assign array_index_72952 = array_update_72021[add_72949 > 32'h0000_0009 ? 4'h9 : add_72949[3:0]];
  assign array_index_72953 = array_update_72950[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_72957 = smul32b_32b_x_32b(array_index_72024[add_72949 > 32'h0000_0009 ? 4'h9 : add_72949[3:0]], array_index_72952[add_72830 > 32'h0000_0009 ? 4'h9 : add_72830[3:0]]);
  assign add_72959 = array_index_72953[add_72830 > 32'h0000_0009 ? 4'h9 : add_72830[3:0]] + smul_72957;
  assign array_update_72960[0] = add_72830 == 32'h0000_0000 ? add_72959 : array_index_72953[0];
  assign array_update_72960[1] = add_72830 == 32'h0000_0001 ? add_72959 : array_index_72953[1];
  assign array_update_72960[2] = add_72830 == 32'h0000_0002 ? add_72959 : array_index_72953[2];
  assign array_update_72960[3] = add_72830 == 32'h0000_0003 ? add_72959 : array_index_72953[3];
  assign array_update_72960[4] = add_72830 == 32'h0000_0004 ? add_72959 : array_index_72953[4];
  assign array_update_72960[5] = add_72830 == 32'h0000_0005 ? add_72959 : array_index_72953[5];
  assign array_update_72960[6] = add_72830 == 32'h0000_0006 ? add_72959 : array_index_72953[6];
  assign array_update_72960[7] = add_72830 == 32'h0000_0007 ? add_72959 : array_index_72953[7];
  assign array_update_72960[8] = add_72830 == 32'h0000_0008 ? add_72959 : array_index_72953[8];
  assign array_update_72960[9] = add_72830 == 32'h0000_0009 ? add_72959 : array_index_72953[9];
  assign array_update_72961[0] = literal_72009 == 32'h0000_0000 ? array_update_72960 : array_update_72950[0];
  assign array_update_72961[1] = literal_72009 == 32'h0000_0001 ? array_update_72960 : array_update_72950[1];
  assign array_update_72961[2] = literal_72009 == 32'h0000_0002 ? array_update_72960 : array_update_72950[2];
  assign array_update_72961[3] = literal_72009 == 32'h0000_0003 ? array_update_72960 : array_update_72950[3];
  assign array_update_72961[4] = literal_72009 == 32'h0000_0004 ? array_update_72960 : array_update_72950[4];
  assign array_update_72961[5] = literal_72009 == 32'h0000_0005 ? array_update_72960 : array_update_72950[5];
  assign array_update_72961[6] = literal_72009 == 32'h0000_0006 ? array_update_72960 : array_update_72950[6];
  assign array_update_72961[7] = literal_72009 == 32'h0000_0007 ? array_update_72960 : array_update_72950[7];
  assign array_update_72961[8] = literal_72009 == 32'h0000_0008 ? array_update_72960 : array_update_72950[8];
  assign array_update_72961[9] = literal_72009 == 32'h0000_0009 ? array_update_72960 : array_update_72950[9];
  assign array_index_72963 = array_update_72961[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign add_72965 = add_72830 + 32'h0000_0001;
  assign array_update_72966[0] = add_72965 == 32'h0000_0000 ? 32'h0000_0000 : array_index_72963[0];
  assign array_update_72966[1] = add_72965 == 32'h0000_0001 ? 32'h0000_0000 : array_index_72963[1];
  assign array_update_72966[2] = add_72965 == 32'h0000_0002 ? 32'h0000_0000 : array_index_72963[2];
  assign array_update_72966[3] = add_72965 == 32'h0000_0003 ? 32'h0000_0000 : array_index_72963[3];
  assign array_update_72966[4] = add_72965 == 32'h0000_0004 ? 32'h0000_0000 : array_index_72963[4];
  assign array_update_72966[5] = add_72965 == 32'h0000_0005 ? 32'h0000_0000 : array_index_72963[5];
  assign array_update_72966[6] = add_72965 == 32'h0000_0006 ? 32'h0000_0000 : array_index_72963[6];
  assign array_update_72966[7] = add_72965 == 32'h0000_0007 ? 32'h0000_0000 : array_index_72963[7];
  assign array_update_72966[8] = add_72965 == 32'h0000_0008 ? 32'h0000_0000 : array_index_72963[8];
  assign array_update_72966[9] = add_72965 == 32'h0000_0009 ? 32'h0000_0000 : array_index_72963[9];
  assign literal_72967 = 32'h0000_0000;
  assign array_update_72968[0] = literal_72009 == 32'h0000_0000 ? array_update_72966 : array_update_72961[0];
  assign array_update_72968[1] = literal_72009 == 32'h0000_0001 ? array_update_72966 : array_update_72961[1];
  assign array_update_72968[2] = literal_72009 == 32'h0000_0002 ? array_update_72966 : array_update_72961[2];
  assign array_update_72968[3] = literal_72009 == 32'h0000_0003 ? array_update_72966 : array_update_72961[3];
  assign array_update_72968[4] = literal_72009 == 32'h0000_0004 ? array_update_72966 : array_update_72961[4];
  assign array_update_72968[5] = literal_72009 == 32'h0000_0005 ? array_update_72966 : array_update_72961[5];
  assign array_update_72968[6] = literal_72009 == 32'h0000_0006 ? array_update_72966 : array_update_72961[6];
  assign array_update_72968[7] = literal_72009 == 32'h0000_0007 ? array_update_72966 : array_update_72961[7];
  assign array_update_72968[8] = literal_72009 == 32'h0000_0008 ? array_update_72966 : array_update_72961[8];
  assign array_update_72968[9] = literal_72009 == 32'h0000_0009 ? array_update_72966 : array_update_72961[9];
  assign array_index_72970 = array_update_72021[literal_72967 > 32'h0000_0009 ? 4'h9 : literal_72967[3:0]];
  assign array_index_72971 = array_update_72968[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_72975 = smul32b_32b_x_32b(array_index_72024[literal_72967 > 32'h0000_0009 ? 4'h9 : literal_72967[3:0]], array_index_72970[add_72965 > 32'h0000_0009 ? 4'h9 : add_72965[3:0]]);
  assign add_72977 = array_index_72971[add_72965 > 32'h0000_0009 ? 4'h9 : add_72965[3:0]] + smul_72975;
  assign array_update_72979[0] = add_72965 == 32'h0000_0000 ? add_72977 : array_index_72971[0];
  assign array_update_72979[1] = add_72965 == 32'h0000_0001 ? add_72977 : array_index_72971[1];
  assign array_update_72979[2] = add_72965 == 32'h0000_0002 ? add_72977 : array_index_72971[2];
  assign array_update_72979[3] = add_72965 == 32'h0000_0003 ? add_72977 : array_index_72971[3];
  assign array_update_72979[4] = add_72965 == 32'h0000_0004 ? add_72977 : array_index_72971[4];
  assign array_update_72979[5] = add_72965 == 32'h0000_0005 ? add_72977 : array_index_72971[5];
  assign array_update_72979[6] = add_72965 == 32'h0000_0006 ? add_72977 : array_index_72971[6];
  assign array_update_72979[7] = add_72965 == 32'h0000_0007 ? add_72977 : array_index_72971[7];
  assign array_update_72979[8] = add_72965 == 32'h0000_0008 ? add_72977 : array_index_72971[8];
  assign array_update_72979[9] = add_72965 == 32'h0000_0009 ? add_72977 : array_index_72971[9];
  assign add_72980 = literal_72967 + 32'h0000_0001;
  assign array_update_72981[0] = literal_72009 == 32'h0000_0000 ? array_update_72979 : array_update_72968[0];
  assign array_update_72981[1] = literal_72009 == 32'h0000_0001 ? array_update_72979 : array_update_72968[1];
  assign array_update_72981[2] = literal_72009 == 32'h0000_0002 ? array_update_72979 : array_update_72968[2];
  assign array_update_72981[3] = literal_72009 == 32'h0000_0003 ? array_update_72979 : array_update_72968[3];
  assign array_update_72981[4] = literal_72009 == 32'h0000_0004 ? array_update_72979 : array_update_72968[4];
  assign array_update_72981[5] = literal_72009 == 32'h0000_0005 ? array_update_72979 : array_update_72968[5];
  assign array_update_72981[6] = literal_72009 == 32'h0000_0006 ? array_update_72979 : array_update_72968[6];
  assign array_update_72981[7] = literal_72009 == 32'h0000_0007 ? array_update_72979 : array_update_72968[7];
  assign array_update_72981[8] = literal_72009 == 32'h0000_0008 ? array_update_72979 : array_update_72968[8];
  assign array_update_72981[9] = literal_72009 == 32'h0000_0009 ? array_update_72979 : array_update_72968[9];
  assign array_index_72983 = array_update_72021[add_72980 > 32'h0000_0009 ? 4'h9 : add_72980[3:0]];
  assign array_index_72984 = array_update_72981[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_72988 = smul32b_32b_x_32b(array_index_72024[add_72980 > 32'h0000_0009 ? 4'h9 : add_72980[3:0]], array_index_72983[add_72965 > 32'h0000_0009 ? 4'h9 : add_72965[3:0]]);
  assign add_72990 = array_index_72984[add_72965 > 32'h0000_0009 ? 4'h9 : add_72965[3:0]] + smul_72988;
  assign array_update_72992[0] = add_72965 == 32'h0000_0000 ? add_72990 : array_index_72984[0];
  assign array_update_72992[1] = add_72965 == 32'h0000_0001 ? add_72990 : array_index_72984[1];
  assign array_update_72992[2] = add_72965 == 32'h0000_0002 ? add_72990 : array_index_72984[2];
  assign array_update_72992[3] = add_72965 == 32'h0000_0003 ? add_72990 : array_index_72984[3];
  assign array_update_72992[4] = add_72965 == 32'h0000_0004 ? add_72990 : array_index_72984[4];
  assign array_update_72992[5] = add_72965 == 32'h0000_0005 ? add_72990 : array_index_72984[5];
  assign array_update_72992[6] = add_72965 == 32'h0000_0006 ? add_72990 : array_index_72984[6];
  assign array_update_72992[7] = add_72965 == 32'h0000_0007 ? add_72990 : array_index_72984[7];
  assign array_update_72992[8] = add_72965 == 32'h0000_0008 ? add_72990 : array_index_72984[8];
  assign array_update_72992[9] = add_72965 == 32'h0000_0009 ? add_72990 : array_index_72984[9];
  assign add_72993 = add_72980 + 32'h0000_0001;
  assign array_update_72994[0] = literal_72009 == 32'h0000_0000 ? array_update_72992 : array_update_72981[0];
  assign array_update_72994[1] = literal_72009 == 32'h0000_0001 ? array_update_72992 : array_update_72981[1];
  assign array_update_72994[2] = literal_72009 == 32'h0000_0002 ? array_update_72992 : array_update_72981[2];
  assign array_update_72994[3] = literal_72009 == 32'h0000_0003 ? array_update_72992 : array_update_72981[3];
  assign array_update_72994[4] = literal_72009 == 32'h0000_0004 ? array_update_72992 : array_update_72981[4];
  assign array_update_72994[5] = literal_72009 == 32'h0000_0005 ? array_update_72992 : array_update_72981[5];
  assign array_update_72994[6] = literal_72009 == 32'h0000_0006 ? array_update_72992 : array_update_72981[6];
  assign array_update_72994[7] = literal_72009 == 32'h0000_0007 ? array_update_72992 : array_update_72981[7];
  assign array_update_72994[8] = literal_72009 == 32'h0000_0008 ? array_update_72992 : array_update_72981[8];
  assign array_update_72994[9] = literal_72009 == 32'h0000_0009 ? array_update_72992 : array_update_72981[9];
  assign array_index_72996 = array_update_72021[add_72993 > 32'h0000_0009 ? 4'h9 : add_72993[3:0]];
  assign array_index_72997 = array_update_72994[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_73001 = smul32b_32b_x_32b(array_index_72024[add_72993 > 32'h0000_0009 ? 4'h9 : add_72993[3:0]], array_index_72996[add_72965 > 32'h0000_0009 ? 4'h9 : add_72965[3:0]]);
  assign add_73003 = array_index_72997[add_72965 > 32'h0000_0009 ? 4'h9 : add_72965[3:0]] + smul_73001;
  assign array_update_73005[0] = add_72965 == 32'h0000_0000 ? add_73003 : array_index_72997[0];
  assign array_update_73005[1] = add_72965 == 32'h0000_0001 ? add_73003 : array_index_72997[1];
  assign array_update_73005[2] = add_72965 == 32'h0000_0002 ? add_73003 : array_index_72997[2];
  assign array_update_73005[3] = add_72965 == 32'h0000_0003 ? add_73003 : array_index_72997[3];
  assign array_update_73005[4] = add_72965 == 32'h0000_0004 ? add_73003 : array_index_72997[4];
  assign array_update_73005[5] = add_72965 == 32'h0000_0005 ? add_73003 : array_index_72997[5];
  assign array_update_73005[6] = add_72965 == 32'h0000_0006 ? add_73003 : array_index_72997[6];
  assign array_update_73005[7] = add_72965 == 32'h0000_0007 ? add_73003 : array_index_72997[7];
  assign array_update_73005[8] = add_72965 == 32'h0000_0008 ? add_73003 : array_index_72997[8];
  assign array_update_73005[9] = add_72965 == 32'h0000_0009 ? add_73003 : array_index_72997[9];
  assign add_73006 = add_72993 + 32'h0000_0001;
  assign array_update_73007[0] = literal_72009 == 32'h0000_0000 ? array_update_73005 : array_update_72994[0];
  assign array_update_73007[1] = literal_72009 == 32'h0000_0001 ? array_update_73005 : array_update_72994[1];
  assign array_update_73007[2] = literal_72009 == 32'h0000_0002 ? array_update_73005 : array_update_72994[2];
  assign array_update_73007[3] = literal_72009 == 32'h0000_0003 ? array_update_73005 : array_update_72994[3];
  assign array_update_73007[4] = literal_72009 == 32'h0000_0004 ? array_update_73005 : array_update_72994[4];
  assign array_update_73007[5] = literal_72009 == 32'h0000_0005 ? array_update_73005 : array_update_72994[5];
  assign array_update_73007[6] = literal_72009 == 32'h0000_0006 ? array_update_73005 : array_update_72994[6];
  assign array_update_73007[7] = literal_72009 == 32'h0000_0007 ? array_update_73005 : array_update_72994[7];
  assign array_update_73007[8] = literal_72009 == 32'h0000_0008 ? array_update_73005 : array_update_72994[8];
  assign array_update_73007[9] = literal_72009 == 32'h0000_0009 ? array_update_73005 : array_update_72994[9];
  assign array_index_73009 = array_update_72021[add_73006 > 32'h0000_0009 ? 4'h9 : add_73006[3:0]];
  assign array_index_73010 = array_update_73007[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_73014 = smul32b_32b_x_32b(array_index_72024[add_73006 > 32'h0000_0009 ? 4'h9 : add_73006[3:0]], array_index_73009[add_72965 > 32'h0000_0009 ? 4'h9 : add_72965[3:0]]);
  assign add_73016 = array_index_73010[add_72965 > 32'h0000_0009 ? 4'h9 : add_72965[3:0]] + smul_73014;
  assign array_update_73018[0] = add_72965 == 32'h0000_0000 ? add_73016 : array_index_73010[0];
  assign array_update_73018[1] = add_72965 == 32'h0000_0001 ? add_73016 : array_index_73010[1];
  assign array_update_73018[2] = add_72965 == 32'h0000_0002 ? add_73016 : array_index_73010[2];
  assign array_update_73018[3] = add_72965 == 32'h0000_0003 ? add_73016 : array_index_73010[3];
  assign array_update_73018[4] = add_72965 == 32'h0000_0004 ? add_73016 : array_index_73010[4];
  assign array_update_73018[5] = add_72965 == 32'h0000_0005 ? add_73016 : array_index_73010[5];
  assign array_update_73018[6] = add_72965 == 32'h0000_0006 ? add_73016 : array_index_73010[6];
  assign array_update_73018[7] = add_72965 == 32'h0000_0007 ? add_73016 : array_index_73010[7];
  assign array_update_73018[8] = add_72965 == 32'h0000_0008 ? add_73016 : array_index_73010[8];
  assign array_update_73018[9] = add_72965 == 32'h0000_0009 ? add_73016 : array_index_73010[9];
  assign add_73019 = add_73006 + 32'h0000_0001;
  assign array_update_73020[0] = literal_72009 == 32'h0000_0000 ? array_update_73018 : array_update_73007[0];
  assign array_update_73020[1] = literal_72009 == 32'h0000_0001 ? array_update_73018 : array_update_73007[1];
  assign array_update_73020[2] = literal_72009 == 32'h0000_0002 ? array_update_73018 : array_update_73007[2];
  assign array_update_73020[3] = literal_72009 == 32'h0000_0003 ? array_update_73018 : array_update_73007[3];
  assign array_update_73020[4] = literal_72009 == 32'h0000_0004 ? array_update_73018 : array_update_73007[4];
  assign array_update_73020[5] = literal_72009 == 32'h0000_0005 ? array_update_73018 : array_update_73007[5];
  assign array_update_73020[6] = literal_72009 == 32'h0000_0006 ? array_update_73018 : array_update_73007[6];
  assign array_update_73020[7] = literal_72009 == 32'h0000_0007 ? array_update_73018 : array_update_73007[7];
  assign array_update_73020[8] = literal_72009 == 32'h0000_0008 ? array_update_73018 : array_update_73007[8];
  assign array_update_73020[9] = literal_72009 == 32'h0000_0009 ? array_update_73018 : array_update_73007[9];
  assign array_index_73022 = array_update_72021[add_73019 > 32'h0000_0009 ? 4'h9 : add_73019[3:0]];
  assign array_index_73023 = array_update_73020[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_73027 = smul32b_32b_x_32b(array_index_72024[add_73019 > 32'h0000_0009 ? 4'h9 : add_73019[3:0]], array_index_73022[add_72965 > 32'h0000_0009 ? 4'h9 : add_72965[3:0]]);
  assign add_73029 = array_index_73023[add_72965 > 32'h0000_0009 ? 4'h9 : add_72965[3:0]] + smul_73027;
  assign array_update_73031[0] = add_72965 == 32'h0000_0000 ? add_73029 : array_index_73023[0];
  assign array_update_73031[1] = add_72965 == 32'h0000_0001 ? add_73029 : array_index_73023[1];
  assign array_update_73031[2] = add_72965 == 32'h0000_0002 ? add_73029 : array_index_73023[2];
  assign array_update_73031[3] = add_72965 == 32'h0000_0003 ? add_73029 : array_index_73023[3];
  assign array_update_73031[4] = add_72965 == 32'h0000_0004 ? add_73029 : array_index_73023[4];
  assign array_update_73031[5] = add_72965 == 32'h0000_0005 ? add_73029 : array_index_73023[5];
  assign array_update_73031[6] = add_72965 == 32'h0000_0006 ? add_73029 : array_index_73023[6];
  assign array_update_73031[7] = add_72965 == 32'h0000_0007 ? add_73029 : array_index_73023[7];
  assign array_update_73031[8] = add_72965 == 32'h0000_0008 ? add_73029 : array_index_73023[8];
  assign array_update_73031[9] = add_72965 == 32'h0000_0009 ? add_73029 : array_index_73023[9];
  assign add_73032 = add_73019 + 32'h0000_0001;
  assign array_update_73033[0] = literal_72009 == 32'h0000_0000 ? array_update_73031 : array_update_73020[0];
  assign array_update_73033[1] = literal_72009 == 32'h0000_0001 ? array_update_73031 : array_update_73020[1];
  assign array_update_73033[2] = literal_72009 == 32'h0000_0002 ? array_update_73031 : array_update_73020[2];
  assign array_update_73033[3] = literal_72009 == 32'h0000_0003 ? array_update_73031 : array_update_73020[3];
  assign array_update_73033[4] = literal_72009 == 32'h0000_0004 ? array_update_73031 : array_update_73020[4];
  assign array_update_73033[5] = literal_72009 == 32'h0000_0005 ? array_update_73031 : array_update_73020[5];
  assign array_update_73033[6] = literal_72009 == 32'h0000_0006 ? array_update_73031 : array_update_73020[6];
  assign array_update_73033[7] = literal_72009 == 32'h0000_0007 ? array_update_73031 : array_update_73020[7];
  assign array_update_73033[8] = literal_72009 == 32'h0000_0008 ? array_update_73031 : array_update_73020[8];
  assign array_update_73033[9] = literal_72009 == 32'h0000_0009 ? array_update_73031 : array_update_73020[9];
  assign array_index_73035 = array_update_72021[add_73032 > 32'h0000_0009 ? 4'h9 : add_73032[3:0]];
  assign array_index_73036 = array_update_73033[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_73040 = smul32b_32b_x_32b(array_index_72024[add_73032 > 32'h0000_0009 ? 4'h9 : add_73032[3:0]], array_index_73035[add_72965 > 32'h0000_0009 ? 4'h9 : add_72965[3:0]]);
  assign add_73042 = array_index_73036[add_72965 > 32'h0000_0009 ? 4'h9 : add_72965[3:0]] + smul_73040;
  assign array_update_73044[0] = add_72965 == 32'h0000_0000 ? add_73042 : array_index_73036[0];
  assign array_update_73044[1] = add_72965 == 32'h0000_0001 ? add_73042 : array_index_73036[1];
  assign array_update_73044[2] = add_72965 == 32'h0000_0002 ? add_73042 : array_index_73036[2];
  assign array_update_73044[3] = add_72965 == 32'h0000_0003 ? add_73042 : array_index_73036[3];
  assign array_update_73044[4] = add_72965 == 32'h0000_0004 ? add_73042 : array_index_73036[4];
  assign array_update_73044[5] = add_72965 == 32'h0000_0005 ? add_73042 : array_index_73036[5];
  assign array_update_73044[6] = add_72965 == 32'h0000_0006 ? add_73042 : array_index_73036[6];
  assign array_update_73044[7] = add_72965 == 32'h0000_0007 ? add_73042 : array_index_73036[7];
  assign array_update_73044[8] = add_72965 == 32'h0000_0008 ? add_73042 : array_index_73036[8];
  assign array_update_73044[9] = add_72965 == 32'h0000_0009 ? add_73042 : array_index_73036[9];
  assign add_73045 = add_73032 + 32'h0000_0001;
  assign array_update_73046[0] = literal_72009 == 32'h0000_0000 ? array_update_73044 : array_update_73033[0];
  assign array_update_73046[1] = literal_72009 == 32'h0000_0001 ? array_update_73044 : array_update_73033[1];
  assign array_update_73046[2] = literal_72009 == 32'h0000_0002 ? array_update_73044 : array_update_73033[2];
  assign array_update_73046[3] = literal_72009 == 32'h0000_0003 ? array_update_73044 : array_update_73033[3];
  assign array_update_73046[4] = literal_72009 == 32'h0000_0004 ? array_update_73044 : array_update_73033[4];
  assign array_update_73046[5] = literal_72009 == 32'h0000_0005 ? array_update_73044 : array_update_73033[5];
  assign array_update_73046[6] = literal_72009 == 32'h0000_0006 ? array_update_73044 : array_update_73033[6];
  assign array_update_73046[7] = literal_72009 == 32'h0000_0007 ? array_update_73044 : array_update_73033[7];
  assign array_update_73046[8] = literal_72009 == 32'h0000_0008 ? array_update_73044 : array_update_73033[8];
  assign array_update_73046[9] = literal_72009 == 32'h0000_0009 ? array_update_73044 : array_update_73033[9];
  assign array_index_73048 = array_update_72021[add_73045 > 32'h0000_0009 ? 4'h9 : add_73045[3:0]];
  assign array_index_73049 = array_update_73046[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_73053 = smul32b_32b_x_32b(array_index_72024[add_73045 > 32'h0000_0009 ? 4'h9 : add_73045[3:0]], array_index_73048[add_72965 > 32'h0000_0009 ? 4'h9 : add_72965[3:0]]);
  assign add_73055 = array_index_73049[add_72965 > 32'h0000_0009 ? 4'h9 : add_72965[3:0]] + smul_73053;
  assign array_update_73057[0] = add_72965 == 32'h0000_0000 ? add_73055 : array_index_73049[0];
  assign array_update_73057[1] = add_72965 == 32'h0000_0001 ? add_73055 : array_index_73049[1];
  assign array_update_73057[2] = add_72965 == 32'h0000_0002 ? add_73055 : array_index_73049[2];
  assign array_update_73057[3] = add_72965 == 32'h0000_0003 ? add_73055 : array_index_73049[3];
  assign array_update_73057[4] = add_72965 == 32'h0000_0004 ? add_73055 : array_index_73049[4];
  assign array_update_73057[5] = add_72965 == 32'h0000_0005 ? add_73055 : array_index_73049[5];
  assign array_update_73057[6] = add_72965 == 32'h0000_0006 ? add_73055 : array_index_73049[6];
  assign array_update_73057[7] = add_72965 == 32'h0000_0007 ? add_73055 : array_index_73049[7];
  assign array_update_73057[8] = add_72965 == 32'h0000_0008 ? add_73055 : array_index_73049[8];
  assign array_update_73057[9] = add_72965 == 32'h0000_0009 ? add_73055 : array_index_73049[9];
  assign add_73058 = add_73045 + 32'h0000_0001;
  assign array_update_73059[0] = literal_72009 == 32'h0000_0000 ? array_update_73057 : array_update_73046[0];
  assign array_update_73059[1] = literal_72009 == 32'h0000_0001 ? array_update_73057 : array_update_73046[1];
  assign array_update_73059[2] = literal_72009 == 32'h0000_0002 ? array_update_73057 : array_update_73046[2];
  assign array_update_73059[3] = literal_72009 == 32'h0000_0003 ? array_update_73057 : array_update_73046[3];
  assign array_update_73059[4] = literal_72009 == 32'h0000_0004 ? array_update_73057 : array_update_73046[4];
  assign array_update_73059[5] = literal_72009 == 32'h0000_0005 ? array_update_73057 : array_update_73046[5];
  assign array_update_73059[6] = literal_72009 == 32'h0000_0006 ? array_update_73057 : array_update_73046[6];
  assign array_update_73059[7] = literal_72009 == 32'h0000_0007 ? array_update_73057 : array_update_73046[7];
  assign array_update_73059[8] = literal_72009 == 32'h0000_0008 ? array_update_73057 : array_update_73046[8];
  assign array_update_73059[9] = literal_72009 == 32'h0000_0009 ? array_update_73057 : array_update_73046[9];
  assign array_index_73061 = array_update_72021[add_73058 > 32'h0000_0009 ? 4'h9 : add_73058[3:0]];
  assign array_index_73062 = array_update_73059[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_73066 = smul32b_32b_x_32b(array_index_72024[add_73058 > 32'h0000_0009 ? 4'h9 : add_73058[3:0]], array_index_73061[add_72965 > 32'h0000_0009 ? 4'h9 : add_72965[3:0]]);
  assign add_73068 = array_index_73062[add_72965 > 32'h0000_0009 ? 4'h9 : add_72965[3:0]] + smul_73066;
  assign array_update_73070[0] = add_72965 == 32'h0000_0000 ? add_73068 : array_index_73062[0];
  assign array_update_73070[1] = add_72965 == 32'h0000_0001 ? add_73068 : array_index_73062[1];
  assign array_update_73070[2] = add_72965 == 32'h0000_0002 ? add_73068 : array_index_73062[2];
  assign array_update_73070[3] = add_72965 == 32'h0000_0003 ? add_73068 : array_index_73062[3];
  assign array_update_73070[4] = add_72965 == 32'h0000_0004 ? add_73068 : array_index_73062[4];
  assign array_update_73070[5] = add_72965 == 32'h0000_0005 ? add_73068 : array_index_73062[5];
  assign array_update_73070[6] = add_72965 == 32'h0000_0006 ? add_73068 : array_index_73062[6];
  assign array_update_73070[7] = add_72965 == 32'h0000_0007 ? add_73068 : array_index_73062[7];
  assign array_update_73070[8] = add_72965 == 32'h0000_0008 ? add_73068 : array_index_73062[8];
  assign array_update_73070[9] = add_72965 == 32'h0000_0009 ? add_73068 : array_index_73062[9];
  assign add_73071 = add_73058 + 32'h0000_0001;
  assign array_update_73072[0] = literal_72009 == 32'h0000_0000 ? array_update_73070 : array_update_73059[0];
  assign array_update_73072[1] = literal_72009 == 32'h0000_0001 ? array_update_73070 : array_update_73059[1];
  assign array_update_73072[2] = literal_72009 == 32'h0000_0002 ? array_update_73070 : array_update_73059[2];
  assign array_update_73072[3] = literal_72009 == 32'h0000_0003 ? array_update_73070 : array_update_73059[3];
  assign array_update_73072[4] = literal_72009 == 32'h0000_0004 ? array_update_73070 : array_update_73059[4];
  assign array_update_73072[5] = literal_72009 == 32'h0000_0005 ? array_update_73070 : array_update_73059[5];
  assign array_update_73072[6] = literal_72009 == 32'h0000_0006 ? array_update_73070 : array_update_73059[6];
  assign array_update_73072[7] = literal_72009 == 32'h0000_0007 ? array_update_73070 : array_update_73059[7];
  assign array_update_73072[8] = literal_72009 == 32'h0000_0008 ? array_update_73070 : array_update_73059[8];
  assign array_update_73072[9] = literal_72009 == 32'h0000_0009 ? array_update_73070 : array_update_73059[9];
  assign array_index_73074 = array_update_72021[add_73071 > 32'h0000_0009 ? 4'h9 : add_73071[3:0]];
  assign array_index_73075 = array_update_73072[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_73079 = smul32b_32b_x_32b(array_index_72024[add_73071 > 32'h0000_0009 ? 4'h9 : add_73071[3:0]], array_index_73074[add_72965 > 32'h0000_0009 ? 4'h9 : add_72965[3:0]]);
  assign add_73081 = array_index_73075[add_72965 > 32'h0000_0009 ? 4'h9 : add_72965[3:0]] + smul_73079;
  assign array_update_73083[0] = add_72965 == 32'h0000_0000 ? add_73081 : array_index_73075[0];
  assign array_update_73083[1] = add_72965 == 32'h0000_0001 ? add_73081 : array_index_73075[1];
  assign array_update_73083[2] = add_72965 == 32'h0000_0002 ? add_73081 : array_index_73075[2];
  assign array_update_73083[3] = add_72965 == 32'h0000_0003 ? add_73081 : array_index_73075[3];
  assign array_update_73083[4] = add_72965 == 32'h0000_0004 ? add_73081 : array_index_73075[4];
  assign array_update_73083[5] = add_72965 == 32'h0000_0005 ? add_73081 : array_index_73075[5];
  assign array_update_73083[6] = add_72965 == 32'h0000_0006 ? add_73081 : array_index_73075[6];
  assign array_update_73083[7] = add_72965 == 32'h0000_0007 ? add_73081 : array_index_73075[7];
  assign array_update_73083[8] = add_72965 == 32'h0000_0008 ? add_73081 : array_index_73075[8];
  assign array_update_73083[9] = add_72965 == 32'h0000_0009 ? add_73081 : array_index_73075[9];
  assign add_73084 = add_73071 + 32'h0000_0001;
  assign array_update_73085[0] = literal_72009 == 32'h0000_0000 ? array_update_73083 : array_update_73072[0];
  assign array_update_73085[1] = literal_72009 == 32'h0000_0001 ? array_update_73083 : array_update_73072[1];
  assign array_update_73085[2] = literal_72009 == 32'h0000_0002 ? array_update_73083 : array_update_73072[2];
  assign array_update_73085[3] = literal_72009 == 32'h0000_0003 ? array_update_73083 : array_update_73072[3];
  assign array_update_73085[4] = literal_72009 == 32'h0000_0004 ? array_update_73083 : array_update_73072[4];
  assign array_update_73085[5] = literal_72009 == 32'h0000_0005 ? array_update_73083 : array_update_73072[5];
  assign array_update_73085[6] = literal_72009 == 32'h0000_0006 ? array_update_73083 : array_update_73072[6];
  assign array_update_73085[7] = literal_72009 == 32'h0000_0007 ? array_update_73083 : array_update_73072[7];
  assign array_update_73085[8] = literal_72009 == 32'h0000_0008 ? array_update_73083 : array_update_73072[8];
  assign array_update_73085[9] = literal_72009 == 32'h0000_0009 ? array_update_73083 : array_update_73072[9];
  assign array_index_73087 = array_update_72021[add_73084 > 32'h0000_0009 ? 4'h9 : add_73084[3:0]];
  assign array_index_73088 = array_update_73085[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_73092 = smul32b_32b_x_32b(array_index_72024[add_73084 > 32'h0000_0009 ? 4'h9 : add_73084[3:0]], array_index_73087[add_72965 > 32'h0000_0009 ? 4'h9 : add_72965[3:0]]);
  assign add_73094 = array_index_73088[add_72965 > 32'h0000_0009 ? 4'h9 : add_72965[3:0]] + smul_73092;
  assign array_update_73095[0] = add_72965 == 32'h0000_0000 ? add_73094 : array_index_73088[0];
  assign array_update_73095[1] = add_72965 == 32'h0000_0001 ? add_73094 : array_index_73088[1];
  assign array_update_73095[2] = add_72965 == 32'h0000_0002 ? add_73094 : array_index_73088[2];
  assign array_update_73095[3] = add_72965 == 32'h0000_0003 ? add_73094 : array_index_73088[3];
  assign array_update_73095[4] = add_72965 == 32'h0000_0004 ? add_73094 : array_index_73088[4];
  assign array_update_73095[5] = add_72965 == 32'h0000_0005 ? add_73094 : array_index_73088[5];
  assign array_update_73095[6] = add_72965 == 32'h0000_0006 ? add_73094 : array_index_73088[6];
  assign array_update_73095[7] = add_72965 == 32'h0000_0007 ? add_73094 : array_index_73088[7];
  assign array_update_73095[8] = add_72965 == 32'h0000_0008 ? add_73094 : array_index_73088[8];
  assign array_update_73095[9] = add_72965 == 32'h0000_0009 ? add_73094 : array_index_73088[9];
  assign array_update_73096[0] = literal_72009 == 32'h0000_0000 ? array_update_73095 : array_update_73085[0];
  assign array_update_73096[1] = literal_72009 == 32'h0000_0001 ? array_update_73095 : array_update_73085[1];
  assign array_update_73096[2] = literal_72009 == 32'h0000_0002 ? array_update_73095 : array_update_73085[2];
  assign array_update_73096[3] = literal_72009 == 32'h0000_0003 ? array_update_73095 : array_update_73085[3];
  assign array_update_73096[4] = literal_72009 == 32'h0000_0004 ? array_update_73095 : array_update_73085[4];
  assign array_update_73096[5] = literal_72009 == 32'h0000_0005 ? array_update_73095 : array_update_73085[5];
  assign array_update_73096[6] = literal_72009 == 32'h0000_0006 ? array_update_73095 : array_update_73085[6];
  assign array_update_73096[7] = literal_72009 == 32'h0000_0007 ? array_update_73095 : array_update_73085[7];
  assign array_update_73096[8] = literal_72009 == 32'h0000_0008 ? array_update_73095 : array_update_73085[8];
  assign array_update_73096[9] = literal_72009 == 32'h0000_0009 ? array_update_73095 : array_update_73085[9];
  assign array_index_73098 = array_update_73096[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign add_73100 = add_72965 + 32'h0000_0001;
  assign array_update_73101[0] = add_73100 == 32'h0000_0000 ? 32'h0000_0000 : array_index_73098[0];
  assign array_update_73101[1] = add_73100 == 32'h0000_0001 ? 32'h0000_0000 : array_index_73098[1];
  assign array_update_73101[2] = add_73100 == 32'h0000_0002 ? 32'h0000_0000 : array_index_73098[2];
  assign array_update_73101[3] = add_73100 == 32'h0000_0003 ? 32'h0000_0000 : array_index_73098[3];
  assign array_update_73101[4] = add_73100 == 32'h0000_0004 ? 32'h0000_0000 : array_index_73098[4];
  assign array_update_73101[5] = add_73100 == 32'h0000_0005 ? 32'h0000_0000 : array_index_73098[5];
  assign array_update_73101[6] = add_73100 == 32'h0000_0006 ? 32'h0000_0000 : array_index_73098[6];
  assign array_update_73101[7] = add_73100 == 32'h0000_0007 ? 32'h0000_0000 : array_index_73098[7];
  assign array_update_73101[8] = add_73100 == 32'h0000_0008 ? 32'h0000_0000 : array_index_73098[8];
  assign array_update_73101[9] = add_73100 == 32'h0000_0009 ? 32'h0000_0000 : array_index_73098[9];
  assign literal_73102 = 32'h0000_0000;
  assign array_update_73103[0] = literal_72009 == 32'h0000_0000 ? array_update_73101 : array_update_73096[0];
  assign array_update_73103[1] = literal_72009 == 32'h0000_0001 ? array_update_73101 : array_update_73096[1];
  assign array_update_73103[2] = literal_72009 == 32'h0000_0002 ? array_update_73101 : array_update_73096[2];
  assign array_update_73103[3] = literal_72009 == 32'h0000_0003 ? array_update_73101 : array_update_73096[3];
  assign array_update_73103[4] = literal_72009 == 32'h0000_0004 ? array_update_73101 : array_update_73096[4];
  assign array_update_73103[5] = literal_72009 == 32'h0000_0005 ? array_update_73101 : array_update_73096[5];
  assign array_update_73103[6] = literal_72009 == 32'h0000_0006 ? array_update_73101 : array_update_73096[6];
  assign array_update_73103[7] = literal_72009 == 32'h0000_0007 ? array_update_73101 : array_update_73096[7];
  assign array_update_73103[8] = literal_72009 == 32'h0000_0008 ? array_update_73101 : array_update_73096[8];
  assign array_update_73103[9] = literal_72009 == 32'h0000_0009 ? array_update_73101 : array_update_73096[9];
  assign array_index_73105 = array_update_72021[literal_73102 > 32'h0000_0009 ? 4'h9 : literal_73102[3:0]];
  assign array_index_73106 = array_update_73103[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_73110 = smul32b_32b_x_32b(array_index_72024[literal_73102 > 32'h0000_0009 ? 4'h9 : literal_73102[3:0]], array_index_73105[add_73100 > 32'h0000_0009 ? 4'h9 : add_73100[3:0]]);
  assign add_73112 = array_index_73106[add_73100 > 32'h0000_0009 ? 4'h9 : add_73100[3:0]] + smul_73110;
  assign array_update_73114[0] = add_73100 == 32'h0000_0000 ? add_73112 : array_index_73106[0];
  assign array_update_73114[1] = add_73100 == 32'h0000_0001 ? add_73112 : array_index_73106[1];
  assign array_update_73114[2] = add_73100 == 32'h0000_0002 ? add_73112 : array_index_73106[2];
  assign array_update_73114[3] = add_73100 == 32'h0000_0003 ? add_73112 : array_index_73106[3];
  assign array_update_73114[4] = add_73100 == 32'h0000_0004 ? add_73112 : array_index_73106[4];
  assign array_update_73114[5] = add_73100 == 32'h0000_0005 ? add_73112 : array_index_73106[5];
  assign array_update_73114[6] = add_73100 == 32'h0000_0006 ? add_73112 : array_index_73106[6];
  assign array_update_73114[7] = add_73100 == 32'h0000_0007 ? add_73112 : array_index_73106[7];
  assign array_update_73114[8] = add_73100 == 32'h0000_0008 ? add_73112 : array_index_73106[8];
  assign array_update_73114[9] = add_73100 == 32'h0000_0009 ? add_73112 : array_index_73106[9];
  assign add_73115 = literal_73102 + 32'h0000_0001;
  assign array_update_73116[0] = literal_72009 == 32'h0000_0000 ? array_update_73114 : array_update_73103[0];
  assign array_update_73116[1] = literal_72009 == 32'h0000_0001 ? array_update_73114 : array_update_73103[1];
  assign array_update_73116[2] = literal_72009 == 32'h0000_0002 ? array_update_73114 : array_update_73103[2];
  assign array_update_73116[3] = literal_72009 == 32'h0000_0003 ? array_update_73114 : array_update_73103[3];
  assign array_update_73116[4] = literal_72009 == 32'h0000_0004 ? array_update_73114 : array_update_73103[4];
  assign array_update_73116[5] = literal_72009 == 32'h0000_0005 ? array_update_73114 : array_update_73103[5];
  assign array_update_73116[6] = literal_72009 == 32'h0000_0006 ? array_update_73114 : array_update_73103[6];
  assign array_update_73116[7] = literal_72009 == 32'h0000_0007 ? array_update_73114 : array_update_73103[7];
  assign array_update_73116[8] = literal_72009 == 32'h0000_0008 ? array_update_73114 : array_update_73103[8];
  assign array_update_73116[9] = literal_72009 == 32'h0000_0009 ? array_update_73114 : array_update_73103[9];
  assign array_index_73118 = array_update_72021[add_73115 > 32'h0000_0009 ? 4'h9 : add_73115[3:0]];
  assign array_index_73119 = array_update_73116[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_73123 = smul32b_32b_x_32b(array_index_72024[add_73115 > 32'h0000_0009 ? 4'h9 : add_73115[3:0]], array_index_73118[add_73100 > 32'h0000_0009 ? 4'h9 : add_73100[3:0]]);
  assign add_73125 = array_index_73119[add_73100 > 32'h0000_0009 ? 4'h9 : add_73100[3:0]] + smul_73123;
  assign array_update_73127[0] = add_73100 == 32'h0000_0000 ? add_73125 : array_index_73119[0];
  assign array_update_73127[1] = add_73100 == 32'h0000_0001 ? add_73125 : array_index_73119[1];
  assign array_update_73127[2] = add_73100 == 32'h0000_0002 ? add_73125 : array_index_73119[2];
  assign array_update_73127[3] = add_73100 == 32'h0000_0003 ? add_73125 : array_index_73119[3];
  assign array_update_73127[4] = add_73100 == 32'h0000_0004 ? add_73125 : array_index_73119[4];
  assign array_update_73127[5] = add_73100 == 32'h0000_0005 ? add_73125 : array_index_73119[5];
  assign array_update_73127[6] = add_73100 == 32'h0000_0006 ? add_73125 : array_index_73119[6];
  assign array_update_73127[7] = add_73100 == 32'h0000_0007 ? add_73125 : array_index_73119[7];
  assign array_update_73127[8] = add_73100 == 32'h0000_0008 ? add_73125 : array_index_73119[8];
  assign array_update_73127[9] = add_73100 == 32'h0000_0009 ? add_73125 : array_index_73119[9];
  assign add_73128 = add_73115 + 32'h0000_0001;
  assign array_update_73129[0] = literal_72009 == 32'h0000_0000 ? array_update_73127 : array_update_73116[0];
  assign array_update_73129[1] = literal_72009 == 32'h0000_0001 ? array_update_73127 : array_update_73116[1];
  assign array_update_73129[2] = literal_72009 == 32'h0000_0002 ? array_update_73127 : array_update_73116[2];
  assign array_update_73129[3] = literal_72009 == 32'h0000_0003 ? array_update_73127 : array_update_73116[3];
  assign array_update_73129[4] = literal_72009 == 32'h0000_0004 ? array_update_73127 : array_update_73116[4];
  assign array_update_73129[5] = literal_72009 == 32'h0000_0005 ? array_update_73127 : array_update_73116[5];
  assign array_update_73129[6] = literal_72009 == 32'h0000_0006 ? array_update_73127 : array_update_73116[6];
  assign array_update_73129[7] = literal_72009 == 32'h0000_0007 ? array_update_73127 : array_update_73116[7];
  assign array_update_73129[8] = literal_72009 == 32'h0000_0008 ? array_update_73127 : array_update_73116[8];
  assign array_update_73129[9] = literal_72009 == 32'h0000_0009 ? array_update_73127 : array_update_73116[9];
  assign array_index_73131 = array_update_72021[add_73128 > 32'h0000_0009 ? 4'h9 : add_73128[3:0]];
  assign array_index_73132 = array_update_73129[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_73136 = smul32b_32b_x_32b(array_index_72024[add_73128 > 32'h0000_0009 ? 4'h9 : add_73128[3:0]], array_index_73131[add_73100 > 32'h0000_0009 ? 4'h9 : add_73100[3:0]]);
  assign add_73138 = array_index_73132[add_73100 > 32'h0000_0009 ? 4'h9 : add_73100[3:0]] + smul_73136;
  assign array_update_73140[0] = add_73100 == 32'h0000_0000 ? add_73138 : array_index_73132[0];
  assign array_update_73140[1] = add_73100 == 32'h0000_0001 ? add_73138 : array_index_73132[1];
  assign array_update_73140[2] = add_73100 == 32'h0000_0002 ? add_73138 : array_index_73132[2];
  assign array_update_73140[3] = add_73100 == 32'h0000_0003 ? add_73138 : array_index_73132[3];
  assign array_update_73140[4] = add_73100 == 32'h0000_0004 ? add_73138 : array_index_73132[4];
  assign array_update_73140[5] = add_73100 == 32'h0000_0005 ? add_73138 : array_index_73132[5];
  assign array_update_73140[6] = add_73100 == 32'h0000_0006 ? add_73138 : array_index_73132[6];
  assign array_update_73140[7] = add_73100 == 32'h0000_0007 ? add_73138 : array_index_73132[7];
  assign array_update_73140[8] = add_73100 == 32'h0000_0008 ? add_73138 : array_index_73132[8];
  assign array_update_73140[9] = add_73100 == 32'h0000_0009 ? add_73138 : array_index_73132[9];
  assign add_73141 = add_73128 + 32'h0000_0001;
  assign array_update_73142[0] = literal_72009 == 32'h0000_0000 ? array_update_73140 : array_update_73129[0];
  assign array_update_73142[1] = literal_72009 == 32'h0000_0001 ? array_update_73140 : array_update_73129[1];
  assign array_update_73142[2] = literal_72009 == 32'h0000_0002 ? array_update_73140 : array_update_73129[2];
  assign array_update_73142[3] = literal_72009 == 32'h0000_0003 ? array_update_73140 : array_update_73129[3];
  assign array_update_73142[4] = literal_72009 == 32'h0000_0004 ? array_update_73140 : array_update_73129[4];
  assign array_update_73142[5] = literal_72009 == 32'h0000_0005 ? array_update_73140 : array_update_73129[5];
  assign array_update_73142[6] = literal_72009 == 32'h0000_0006 ? array_update_73140 : array_update_73129[6];
  assign array_update_73142[7] = literal_72009 == 32'h0000_0007 ? array_update_73140 : array_update_73129[7];
  assign array_update_73142[8] = literal_72009 == 32'h0000_0008 ? array_update_73140 : array_update_73129[8];
  assign array_update_73142[9] = literal_72009 == 32'h0000_0009 ? array_update_73140 : array_update_73129[9];
  assign array_index_73144 = array_update_72021[add_73141 > 32'h0000_0009 ? 4'h9 : add_73141[3:0]];
  assign array_index_73145 = array_update_73142[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_73149 = smul32b_32b_x_32b(array_index_72024[add_73141 > 32'h0000_0009 ? 4'h9 : add_73141[3:0]], array_index_73144[add_73100 > 32'h0000_0009 ? 4'h9 : add_73100[3:0]]);
  assign add_73151 = array_index_73145[add_73100 > 32'h0000_0009 ? 4'h9 : add_73100[3:0]] + smul_73149;
  assign array_update_73153[0] = add_73100 == 32'h0000_0000 ? add_73151 : array_index_73145[0];
  assign array_update_73153[1] = add_73100 == 32'h0000_0001 ? add_73151 : array_index_73145[1];
  assign array_update_73153[2] = add_73100 == 32'h0000_0002 ? add_73151 : array_index_73145[2];
  assign array_update_73153[3] = add_73100 == 32'h0000_0003 ? add_73151 : array_index_73145[3];
  assign array_update_73153[4] = add_73100 == 32'h0000_0004 ? add_73151 : array_index_73145[4];
  assign array_update_73153[5] = add_73100 == 32'h0000_0005 ? add_73151 : array_index_73145[5];
  assign array_update_73153[6] = add_73100 == 32'h0000_0006 ? add_73151 : array_index_73145[6];
  assign array_update_73153[7] = add_73100 == 32'h0000_0007 ? add_73151 : array_index_73145[7];
  assign array_update_73153[8] = add_73100 == 32'h0000_0008 ? add_73151 : array_index_73145[8];
  assign array_update_73153[9] = add_73100 == 32'h0000_0009 ? add_73151 : array_index_73145[9];
  assign add_73154 = add_73141 + 32'h0000_0001;
  assign array_update_73155[0] = literal_72009 == 32'h0000_0000 ? array_update_73153 : array_update_73142[0];
  assign array_update_73155[1] = literal_72009 == 32'h0000_0001 ? array_update_73153 : array_update_73142[1];
  assign array_update_73155[2] = literal_72009 == 32'h0000_0002 ? array_update_73153 : array_update_73142[2];
  assign array_update_73155[3] = literal_72009 == 32'h0000_0003 ? array_update_73153 : array_update_73142[3];
  assign array_update_73155[4] = literal_72009 == 32'h0000_0004 ? array_update_73153 : array_update_73142[4];
  assign array_update_73155[5] = literal_72009 == 32'h0000_0005 ? array_update_73153 : array_update_73142[5];
  assign array_update_73155[6] = literal_72009 == 32'h0000_0006 ? array_update_73153 : array_update_73142[6];
  assign array_update_73155[7] = literal_72009 == 32'h0000_0007 ? array_update_73153 : array_update_73142[7];
  assign array_update_73155[8] = literal_72009 == 32'h0000_0008 ? array_update_73153 : array_update_73142[8];
  assign array_update_73155[9] = literal_72009 == 32'h0000_0009 ? array_update_73153 : array_update_73142[9];
  assign array_index_73157 = array_update_72021[add_73154 > 32'h0000_0009 ? 4'h9 : add_73154[3:0]];
  assign array_index_73158 = array_update_73155[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_73162 = smul32b_32b_x_32b(array_index_72024[add_73154 > 32'h0000_0009 ? 4'h9 : add_73154[3:0]], array_index_73157[add_73100 > 32'h0000_0009 ? 4'h9 : add_73100[3:0]]);
  assign add_73164 = array_index_73158[add_73100 > 32'h0000_0009 ? 4'h9 : add_73100[3:0]] + smul_73162;
  assign array_update_73166[0] = add_73100 == 32'h0000_0000 ? add_73164 : array_index_73158[0];
  assign array_update_73166[1] = add_73100 == 32'h0000_0001 ? add_73164 : array_index_73158[1];
  assign array_update_73166[2] = add_73100 == 32'h0000_0002 ? add_73164 : array_index_73158[2];
  assign array_update_73166[3] = add_73100 == 32'h0000_0003 ? add_73164 : array_index_73158[3];
  assign array_update_73166[4] = add_73100 == 32'h0000_0004 ? add_73164 : array_index_73158[4];
  assign array_update_73166[5] = add_73100 == 32'h0000_0005 ? add_73164 : array_index_73158[5];
  assign array_update_73166[6] = add_73100 == 32'h0000_0006 ? add_73164 : array_index_73158[6];
  assign array_update_73166[7] = add_73100 == 32'h0000_0007 ? add_73164 : array_index_73158[7];
  assign array_update_73166[8] = add_73100 == 32'h0000_0008 ? add_73164 : array_index_73158[8];
  assign array_update_73166[9] = add_73100 == 32'h0000_0009 ? add_73164 : array_index_73158[9];
  assign add_73167 = add_73154 + 32'h0000_0001;
  assign array_update_73168[0] = literal_72009 == 32'h0000_0000 ? array_update_73166 : array_update_73155[0];
  assign array_update_73168[1] = literal_72009 == 32'h0000_0001 ? array_update_73166 : array_update_73155[1];
  assign array_update_73168[2] = literal_72009 == 32'h0000_0002 ? array_update_73166 : array_update_73155[2];
  assign array_update_73168[3] = literal_72009 == 32'h0000_0003 ? array_update_73166 : array_update_73155[3];
  assign array_update_73168[4] = literal_72009 == 32'h0000_0004 ? array_update_73166 : array_update_73155[4];
  assign array_update_73168[5] = literal_72009 == 32'h0000_0005 ? array_update_73166 : array_update_73155[5];
  assign array_update_73168[6] = literal_72009 == 32'h0000_0006 ? array_update_73166 : array_update_73155[6];
  assign array_update_73168[7] = literal_72009 == 32'h0000_0007 ? array_update_73166 : array_update_73155[7];
  assign array_update_73168[8] = literal_72009 == 32'h0000_0008 ? array_update_73166 : array_update_73155[8];
  assign array_update_73168[9] = literal_72009 == 32'h0000_0009 ? array_update_73166 : array_update_73155[9];
  assign array_index_73170 = array_update_72021[add_73167 > 32'h0000_0009 ? 4'h9 : add_73167[3:0]];
  assign array_index_73171 = array_update_73168[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_73175 = smul32b_32b_x_32b(array_index_72024[add_73167 > 32'h0000_0009 ? 4'h9 : add_73167[3:0]], array_index_73170[add_73100 > 32'h0000_0009 ? 4'h9 : add_73100[3:0]]);
  assign add_73177 = array_index_73171[add_73100 > 32'h0000_0009 ? 4'h9 : add_73100[3:0]] + smul_73175;
  assign array_update_73179[0] = add_73100 == 32'h0000_0000 ? add_73177 : array_index_73171[0];
  assign array_update_73179[1] = add_73100 == 32'h0000_0001 ? add_73177 : array_index_73171[1];
  assign array_update_73179[2] = add_73100 == 32'h0000_0002 ? add_73177 : array_index_73171[2];
  assign array_update_73179[3] = add_73100 == 32'h0000_0003 ? add_73177 : array_index_73171[3];
  assign array_update_73179[4] = add_73100 == 32'h0000_0004 ? add_73177 : array_index_73171[4];
  assign array_update_73179[5] = add_73100 == 32'h0000_0005 ? add_73177 : array_index_73171[5];
  assign array_update_73179[6] = add_73100 == 32'h0000_0006 ? add_73177 : array_index_73171[6];
  assign array_update_73179[7] = add_73100 == 32'h0000_0007 ? add_73177 : array_index_73171[7];
  assign array_update_73179[8] = add_73100 == 32'h0000_0008 ? add_73177 : array_index_73171[8];
  assign array_update_73179[9] = add_73100 == 32'h0000_0009 ? add_73177 : array_index_73171[9];
  assign add_73180 = add_73167 + 32'h0000_0001;
  assign array_update_73181[0] = literal_72009 == 32'h0000_0000 ? array_update_73179 : array_update_73168[0];
  assign array_update_73181[1] = literal_72009 == 32'h0000_0001 ? array_update_73179 : array_update_73168[1];
  assign array_update_73181[2] = literal_72009 == 32'h0000_0002 ? array_update_73179 : array_update_73168[2];
  assign array_update_73181[3] = literal_72009 == 32'h0000_0003 ? array_update_73179 : array_update_73168[3];
  assign array_update_73181[4] = literal_72009 == 32'h0000_0004 ? array_update_73179 : array_update_73168[4];
  assign array_update_73181[5] = literal_72009 == 32'h0000_0005 ? array_update_73179 : array_update_73168[5];
  assign array_update_73181[6] = literal_72009 == 32'h0000_0006 ? array_update_73179 : array_update_73168[6];
  assign array_update_73181[7] = literal_72009 == 32'h0000_0007 ? array_update_73179 : array_update_73168[7];
  assign array_update_73181[8] = literal_72009 == 32'h0000_0008 ? array_update_73179 : array_update_73168[8];
  assign array_update_73181[9] = literal_72009 == 32'h0000_0009 ? array_update_73179 : array_update_73168[9];
  assign array_index_73183 = array_update_72021[add_73180 > 32'h0000_0009 ? 4'h9 : add_73180[3:0]];
  assign array_index_73184 = array_update_73181[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_73188 = smul32b_32b_x_32b(array_index_72024[add_73180 > 32'h0000_0009 ? 4'h9 : add_73180[3:0]], array_index_73183[add_73100 > 32'h0000_0009 ? 4'h9 : add_73100[3:0]]);
  assign add_73190 = array_index_73184[add_73100 > 32'h0000_0009 ? 4'h9 : add_73100[3:0]] + smul_73188;
  assign array_update_73192[0] = add_73100 == 32'h0000_0000 ? add_73190 : array_index_73184[0];
  assign array_update_73192[1] = add_73100 == 32'h0000_0001 ? add_73190 : array_index_73184[1];
  assign array_update_73192[2] = add_73100 == 32'h0000_0002 ? add_73190 : array_index_73184[2];
  assign array_update_73192[3] = add_73100 == 32'h0000_0003 ? add_73190 : array_index_73184[3];
  assign array_update_73192[4] = add_73100 == 32'h0000_0004 ? add_73190 : array_index_73184[4];
  assign array_update_73192[5] = add_73100 == 32'h0000_0005 ? add_73190 : array_index_73184[5];
  assign array_update_73192[6] = add_73100 == 32'h0000_0006 ? add_73190 : array_index_73184[6];
  assign array_update_73192[7] = add_73100 == 32'h0000_0007 ? add_73190 : array_index_73184[7];
  assign array_update_73192[8] = add_73100 == 32'h0000_0008 ? add_73190 : array_index_73184[8];
  assign array_update_73192[9] = add_73100 == 32'h0000_0009 ? add_73190 : array_index_73184[9];
  assign add_73193 = add_73180 + 32'h0000_0001;
  assign array_update_73194[0] = literal_72009 == 32'h0000_0000 ? array_update_73192 : array_update_73181[0];
  assign array_update_73194[1] = literal_72009 == 32'h0000_0001 ? array_update_73192 : array_update_73181[1];
  assign array_update_73194[2] = literal_72009 == 32'h0000_0002 ? array_update_73192 : array_update_73181[2];
  assign array_update_73194[3] = literal_72009 == 32'h0000_0003 ? array_update_73192 : array_update_73181[3];
  assign array_update_73194[4] = literal_72009 == 32'h0000_0004 ? array_update_73192 : array_update_73181[4];
  assign array_update_73194[5] = literal_72009 == 32'h0000_0005 ? array_update_73192 : array_update_73181[5];
  assign array_update_73194[6] = literal_72009 == 32'h0000_0006 ? array_update_73192 : array_update_73181[6];
  assign array_update_73194[7] = literal_72009 == 32'h0000_0007 ? array_update_73192 : array_update_73181[7];
  assign array_update_73194[8] = literal_72009 == 32'h0000_0008 ? array_update_73192 : array_update_73181[8];
  assign array_update_73194[9] = literal_72009 == 32'h0000_0009 ? array_update_73192 : array_update_73181[9];
  assign array_index_73196 = array_update_72021[add_73193 > 32'h0000_0009 ? 4'h9 : add_73193[3:0]];
  assign array_index_73197 = array_update_73194[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_73201 = smul32b_32b_x_32b(array_index_72024[add_73193 > 32'h0000_0009 ? 4'h9 : add_73193[3:0]], array_index_73196[add_73100 > 32'h0000_0009 ? 4'h9 : add_73100[3:0]]);
  assign add_73203 = array_index_73197[add_73100 > 32'h0000_0009 ? 4'h9 : add_73100[3:0]] + smul_73201;
  assign array_update_73205[0] = add_73100 == 32'h0000_0000 ? add_73203 : array_index_73197[0];
  assign array_update_73205[1] = add_73100 == 32'h0000_0001 ? add_73203 : array_index_73197[1];
  assign array_update_73205[2] = add_73100 == 32'h0000_0002 ? add_73203 : array_index_73197[2];
  assign array_update_73205[3] = add_73100 == 32'h0000_0003 ? add_73203 : array_index_73197[3];
  assign array_update_73205[4] = add_73100 == 32'h0000_0004 ? add_73203 : array_index_73197[4];
  assign array_update_73205[5] = add_73100 == 32'h0000_0005 ? add_73203 : array_index_73197[5];
  assign array_update_73205[6] = add_73100 == 32'h0000_0006 ? add_73203 : array_index_73197[6];
  assign array_update_73205[7] = add_73100 == 32'h0000_0007 ? add_73203 : array_index_73197[7];
  assign array_update_73205[8] = add_73100 == 32'h0000_0008 ? add_73203 : array_index_73197[8];
  assign array_update_73205[9] = add_73100 == 32'h0000_0009 ? add_73203 : array_index_73197[9];
  assign add_73206 = add_73193 + 32'h0000_0001;
  assign array_update_73207[0] = literal_72009 == 32'h0000_0000 ? array_update_73205 : array_update_73194[0];
  assign array_update_73207[1] = literal_72009 == 32'h0000_0001 ? array_update_73205 : array_update_73194[1];
  assign array_update_73207[2] = literal_72009 == 32'h0000_0002 ? array_update_73205 : array_update_73194[2];
  assign array_update_73207[3] = literal_72009 == 32'h0000_0003 ? array_update_73205 : array_update_73194[3];
  assign array_update_73207[4] = literal_72009 == 32'h0000_0004 ? array_update_73205 : array_update_73194[4];
  assign array_update_73207[5] = literal_72009 == 32'h0000_0005 ? array_update_73205 : array_update_73194[5];
  assign array_update_73207[6] = literal_72009 == 32'h0000_0006 ? array_update_73205 : array_update_73194[6];
  assign array_update_73207[7] = literal_72009 == 32'h0000_0007 ? array_update_73205 : array_update_73194[7];
  assign array_update_73207[8] = literal_72009 == 32'h0000_0008 ? array_update_73205 : array_update_73194[8];
  assign array_update_73207[9] = literal_72009 == 32'h0000_0009 ? array_update_73205 : array_update_73194[9];
  assign array_index_73209 = array_update_72021[add_73206 > 32'h0000_0009 ? 4'h9 : add_73206[3:0]];
  assign array_index_73210 = array_update_73207[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_73214 = smul32b_32b_x_32b(array_index_72024[add_73206 > 32'h0000_0009 ? 4'h9 : add_73206[3:0]], array_index_73209[add_73100 > 32'h0000_0009 ? 4'h9 : add_73100[3:0]]);
  assign add_73216 = array_index_73210[add_73100 > 32'h0000_0009 ? 4'h9 : add_73100[3:0]] + smul_73214;
  assign array_update_73218[0] = add_73100 == 32'h0000_0000 ? add_73216 : array_index_73210[0];
  assign array_update_73218[1] = add_73100 == 32'h0000_0001 ? add_73216 : array_index_73210[1];
  assign array_update_73218[2] = add_73100 == 32'h0000_0002 ? add_73216 : array_index_73210[2];
  assign array_update_73218[3] = add_73100 == 32'h0000_0003 ? add_73216 : array_index_73210[3];
  assign array_update_73218[4] = add_73100 == 32'h0000_0004 ? add_73216 : array_index_73210[4];
  assign array_update_73218[5] = add_73100 == 32'h0000_0005 ? add_73216 : array_index_73210[5];
  assign array_update_73218[6] = add_73100 == 32'h0000_0006 ? add_73216 : array_index_73210[6];
  assign array_update_73218[7] = add_73100 == 32'h0000_0007 ? add_73216 : array_index_73210[7];
  assign array_update_73218[8] = add_73100 == 32'h0000_0008 ? add_73216 : array_index_73210[8];
  assign array_update_73218[9] = add_73100 == 32'h0000_0009 ? add_73216 : array_index_73210[9];
  assign add_73219 = add_73206 + 32'h0000_0001;
  assign array_update_73220[0] = literal_72009 == 32'h0000_0000 ? array_update_73218 : array_update_73207[0];
  assign array_update_73220[1] = literal_72009 == 32'h0000_0001 ? array_update_73218 : array_update_73207[1];
  assign array_update_73220[2] = literal_72009 == 32'h0000_0002 ? array_update_73218 : array_update_73207[2];
  assign array_update_73220[3] = literal_72009 == 32'h0000_0003 ? array_update_73218 : array_update_73207[3];
  assign array_update_73220[4] = literal_72009 == 32'h0000_0004 ? array_update_73218 : array_update_73207[4];
  assign array_update_73220[5] = literal_72009 == 32'h0000_0005 ? array_update_73218 : array_update_73207[5];
  assign array_update_73220[6] = literal_72009 == 32'h0000_0006 ? array_update_73218 : array_update_73207[6];
  assign array_update_73220[7] = literal_72009 == 32'h0000_0007 ? array_update_73218 : array_update_73207[7];
  assign array_update_73220[8] = literal_72009 == 32'h0000_0008 ? array_update_73218 : array_update_73207[8];
  assign array_update_73220[9] = literal_72009 == 32'h0000_0009 ? array_update_73218 : array_update_73207[9];
  assign array_index_73222 = array_update_72021[add_73219 > 32'h0000_0009 ? 4'h9 : add_73219[3:0]];
  assign array_index_73223 = array_update_73220[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_73227 = smul32b_32b_x_32b(array_index_72024[add_73219 > 32'h0000_0009 ? 4'h9 : add_73219[3:0]], array_index_73222[add_73100 > 32'h0000_0009 ? 4'h9 : add_73100[3:0]]);
  assign add_73229 = array_index_73223[add_73100 > 32'h0000_0009 ? 4'h9 : add_73100[3:0]] + smul_73227;
  assign array_update_73230[0] = add_73100 == 32'h0000_0000 ? add_73229 : array_index_73223[0];
  assign array_update_73230[1] = add_73100 == 32'h0000_0001 ? add_73229 : array_index_73223[1];
  assign array_update_73230[2] = add_73100 == 32'h0000_0002 ? add_73229 : array_index_73223[2];
  assign array_update_73230[3] = add_73100 == 32'h0000_0003 ? add_73229 : array_index_73223[3];
  assign array_update_73230[4] = add_73100 == 32'h0000_0004 ? add_73229 : array_index_73223[4];
  assign array_update_73230[5] = add_73100 == 32'h0000_0005 ? add_73229 : array_index_73223[5];
  assign array_update_73230[6] = add_73100 == 32'h0000_0006 ? add_73229 : array_index_73223[6];
  assign array_update_73230[7] = add_73100 == 32'h0000_0007 ? add_73229 : array_index_73223[7];
  assign array_update_73230[8] = add_73100 == 32'h0000_0008 ? add_73229 : array_index_73223[8];
  assign array_update_73230[9] = add_73100 == 32'h0000_0009 ? add_73229 : array_index_73223[9];
  assign array_update_73231[0] = literal_72009 == 32'h0000_0000 ? array_update_73230 : array_update_73220[0];
  assign array_update_73231[1] = literal_72009 == 32'h0000_0001 ? array_update_73230 : array_update_73220[1];
  assign array_update_73231[2] = literal_72009 == 32'h0000_0002 ? array_update_73230 : array_update_73220[2];
  assign array_update_73231[3] = literal_72009 == 32'h0000_0003 ? array_update_73230 : array_update_73220[3];
  assign array_update_73231[4] = literal_72009 == 32'h0000_0004 ? array_update_73230 : array_update_73220[4];
  assign array_update_73231[5] = literal_72009 == 32'h0000_0005 ? array_update_73230 : array_update_73220[5];
  assign array_update_73231[6] = literal_72009 == 32'h0000_0006 ? array_update_73230 : array_update_73220[6];
  assign array_update_73231[7] = literal_72009 == 32'h0000_0007 ? array_update_73230 : array_update_73220[7];
  assign array_update_73231[8] = literal_72009 == 32'h0000_0008 ? array_update_73230 : array_update_73220[8];
  assign array_update_73231[9] = literal_72009 == 32'h0000_0009 ? array_update_73230 : array_update_73220[9];
  assign array_index_73233 = array_update_73231[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign add_73235 = add_73100 + 32'h0000_0001;
  assign array_update_73236[0] = add_73235 == 32'h0000_0000 ? 32'h0000_0000 : array_index_73233[0];
  assign array_update_73236[1] = add_73235 == 32'h0000_0001 ? 32'h0000_0000 : array_index_73233[1];
  assign array_update_73236[2] = add_73235 == 32'h0000_0002 ? 32'h0000_0000 : array_index_73233[2];
  assign array_update_73236[3] = add_73235 == 32'h0000_0003 ? 32'h0000_0000 : array_index_73233[3];
  assign array_update_73236[4] = add_73235 == 32'h0000_0004 ? 32'h0000_0000 : array_index_73233[4];
  assign array_update_73236[5] = add_73235 == 32'h0000_0005 ? 32'h0000_0000 : array_index_73233[5];
  assign array_update_73236[6] = add_73235 == 32'h0000_0006 ? 32'h0000_0000 : array_index_73233[6];
  assign array_update_73236[7] = add_73235 == 32'h0000_0007 ? 32'h0000_0000 : array_index_73233[7];
  assign array_update_73236[8] = add_73235 == 32'h0000_0008 ? 32'h0000_0000 : array_index_73233[8];
  assign array_update_73236[9] = add_73235 == 32'h0000_0009 ? 32'h0000_0000 : array_index_73233[9];
  assign literal_73237 = 32'h0000_0000;
  assign array_update_73238[0] = literal_72009 == 32'h0000_0000 ? array_update_73236 : array_update_73231[0];
  assign array_update_73238[1] = literal_72009 == 32'h0000_0001 ? array_update_73236 : array_update_73231[1];
  assign array_update_73238[2] = literal_72009 == 32'h0000_0002 ? array_update_73236 : array_update_73231[2];
  assign array_update_73238[3] = literal_72009 == 32'h0000_0003 ? array_update_73236 : array_update_73231[3];
  assign array_update_73238[4] = literal_72009 == 32'h0000_0004 ? array_update_73236 : array_update_73231[4];
  assign array_update_73238[5] = literal_72009 == 32'h0000_0005 ? array_update_73236 : array_update_73231[5];
  assign array_update_73238[6] = literal_72009 == 32'h0000_0006 ? array_update_73236 : array_update_73231[6];
  assign array_update_73238[7] = literal_72009 == 32'h0000_0007 ? array_update_73236 : array_update_73231[7];
  assign array_update_73238[8] = literal_72009 == 32'h0000_0008 ? array_update_73236 : array_update_73231[8];
  assign array_update_73238[9] = literal_72009 == 32'h0000_0009 ? array_update_73236 : array_update_73231[9];
  assign array_index_73240 = array_update_72021[literal_73237 > 32'h0000_0009 ? 4'h9 : literal_73237[3:0]];
  assign array_index_73241 = array_update_73238[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_73245 = smul32b_32b_x_32b(array_index_72024[literal_73237 > 32'h0000_0009 ? 4'h9 : literal_73237[3:0]], array_index_73240[add_73235 > 32'h0000_0009 ? 4'h9 : add_73235[3:0]]);
  assign add_73247 = array_index_73241[add_73235 > 32'h0000_0009 ? 4'h9 : add_73235[3:0]] + smul_73245;
  assign array_update_73249[0] = add_73235 == 32'h0000_0000 ? add_73247 : array_index_73241[0];
  assign array_update_73249[1] = add_73235 == 32'h0000_0001 ? add_73247 : array_index_73241[1];
  assign array_update_73249[2] = add_73235 == 32'h0000_0002 ? add_73247 : array_index_73241[2];
  assign array_update_73249[3] = add_73235 == 32'h0000_0003 ? add_73247 : array_index_73241[3];
  assign array_update_73249[4] = add_73235 == 32'h0000_0004 ? add_73247 : array_index_73241[4];
  assign array_update_73249[5] = add_73235 == 32'h0000_0005 ? add_73247 : array_index_73241[5];
  assign array_update_73249[6] = add_73235 == 32'h0000_0006 ? add_73247 : array_index_73241[6];
  assign array_update_73249[7] = add_73235 == 32'h0000_0007 ? add_73247 : array_index_73241[7];
  assign array_update_73249[8] = add_73235 == 32'h0000_0008 ? add_73247 : array_index_73241[8];
  assign array_update_73249[9] = add_73235 == 32'h0000_0009 ? add_73247 : array_index_73241[9];
  assign add_73250 = literal_73237 + 32'h0000_0001;
  assign array_update_73251[0] = literal_72009 == 32'h0000_0000 ? array_update_73249 : array_update_73238[0];
  assign array_update_73251[1] = literal_72009 == 32'h0000_0001 ? array_update_73249 : array_update_73238[1];
  assign array_update_73251[2] = literal_72009 == 32'h0000_0002 ? array_update_73249 : array_update_73238[2];
  assign array_update_73251[3] = literal_72009 == 32'h0000_0003 ? array_update_73249 : array_update_73238[3];
  assign array_update_73251[4] = literal_72009 == 32'h0000_0004 ? array_update_73249 : array_update_73238[4];
  assign array_update_73251[5] = literal_72009 == 32'h0000_0005 ? array_update_73249 : array_update_73238[5];
  assign array_update_73251[6] = literal_72009 == 32'h0000_0006 ? array_update_73249 : array_update_73238[6];
  assign array_update_73251[7] = literal_72009 == 32'h0000_0007 ? array_update_73249 : array_update_73238[7];
  assign array_update_73251[8] = literal_72009 == 32'h0000_0008 ? array_update_73249 : array_update_73238[8];
  assign array_update_73251[9] = literal_72009 == 32'h0000_0009 ? array_update_73249 : array_update_73238[9];
  assign array_index_73253 = array_update_72021[add_73250 > 32'h0000_0009 ? 4'h9 : add_73250[3:0]];
  assign array_index_73254 = array_update_73251[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_73258 = smul32b_32b_x_32b(array_index_72024[add_73250 > 32'h0000_0009 ? 4'h9 : add_73250[3:0]], array_index_73253[add_73235 > 32'h0000_0009 ? 4'h9 : add_73235[3:0]]);
  assign add_73260 = array_index_73254[add_73235 > 32'h0000_0009 ? 4'h9 : add_73235[3:0]] + smul_73258;
  assign array_update_73262[0] = add_73235 == 32'h0000_0000 ? add_73260 : array_index_73254[0];
  assign array_update_73262[1] = add_73235 == 32'h0000_0001 ? add_73260 : array_index_73254[1];
  assign array_update_73262[2] = add_73235 == 32'h0000_0002 ? add_73260 : array_index_73254[2];
  assign array_update_73262[3] = add_73235 == 32'h0000_0003 ? add_73260 : array_index_73254[3];
  assign array_update_73262[4] = add_73235 == 32'h0000_0004 ? add_73260 : array_index_73254[4];
  assign array_update_73262[5] = add_73235 == 32'h0000_0005 ? add_73260 : array_index_73254[5];
  assign array_update_73262[6] = add_73235 == 32'h0000_0006 ? add_73260 : array_index_73254[6];
  assign array_update_73262[7] = add_73235 == 32'h0000_0007 ? add_73260 : array_index_73254[7];
  assign array_update_73262[8] = add_73235 == 32'h0000_0008 ? add_73260 : array_index_73254[8];
  assign array_update_73262[9] = add_73235 == 32'h0000_0009 ? add_73260 : array_index_73254[9];
  assign add_73263 = add_73250 + 32'h0000_0001;
  assign array_update_73264[0] = literal_72009 == 32'h0000_0000 ? array_update_73262 : array_update_73251[0];
  assign array_update_73264[1] = literal_72009 == 32'h0000_0001 ? array_update_73262 : array_update_73251[1];
  assign array_update_73264[2] = literal_72009 == 32'h0000_0002 ? array_update_73262 : array_update_73251[2];
  assign array_update_73264[3] = literal_72009 == 32'h0000_0003 ? array_update_73262 : array_update_73251[3];
  assign array_update_73264[4] = literal_72009 == 32'h0000_0004 ? array_update_73262 : array_update_73251[4];
  assign array_update_73264[5] = literal_72009 == 32'h0000_0005 ? array_update_73262 : array_update_73251[5];
  assign array_update_73264[6] = literal_72009 == 32'h0000_0006 ? array_update_73262 : array_update_73251[6];
  assign array_update_73264[7] = literal_72009 == 32'h0000_0007 ? array_update_73262 : array_update_73251[7];
  assign array_update_73264[8] = literal_72009 == 32'h0000_0008 ? array_update_73262 : array_update_73251[8];
  assign array_update_73264[9] = literal_72009 == 32'h0000_0009 ? array_update_73262 : array_update_73251[9];
  assign array_index_73266 = array_update_72021[add_73263 > 32'h0000_0009 ? 4'h9 : add_73263[3:0]];
  assign array_index_73267 = array_update_73264[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_73271 = smul32b_32b_x_32b(array_index_72024[add_73263 > 32'h0000_0009 ? 4'h9 : add_73263[3:0]], array_index_73266[add_73235 > 32'h0000_0009 ? 4'h9 : add_73235[3:0]]);
  assign add_73273 = array_index_73267[add_73235 > 32'h0000_0009 ? 4'h9 : add_73235[3:0]] + smul_73271;
  assign array_update_73275[0] = add_73235 == 32'h0000_0000 ? add_73273 : array_index_73267[0];
  assign array_update_73275[1] = add_73235 == 32'h0000_0001 ? add_73273 : array_index_73267[1];
  assign array_update_73275[2] = add_73235 == 32'h0000_0002 ? add_73273 : array_index_73267[2];
  assign array_update_73275[3] = add_73235 == 32'h0000_0003 ? add_73273 : array_index_73267[3];
  assign array_update_73275[4] = add_73235 == 32'h0000_0004 ? add_73273 : array_index_73267[4];
  assign array_update_73275[5] = add_73235 == 32'h0000_0005 ? add_73273 : array_index_73267[5];
  assign array_update_73275[6] = add_73235 == 32'h0000_0006 ? add_73273 : array_index_73267[6];
  assign array_update_73275[7] = add_73235 == 32'h0000_0007 ? add_73273 : array_index_73267[7];
  assign array_update_73275[8] = add_73235 == 32'h0000_0008 ? add_73273 : array_index_73267[8];
  assign array_update_73275[9] = add_73235 == 32'h0000_0009 ? add_73273 : array_index_73267[9];
  assign add_73276 = add_73263 + 32'h0000_0001;
  assign array_update_73277[0] = literal_72009 == 32'h0000_0000 ? array_update_73275 : array_update_73264[0];
  assign array_update_73277[1] = literal_72009 == 32'h0000_0001 ? array_update_73275 : array_update_73264[1];
  assign array_update_73277[2] = literal_72009 == 32'h0000_0002 ? array_update_73275 : array_update_73264[2];
  assign array_update_73277[3] = literal_72009 == 32'h0000_0003 ? array_update_73275 : array_update_73264[3];
  assign array_update_73277[4] = literal_72009 == 32'h0000_0004 ? array_update_73275 : array_update_73264[4];
  assign array_update_73277[5] = literal_72009 == 32'h0000_0005 ? array_update_73275 : array_update_73264[5];
  assign array_update_73277[6] = literal_72009 == 32'h0000_0006 ? array_update_73275 : array_update_73264[6];
  assign array_update_73277[7] = literal_72009 == 32'h0000_0007 ? array_update_73275 : array_update_73264[7];
  assign array_update_73277[8] = literal_72009 == 32'h0000_0008 ? array_update_73275 : array_update_73264[8];
  assign array_update_73277[9] = literal_72009 == 32'h0000_0009 ? array_update_73275 : array_update_73264[9];
  assign array_index_73279 = array_update_72021[add_73276 > 32'h0000_0009 ? 4'h9 : add_73276[3:0]];
  assign array_index_73280 = array_update_73277[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_73284 = smul32b_32b_x_32b(array_index_72024[add_73276 > 32'h0000_0009 ? 4'h9 : add_73276[3:0]], array_index_73279[add_73235 > 32'h0000_0009 ? 4'h9 : add_73235[3:0]]);
  assign add_73286 = array_index_73280[add_73235 > 32'h0000_0009 ? 4'h9 : add_73235[3:0]] + smul_73284;
  assign array_update_73288[0] = add_73235 == 32'h0000_0000 ? add_73286 : array_index_73280[0];
  assign array_update_73288[1] = add_73235 == 32'h0000_0001 ? add_73286 : array_index_73280[1];
  assign array_update_73288[2] = add_73235 == 32'h0000_0002 ? add_73286 : array_index_73280[2];
  assign array_update_73288[3] = add_73235 == 32'h0000_0003 ? add_73286 : array_index_73280[3];
  assign array_update_73288[4] = add_73235 == 32'h0000_0004 ? add_73286 : array_index_73280[4];
  assign array_update_73288[5] = add_73235 == 32'h0000_0005 ? add_73286 : array_index_73280[5];
  assign array_update_73288[6] = add_73235 == 32'h0000_0006 ? add_73286 : array_index_73280[6];
  assign array_update_73288[7] = add_73235 == 32'h0000_0007 ? add_73286 : array_index_73280[7];
  assign array_update_73288[8] = add_73235 == 32'h0000_0008 ? add_73286 : array_index_73280[8];
  assign array_update_73288[9] = add_73235 == 32'h0000_0009 ? add_73286 : array_index_73280[9];
  assign add_73289 = add_73276 + 32'h0000_0001;
  assign array_update_73290[0] = literal_72009 == 32'h0000_0000 ? array_update_73288 : array_update_73277[0];
  assign array_update_73290[1] = literal_72009 == 32'h0000_0001 ? array_update_73288 : array_update_73277[1];
  assign array_update_73290[2] = literal_72009 == 32'h0000_0002 ? array_update_73288 : array_update_73277[2];
  assign array_update_73290[3] = literal_72009 == 32'h0000_0003 ? array_update_73288 : array_update_73277[3];
  assign array_update_73290[4] = literal_72009 == 32'h0000_0004 ? array_update_73288 : array_update_73277[4];
  assign array_update_73290[5] = literal_72009 == 32'h0000_0005 ? array_update_73288 : array_update_73277[5];
  assign array_update_73290[6] = literal_72009 == 32'h0000_0006 ? array_update_73288 : array_update_73277[6];
  assign array_update_73290[7] = literal_72009 == 32'h0000_0007 ? array_update_73288 : array_update_73277[7];
  assign array_update_73290[8] = literal_72009 == 32'h0000_0008 ? array_update_73288 : array_update_73277[8];
  assign array_update_73290[9] = literal_72009 == 32'h0000_0009 ? array_update_73288 : array_update_73277[9];
  assign array_index_73292 = array_update_72021[add_73289 > 32'h0000_0009 ? 4'h9 : add_73289[3:0]];
  assign array_index_73293 = array_update_73290[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_73297 = smul32b_32b_x_32b(array_index_72024[add_73289 > 32'h0000_0009 ? 4'h9 : add_73289[3:0]], array_index_73292[add_73235 > 32'h0000_0009 ? 4'h9 : add_73235[3:0]]);
  assign add_73299 = array_index_73293[add_73235 > 32'h0000_0009 ? 4'h9 : add_73235[3:0]] + smul_73297;
  assign array_update_73301[0] = add_73235 == 32'h0000_0000 ? add_73299 : array_index_73293[0];
  assign array_update_73301[1] = add_73235 == 32'h0000_0001 ? add_73299 : array_index_73293[1];
  assign array_update_73301[2] = add_73235 == 32'h0000_0002 ? add_73299 : array_index_73293[2];
  assign array_update_73301[3] = add_73235 == 32'h0000_0003 ? add_73299 : array_index_73293[3];
  assign array_update_73301[4] = add_73235 == 32'h0000_0004 ? add_73299 : array_index_73293[4];
  assign array_update_73301[5] = add_73235 == 32'h0000_0005 ? add_73299 : array_index_73293[5];
  assign array_update_73301[6] = add_73235 == 32'h0000_0006 ? add_73299 : array_index_73293[6];
  assign array_update_73301[7] = add_73235 == 32'h0000_0007 ? add_73299 : array_index_73293[7];
  assign array_update_73301[8] = add_73235 == 32'h0000_0008 ? add_73299 : array_index_73293[8];
  assign array_update_73301[9] = add_73235 == 32'h0000_0009 ? add_73299 : array_index_73293[9];
  assign add_73302 = add_73289 + 32'h0000_0001;
  assign array_update_73303[0] = literal_72009 == 32'h0000_0000 ? array_update_73301 : array_update_73290[0];
  assign array_update_73303[1] = literal_72009 == 32'h0000_0001 ? array_update_73301 : array_update_73290[1];
  assign array_update_73303[2] = literal_72009 == 32'h0000_0002 ? array_update_73301 : array_update_73290[2];
  assign array_update_73303[3] = literal_72009 == 32'h0000_0003 ? array_update_73301 : array_update_73290[3];
  assign array_update_73303[4] = literal_72009 == 32'h0000_0004 ? array_update_73301 : array_update_73290[4];
  assign array_update_73303[5] = literal_72009 == 32'h0000_0005 ? array_update_73301 : array_update_73290[5];
  assign array_update_73303[6] = literal_72009 == 32'h0000_0006 ? array_update_73301 : array_update_73290[6];
  assign array_update_73303[7] = literal_72009 == 32'h0000_0007 ? array_update_73301 : array_update_73290[7];
  assign array_update_73303[8] = literal_72009 == 32'h0000_0008 ? array_update_73301 : array_update_73290[8];
  assign array_update_73303[9] = literal_72009 == 32'h0000_0009 ? array_update_73301 : array_update_73290[9];
  assign array_index_73305 = array_update_72021[add_73302 > 32'h0000_0009 ? 4'h9 : add_73302[3:0]];
  assign array_index_73306 = array_update_73303[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_73310 = smul32b_32b_x_32b(array_index_72024[add_73302 > 32'h0000_0009 ? 4'h9 : add_73302[3:0]], array_index_73305[add_73235 > 32'h0000_0009 ? 4'h9 : add_73235[3:0]]);
  assign add_73312 = array_index_73306[add_73235 > 32'h0000_0009 ? 4'h9 : add_73235[3:0]] + smul_73310;
  assign array_update_73314[0] = add_73235 == 32'h0000_0000 ? add_73312 : array_index_73306[0];
  assign array_update_73314[1] = add_73235 == 32'h0000_0001 ? add_73312 : array_index_73306[1];
  assign array_update_73314[2] = add_73235 == 32'h0000_0002 ? add_73312 : array_index_73306[2];
  assign array_update_73314[3] = add_73235 == 32'h0000_0003 ? add_73312 : array_index_73306[3];
  assign array_update_73314[4] = add_73235 == 32'h0000_0004 ? add_73312 : array_index_73306[4];
  assign array_update_73314[5] = add_73235 == 32'h0000_0005 ? add_73312 : array_index_73306[5];
  assign array_update_73314[6] = add_73235 == 32'h0000_0006 ? add_73312 : array_index_73306[6];
  assign array_update_73314[7] = add_73235 == 32'h0000_0007 ? add_73312 : array_index_73306[7];
  assign array_update_73314[8] = add_73235 == 32'h0000_0008 ? add_73312 : array_index_73306[8];
  assign array_update_73314[9] = add_73235 == 32'h0000_0009 ? add_73312 : array_index_73306[9];
  assign add_73315 = add_73302 + 32'h0000_0001;
  assign array_update_73316[0] = literal_72009 == 32'h0000_0000 ? array_update_73314 : array_update_73303[0];
  assign array_update_73316[1] = literal_72009 == 32'h0000_0001 ? array_update_73314 : array_update_73303[1];
  assign array_update_73316[2] = literal_72009 == 32'h0000_0002 ? array_update_73314 : array_update_73303[2];
  assign array_update_73316[3] = literal_72009 == 32'h0000_0003 ? array_update_73314 : array_update_73303[3];
  assign array_update_73316[4] = literal_72009 == 32'h0000_0004 ? array_update_73314 : array_update_73303[4];
  assign array_update_73316[5] = literal_72009 == 32'h0000_0005 ? array_update_73314 : array_update_73303[5];
  assign array_update_73316[6] = literal_72009 == 32'h0000_0006 ? array_update_73314 : array_update_73303[6];
  assign array_update_73316[7] = literal_72009 == 32'h0000_0007 ? array_update_73314 : array_update_73303[7];
  assign array_update_73316[8] = literal_72009 == 32'h0000_0008 ? array_update_73314 : array_update_73303[8];
  assign array_update_73316[9] = literal_72009 == 32'h0000_0009 ? array_update_73314 : array_update_73303[9];
  assign array_index_73318 = array_update_72021[add_73315 > 32'h0000_0009 ? 4'h9 : add_73315[3:0]];
  assign array_index_73319 = array_update_73316[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_73323 = smul32b_32b_x_32b(array_index_72024[add_73315 > 32'h0000_0009 ? 4'h9 : add_73315[3:0]], array_index_73318[add_73235 > 32'h0000_0009 ? 4'h9 : add_73235[3:0]]);
  assign add_73325 = array_index_73319[add_73235 > 32'h0000_0009 ? 4'h9 : add_73235[3:0]] + smul_73323;
  assign array_update_73327[0] = add_73235 == 32'h0000_0000 ? add_73325 : array_index_73319[0];
  assign array_update_73327[1] = add_73235 == 32'h0000_0001 ? add_73325 : array_index_73319[1];
  assign array_update_73327[2] = add_73235 == 32'h0000_0002 ? add_73325 : array_index_73319[2];
  assign array_update_73327[3] = add_73235 == 32'h0000_0003 ? add_73325 : array_index_73319[3];
  assign array_update_73327[4] = add_73235 == 32'h0000_0004 ? add_73325 : array_index_73319[4];
  assign array_update_73327[5] = add_73235 == 32'h0000_0005 ? add_73325 : array_index_73319[5];
  assign array_update_73327[6] = add_73235 == 32'h0000_0006 ? add_73325 : array_index_73319[6];
  assign array_update_73327[7] = add_73235 == 32'h0000_0007 ? add_73325 : array_index_73319[7];
  assign array_update_73327[8] = add_73235 == 32'h0000_0008 ? add_73325 : array_index_73319[8];
  assign array_update_73327[9] = add_73235 == 32'h0000_0009 ? add_73325 : array_index_73319[9];
  assign add_73328 = add_73315 + 32'h0000_0001;
  assign array_update_73329[0] = literal_72009 == 32'h0000_0000 ? array_update_73327 : array_update_73316[0];
  assign array_update_73329[1] = literal_72009 == 32'h0000_0001 ? array_update_73327 : array_update_73316[1];
  assign array_update_73329[2] = literal_72009 == 32'h0000_0002 ? array_update_73327 : array_update_73316[2];
  assign array_update_73329[3] = literal_72009 == 32'h0000_0003 ? array_update_73327 : array_update_73316[3];
  assign array_update_73329[4] = literal_72009 == 32'h0000_0004 ? array_update_73327 : array_update_73316[4];
  assign array_update_73329[5] = literal_72009 == 32'h0000_0005 ? array_update_73327 : array_update_73316[5];
  assign array_update_73329[6] = literal_72009 == 32'h0000_0006 ? array_update_73327 : array_update_73316[6];
  assign array_update_73329[7] = literal_72009 == 32'h0000_0007 ? array_update_73327 : array_update_73316[7];
  assign array_update_73329[8] = literal_72009 == 32'h0000_0008 ? array_update_73327 : array_update_73316[8];
  assign array_update_73329[9] = literal_72009 == 32'h0000_0009 ? array_update_73327 : array_update_73316[9];
  assign array_index_73331 = array_update_72021[add_73328 > 32'h0000_0009 ? 4'h9 : add_73328[3:0]];
  assign array_index_73332 = array_update_73329[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_73336 = smul32b_32b_x_32b(array_index_72024[add_73328 > 32'h0000_0009 ? 4'h9 : add_73328[3:0]], array_index_73331[add_73235 > 32'h0000_0009 ? 4'h9 : add_73235[3:0]]);
  assign add_73338 = array_index_73332[add_73235 > 32'h0000_0009 ? 4'h9 : add_73235[3:0]] + smul_73336;
  assign array_update_73340[0] = add_73235 == 32'h0000_0000 ? add_73338 : array_index_73332[0];
  assign array_update_73340[1] = add_73235 == 32'h0000_0001 ? add_73338 : array_index_73332[1];
  assign array_update_73340[2] = add_73235 == 32'h0000_0002 ? add_73338 : array_index_73332[2];
  assign array_update_73340[3] = add_73235 == 32'h0000_0003 ? add_73338 : array_index_73332[3];
  assign array_update_73340[4] = add_73235 == 32'h0000_0004 ? add_73338 : array_index_73332[4];
  assign array_update_73340[5] = add_73235 == 32'h0000_0005 ? add_73338 : array_index_73332[5];
  assign array_update_73340[6] = add_73235 == 32'h0000_0006 ? add_73338 : array_index_73332[6];
  assign array_update_73340[7] = add_73235 == 32'h0000_0007 ? add_73338 : array_index_73332[7];
  assign array_update_73340[8] = add_73235 == 32'h0000_0008 ? add_73338 : array_index_73332[8];
  assign array_update_73340[9] = add_73235 == 32'h0000_0009 ? add_73338 : array_index_73332[9];
  assign add_73341 = add_73328 + 32'h0000_0001;
  assign array_update_73342[0] = literal_72009 == 32'h0000_0000 ? array_update_73340 : array_update_73329[0];
  assign array_update_73342[1] = literal_72009 == 32'h0000_0001 ? array_update_73340 : array_update_73329[1];
  assign array_update_73342[2] = literal_72009 == 32'h0000_0002 ? array_update_73340 : array_update_73329[2];
  assign array_update_73342[3] = literal_72009 == 32'h0000_0003 ? array_update_73340 : array_update_73329[3];
  assign array_update_73342[4] = literal_72009 == 32'h0000_0004 ? array_update_73340 : array_update_73329[4];
  assign array_update_73342[5] = literal_72009 == 32'h0000_0005 ? array_update_73340 : array_update_73329[5];
  assign array_update_73342[6] = literal_72009 == 32'h0000_0006 ? array_update_73340 : array_update_73329[6];
  assign array_update_73342[7] = literal_72009 == 32'h0000_0007 ? array_update_73340 : array_update_73329[7];
  assign array_update_73342[8] = literal_72009 == 32'h0000_0008 ? array_update_73340 : array_update_73329[8];
  assign array_update_73342[9] = literal_72009 == 32'h0000_0009 ? array_update_73340 : array_update_73329[9];
  assign array_index_73344 = array_update_72021[add_73341 > 32'h0000_0009 ? 4'h9 : add_73341[3:0]];
  assign array_index_73345 = array_update_73342[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_73349 = smul32b_32b_x_32b(array_index_72024[add_73341 > 32'h0000_0009 ? 4'h9 : add_73341[3:0]], array_index_73344[add_73235 > 32'h0000_0009 ? 4'h9 : add_73235[3:0]]);
  assign add_73351 = array_index_73345[add_73235 > 32'h0000_0009 ? 4'h9 : add_73235[3:0]] + smul_73349;
  assign array_update_73353[0] = add_73235 == 32'h0000_0000 ? add_73351 : array_index_73345[0];
  assign array_update_73353[1] = add_73235 == 32'h0000_0001 ? add_73351 : array_index_73345[1];
  assign array_update_73353[2] = add_73235 == 32'h0000_0002 ? add_73351 : array_index_73345[2];
  assign array_update_73353[3] = add_73235 == 32'h0000_0003 ? add_73351 : array_index_73345[3];
  assign array_update_73353[4] = add_73235 == 32'h0000_0004 ? add_73351 : array_index_73345[4];
  assign array_update_73353[5] = add_73235 == 32'h0000_0005 ? add_73351 : array_index_73345[5];
  assign array_update_73353[6] = add_73235 == 32'h0000_0006 ? add_73351 : array_index_73345[6];
  assign array_update_73353[7] = add_73235 == 32'h0000_0007 ? add_73351 : array_index_73345[7];
  assign array_update_73353[8] = add_73235 == 32'h0000_0008 ? add_73351 : array_index_73345[8];
  assign array_update_73353[9] = add_73235 == 32'h0000_0009 ? add_73351 : array_index_73345[9];
  assign add_73354 = add_73341 + 32'h0000_0001;
  assign array_update_73355[0] = literal_72009 == 32'h0000_0000 ? array_update_73353 : array_update_73342[0];
  assign array_update_73355[1] = literal_72009 == 32'h0000_0001 ? array_update_73353 : array_update_73342[1];
  assign array_update_73355[2] = literal_72009 == 32'h0000_0002 ? array_update_73353 : array_update_73342[2];
  assign array_update_73355[3] = literal_72009 == 32'h0000_0003 ? array_update_73353 : array_update_73342[3];
  assign array_update_73355[4] = literal_72009 == 32'h0000_0004 ? array_update_73353 : array_update_73342[4];
  assign array_update_73355[5] = literal_72009 == 32'h0000_0005 ? array_update_73353 : array_update_73342[5];
  assign array_update_73355[6] = literal_72009 == 32'h0000_0006 ? array_update_73353 : array_update_73342[6];
  assign array_update_73355[7] = literal_72009 == 32'h0000_0007 ? array_update_73353 : array_update_73342[7];
  assign array_update_73355[8] = literal_72009 == 32'h0000_0008 ? array_update_73353 : array_update_73342[8];
  assign array_update_73355[9] = literal_72009 == 32'h0000_0009 ? array_update_73353 : array_update_73342[9];
  assign array_index_73357 = array_update_72021[add_73354 > 32'h0000_0009 ? 4'h9 : add_73354[3:0]];
  assign array_index_73358 = array_update_73355[literal_72009 > 32'h0000_0009 ? 4'h9 : literal_72009[3:0]];
  assign smul_73362 = smul32b_32b_x_32b(array_index_72024[add_73354 > 32'h0000_0009 ? 4'h9 : add_73354[3:0]], array_index_73357[add_73235 > 32'h0000_0009 ? 4'h9 : add_73235[3:0]]);
  assign add_73364 = array_index_73358[add_73235 > 32'h0000_0009 ? 4'h9 : add_73235[3:0]] + smul_73362;
  assign array_update_73365[0] = add_73235 == 32'h0000_0000 ? add_73364 : array_index_73358[0];
  assign array_update_73365[1] = add_73235 == 32'h0000_0001 ? add_73364 : array_index_73358[1];
  assign array_update_73365[2] = add_73235 == 32'h0000_0002 ? add_73364 : array_index_73358[2];
  assign array_update_73365[3] = add_73235 == 32'h0000_0003 ? add_73364 : array_index_73358[3];
  assign array_update_73365[4] = add_73235 == 32'h0000_0004 ? add_73364 : array_index_73358[4];
  assign array_update_73365[5] = add_73235 == 32'h0000_0005 ? add_73364 : array_index_73358[5];
  assign array_update_73365[6] = add_73235 == 32'h0000_0006 ? add_73364 : array_index_73358[6];
  assign array_update_73365[7] = add_73235 == 32'h0000_0007 ? add_73364 : array_index_73358[7];
  assign array_update_73365[8] = add_73235 == 32'h0000_0008 ? add_73364 : array_index_73358[8];
  assign array_update_73365[9] = add_73235 == 32'h0000_0009 ? add_73364 : array_index_73358[9];
  assign array_update_73367[0] = literal_72009 == 32'h0000_0000 ? array_update_73365 : array_update_73355[0];
  assign array_update_73367[1] = literal_72009 == 32'h0000_0001 ? array_update_73365 : array_update_73355[1];
  assign array_update_73367[2] = literal_72009 == 32'h0000_0002 ? array_update_73365 : array_update_73355[2];
  assign array_update_73367[3] = literal_72009 == 32'h0000_0003 ? array_update_73365 : array_update_73355[3];
  assign array_update_73367[4] = literal_72009 == 32'h0000_0004 ? array_update_73365 : array_update_73355[4];
  assign array_update_73367[5] = literal_72009 == 32'h0000_0005 ? array_update_73365 : array_update_73355[5];
  assign array_update_73367[6] = literal_72009 == 32'h0000_0006 ? array_update_73365 : array_update_73355[6];
  assign array_update_73367[7] = literal_72009 == 32'h0000_0007 ? array_update_73365 : array_update_73355[7];
  assign array_update_73367[8] = literal_72009 == 32'h0000_0008 ? array_update_73365 : array_update_73355[8];
  assign array_update_73367[9] = literal_72009 == 32'h0000_0009 ? array_update_73365 : array_update_73355[9];
  assign add_73368 = literal_72009 + 32'h0000_0001;
  assign array_index_73369 = array_update_73367[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign literal_73371 = 32'h0000_0000;
  assign array_update_73372[0] = literal_73371 == 32'h0000_0000 ? 32'h0000_0000 : array_index_73369[0];
  assign array_update_73372[1] = literal_73371 == 32'h0000_0001 ? 32'h0000_0000 : array_index_73369[1];
  assign array_update_73372[2] = literal_73371 == 32'h0000_0002 ? 32'h0000_0000 : array_index_73369[2];
  assign array_update_73372[3] = literal_73371 == 32'h0000_0003 ? 32'h0000_0000 : array_index_73369[3];
  assign array_update_73372[4] = literal_73371 == 32'h0000_0004 ? 32'h0000_0000 : array_index_73369[4];
  assign array_update_73372[5] = literal_73371 == 32'h0000_0005 ? 32'h0000_0000 : array_index_73369[5];
  assign array_update_73372[6] = literal_73371 == 32'h0000_0006 ? 32'h0000_0000 : array_index_73369[6];
  assign array_update_73372[7] = literal_73371 == 32'h0000_0007 ? 32'h0000_0000 : array_index_73369[7];
  assign array_update_73372[8] = literal_73371 == 32'h0000_0008 ? 32'h0000_0000 : array_index_73369[8];
  assign array_update_73372[9] = literal_73371 == 32'h0000_0009 ? 32'h0000_0000 : array_index_73369[9];
  assign literal_73373 = 32'h0000_0000;
  assign array_update_73374[0] = add_73368 == 32'h0000_0000 ? array_update_73372 : array_update_73367[0];
  assign array_update_73374[1] = add_73368 == 32'h0000_0001 ? array_update_73372 : array_update_73367[1];
  assign array_update_73374[2] = add_73368 == 32'h0000_0002 ? array_update_73372 : array_update_73367[2];
  assign array_update_73374[3] = add_73368 == 32'h0000_0003 ? array_update_73372 : array_update_73367[3];
  assign array_update_73374[4] = add_73368 == 32'h0000_0004 ? array_update_73372 : array_update_73367[4];
  assign array_update_73374[5] = add_73368 == 32'h0000_0005 ? array_update_73372 : array_update_73367[5];
  assign array_update_73374[6] = add_73368 == 32'h0000_0006 ? array_update_73372 : array_update_73367[6];
  assign array_update_73374[7] = add_73368 == 32'h0000_0007 ? array_update_73372 : array_update_73367[7];
  assign array_update_73374[8] = add_73368 == 32'h0000_0008 ? array_update_73372 : array_update_73367[8];
  assign array_update_73374[9] = add_73368 == 32'h0000_0009 ? array_update_73372 : array_update_73367[9];
  assign array_index_73375 = array_update_72020[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign array_index_73376 = array_update_72021[literal_73373 > 32'h0000_0009 ? 4'h9 : literal_73373[3:0]];
  assign array_index_73377 = array_update_73374[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_73381 = smul32b_32b_x_32b(array_index_73375[literal_73373 > 32'h0000_0009 ? 4'h9 : literal_73373[3:0]], array_index_73376[literal_73371 > 32'h0000_0009 ? 4'h9 : literal_73371[3:0]]);
  assign add_73383 = array_index_73377[literal_73371 > 32'h0000_0009 ? 4'h9 : literal_73371[3:0]] + smul_73381;
  assign array_update_73385[0] = literal_73371 == 32'h0000_0000 ? add_73383 : array_index_73377[0];
  assign array_update_73385[1] = literal_73371 == 32'h0000_0001 ? add_73383 : array_index_73377[1];
  assign array_update_73385[2] = literal_73371 == 32'h0000_0002 ? add_73383 : array_index_73377[2];
  assign array_update_73385[3] = literal_73371 == 32'h0000_0003 ? add_73383 : array_index_73377[3];
  assign array_update_73385[4] = literal_73371 == 32'h0000_0004 ? add_73383 : array_index_73377[4];
  assign array_update_73385[5] = literal_73371 == 32'h0000_0005 ? add_73383 : array_index_73377[5];
  assign array_update_73385[6] = literal_73371 == 32'h0000_0006 ? add_73383 : array_index_73377[6];
  assign array_update_73385[7] = literal_73371 == 32'h0000_0007 ? add_73383 : array_index_73377[7];
  assign array_update_73385[8] = literal_73371 == 32'h0000_0008 ? add_73383 : array_index_73377[8];
  assign array_update_73385[9] = literal_73371 == 32'h0000_0009 ? add_73383 : array_index_73377[9];
  assign add_73386 = literal_73373 + 32'h0000_0001;
  assign array_update_73387[0] = add_73368 == 32'h0000_0000 ? array_update_73385 : array_update_73374[0];
  assign array_update_73387[1] = add_73368 == 32'h0000_0001 ? array_update_73385 : array_update_73374[1];
  assign array_update_73387[2] = add_73368 == 32'h0000_0002 ? array_update_73385 : array_update_73374[2];
  assign array_update_73387[3] = add_73368 == 32'h0000_0003 ? array_update_73385 : array_update_73374[3];
  assign array_update_73387[4] = add_73368 == 32'h0000_0004 ? array_update_73385 : array_update_73374[4];
  assign array_update_73387[5] = add_73368 == 32'h0000_0005 ? array_update_73385 : array_update_73374[5];
  assign array_update_73387[6] = add_73368 == 32'h0000_0006 ? array_update_73385 : array_update_73374[6];
  assign array_update_73387[7] = add_73368 == 32'h0000_0007 ? array_update_73385 : array_update_73374[7];
  assign array_update_73387[8] = add_73368 == 32'h0000_0008 ? array_update_73385 : array_update_73374[8];
  assign array_update_73387[9] = add_73368 == 32'h0000_0009 ? array_update_73385 : array_update_73374[9];
  assign array_index_73389 = array_update_72021[add_73386 > 32'h0000_0009 ? 4'h9 : add_73386[3:0]];
  assign array_index_73390 = array_update_73387[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_73394 = smul32b_32b_x_32b(array_index_73375[add_73386 > 32'h0000_0009 ? 4'h9 : add_73386[3:0]], array_index_73389[literal_73371 > 32'h0000_0009 ? 4'h9 : literal_73371[3:0]]);
  assign add_73396 = array_index_73390[literal_73371 > 32'h0000_0009 ? 4'h9 : literal_73371[3:0]] + smul_73394;
  assign array_update_73398[0] = literal_73371 == 32'h0000_0000 ? add_73396 : array_index_73390[0];
  assign array_update_73398[1] = literal_73371 == 32'h0000_0001 ? add_73396 : array_index_73390[1];
  assign array_update_73398[2] = literal_73371 == 32'h0000_0002 ? add_73396 : array_index_73390[2];
  assign array_update_73398[3] = literal_73371 == 32'h0000_0003 ? add_73396 : array_index_73390[3];
  assign array_update_73398[4] = literal_73371 == 32'h0000_0004 ? add_73396 : array_index_73390[4];
  assign array_update_73398[5] = literal_73371 == 32'h0000_0005 ? add_73396 : array_index_73390[5];
  assign array_update_73398[6] = literal_73371 == 32'h0000_0006 ? add_73396 : array_index_73390[6];
  assign array_update_73398[7] = literal_73371 == 32'h0000_0007 ? add_73396 : array_index_73390[7];
  assign array_update_73398[8] = literal_73371 == 32'h0000_0008 ? add_73396 : array_index_73390[8];
  assign array_update_73398[9] = literal_73371 == 32'h0000_0009 ? add_73396 : array_index_73390[9];
  assign add_73399 = add_73386 + 32'h0000_0001;
  assign array_update_73400[0] = add_73368 == 32'h0000_0000 ? array_update_73398 : array_update_73387[0];
  assign array_update_73400[1] = add_73368 == 32'h0000_0001 ? array_update_73398 : array_update_73387[1];
  assign array_update_73400[2] = add_73368 == 32'h0000_0002 ? array_update_73398 : array_update_73387[2];
  assign array_update_73400[3] = add_73368 == 32'h0000_0003 ? array_update_73398 : array_update_73387[3];
  assign array_update_73400[4] = add_73368 == 32'h0000_0004 ? array_update_73398 : array_update_73387[4];
  assign array_update_73400[5] = add_73368 == 32'h0000_0005 ? array_update_73398 : array_update_73387[5];
  assign array_update_73400[6] = add_73368 == 32'h0000_0006 ? array_update_73398 : array_update_73387[6];
  assign array_update_73400[7] = add_73368 == 32'h0000_0007 ? array_update_73398 : array_update_73387[7];
  assign array_update_73400[8] = add_73368 == 32'h0000_0008 ? array_update_73398 : array_update_73387[8];
  assign array_update_73400[9] = add_73368 == 32'h0000_0009 ? array_update_73398 : array_update_73387[9];
  assign array_index_73402 = array_update_72021[add_73399 > 32'h0000_0009 ? 4'h9 : add_73399[3:0]];
  assign array_index_73403 = array_update_73400[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_73407 = smul32b_32b_x_32b(array_index_73375[add_73399 > 32'h0000_0009 ? 4'h9 : add_73399[3:0]], array_index_73402[literal_73371 > 32'h0000_0009 ? 4'h9 : literal_73371[3:0]]);
  assign add_73409 = array_index_73403[literal_73371 > 32'h0000_0009 ? 4'h9 : literal_73371[3:0]] + smul_73407;
  assign array_update_73411[0] = literal_73371 == 32'h0000_0000 ? add_73409 : array_index_73403[0];
  assign array_update_73411[1] = literal_73371 == 32'h0000_0001 ? add_73409 : array_index_73403[1];
  assign array_update_73411[2] = literal_73371 == 32'h0000_0002 ? add_73409 : array_index_73403[2];
  assign array_update_73411[3] = literal_73371 == 32'h0000_0003 ? add_73409 : array_index_73403[3];
  assign array_update_73411[4] = literal_73371 == 32'h0000_0004 ? add_73409 : array_index_73403[4];
  assign array_update_73411[5] = literal_73371 == 32'h0000_0005 ? add_73409 : array_index_73403[5];
  assign array_update_73411[6] = literal_73371 == 32'h0000_0006 ? add_73409 : array_index_73403[6];
  assign array_update_73411[7] = literal_73371 == 32'h0000_0007 ? add_73409 : array_index_73403[7];
  assign array_update_73411[8] = literal_73371 == 32'h0000_0008 ? add_73409 : array_index_73403[8];
  assign array_update_73411[9] = literal_73371 == 32'h0000_0009 ? add_73409 : array_index_73403[9];
  assign add_73412 = add_73399 + 32'h0000_0001;
  assign array_update_73413[0] = add_73368 == 32'h0000_0000 ? array_update_73411 : array_update_73400[0];
  assign array_update_73413[1] = add_73368 == 32'h0000_0001 ? array_update_73411 : array_update_73400[1];
  assign array_update_73413[2] = add_73368 == 32'h0000_0002 ? array_update_73411 : array_update_73400[2];
  assign array_update_73413[3] = add_73368 == 32'h0000_0003 ? array_update_73411 : array_update_73400[3];
  assign array_update_73413[4] = add_73368 == 32'h0000_0004 ? array_update_73411 : array_update_73400[4];
  assign array_update_73413[5] = add_73368 == 32'h0000_0005 ? array_update_73411 : array_update_73400[5];
  assign array_update_73413[6] = add_73368 == 32'h0000_0006 ? array_update_73411 : array_update_73400[6];
  assign array_update_73413[7] = add_73368 == 32'h0000_0007 ? array_update_73411 : array_update_73400[7];
  assign array_update_73413[8] = add_73368 == 32'h0000_0008 ? array_update_73411 : array_update_73400[8];
  assign array_update_73413[9] = add_73368 == 32'h0000_0009 ? array_update_73411 : array_update_73400[9];
  assign array_index_73415 = array_update_72021[add_73412 > 32'h0000_0009 ? 4'h9 : add_73412[3:0]];
  assign array_index_73416 = array_update_73413[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_73420 = smul32b_32b_x_32b(array_index_73375[add_73412 > 32'h0000_0009 ? 4'h9 : add_73412[3:0]], array_index_73415[literal_73371 > 32'h0000_0009 ? 4'h9 : literal_73371[3:0]]);
  assign add_73422 = array_index_73416[literal_73371 > 32'h0000_0009 ? 4'h9 : literal_73371[3:0]] + smul_73420;
  assign array_update_73424[0] = literal_73371 == 32'h0000_0000 ? add_73422 : array_index_73416[0];
  assign array_update_73424[1] = literal_73371 == 32'h0000_0001 ? add_73422 : array_index_73416[1];
  assign array_update_73424[2] = literal_73371 == 32'h0000_0002 ? add_73422 : array_index_73416[2];
  assign array_update_73424[3] = literal_73371 == 32'h0000_0003 ? add_73422 : array_index_73416[3];
  assign array_update_73424[4] = literal_73371 == 32'h0000_0004 ? add_73422 : array_index_73416[4];
  assign array_update_73424[5] = literal_73371 == 32'h0000_0005 ? add_73422 : array_index_73416[5];
  assign array_update_73424[6] = literal_73371 == 32'h0000_0006 ? add_73422 : array_index_73416[6];
  assign array_update_73424[7] = literal_73371 == 32'h0000_0007 ? add_73422 : array_index_73416[7];
  assign array_update_73424[8] = literal_73371 == 32'h0000_0008 ? add_73422 : array_index_73416[8];
  assign array_update_73424[9] = literal_73371 == 32'h0000_0009 ? add_73422 : array_index_73416[9];
  assign add_73425 = add_73412 + 32'h0000_0001;
  assign array_update_73426[0] = add_73368 == 32'h0000_0000 ? array_update_73424 : array_update_73413[0];
  assign array_update_73426[1] = add_73368 == 32'h0000_0001 ? array_update_73424 : array_update_73413[1];
  assign array_update_73426[2] = add_73368 == 32'h0000_0002 ? array_update_73424 : array_update_73413[2];
  assign array_update_73426[3] = add_73368 == 32'h0000_0003 ? array_update_73424 : array_update_73413[3];
  assign array_update_73426[4] = add_73368 == 32'h0000_0004 ? array_update_73424 : array_update_73413[4];
  assign array_update_73426[5] = add_73368 == 32'h0000_0005 ? array_update_73424 : array_update_73413[5];
  assign array_update_73426[6] = add_73368 == 32'h0000_0006 ? array_update_73424 : array_update_73413[6];
  assign array_update_73426[7] = add_73368 == 32'h0000_0007 ? array_update_73424 : array_update_73413[7];
  assign array_update_73426[8] = add_73368 == 32'h0000_0008 ? array_update_73424 : array_update_73413[8];
  assign array_update_73426[9] = add_73368 == 32'h0000_0009 ? array_update_73424 : array_update_73413[9];
  assign array_index_73428 = array_update_72021[add_73425 > 32'h0000_0009 ? 4'h9 : add_73425[3:0]];
  assign array_index_73429 = array_update_73426[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_73433 = smul32b_32b_x_32b(array_index_73375[add_73425 > 32'h0000_0009 ? 4'h9 : add_73425[3:0]], array_index_73428[literal_73371 > 32'h0000_0009 ? 4'h9 : literal_73371[3:0]]);
  assign add_73435 = array_index_73429[literal_73371 > 32'h0000_0009 ? 4'h9 : literal_73371[3:0]] + smul_73433;
  assign array_update_73437[0] = literal_73371 == 32'h0000_0000 ? add_73435 : array_index_73429[0];
  assign array_update_73437[1] = literal_73371 == 32'h0000_0001 ? add_73435 : array_index_73429[1];
  assign array_update_73437[2] = literal_73371 == 32'h0000_0002 ? add_73435 : array_index_73429[2];
  assign array_update_73437[3] = literal_73371 == 32'h0000_0003 ? add_73435 : array_index_73429[3];
  assign array_update_73437[4] = literal_73371 == 32'h0000_0004 ? add_73435 : array_index_73429[4];
  assign array_update_73437[5] = literal_73371 == 32'h0000_0005 ? add_73435 : array_index_73429[5];
  assign array_update_73437[6] = literal_73371 == 32'h0000_0006 ? add_73435 : array_index_73429[6];
  assign array_update_73437[7] = literal_73371 == 32'h0000_0007 ? add_73435 : array_index_73429[7];
  assign array_update_73437[8] = literal_73371 == 32'h0000_0008 ? add_73435 : array_index_73429[8];
  assign array_update_73437[9] = literal_73371 == 32'h0000_0009 ? add_73435 : array_index_73429[9];
  assign add_73438 = add_73425 + 32'h0000_0001;
  assign array_update_73439[0] = add_73368 == 32'h0000_0000 ? array_update_73437 : array_update_73426[0];
  assign array_update_73439[1] = add_73368 == 32'h0000_0001 ? array_update_73437 : array_update_73426[1];
  assign array_update_73439[2] = add_73368 == 32'h0000_0002 ? array_update_73437 : array_update_73426[2];
  assign array_update_73439[3] = add_73368 == 32'h0000_0003 ? array_update_73437 : array_update_73426[3];
  assign array_update_73439[4] = add_73368 == 32'h0000_0004 ? array_update_73437 : array_update_73426[4];
  assign array_update_73439[5] = add_73368 == 32'h0000_0005 ? array_update_73437 : array_update_73426[5];
  assign array_update_73439[6] = add_73368 == 32'h0000_0006 ? array_update_73437 : array_update_73426[6];
  assign array_update_73439[7] = add_73368 == 32'h0000_0007 ? array_update_73437 : array_update_73426[7];
  assign array_update_73439[8] = add_73368 == 32'h0000_0008 ? array_update_73437 : array_update_73426[8];
  assign array_update_73439[9] = add_73368 == 32'h0000_0009 ? array_update_73437 : array_update_73426[9];
  assign array_index_73441 = array_update_72021[add_73438 > 32'h0000_0009 ? 4'h9 : add_73438[3:0]];
  assign array_index_73442 = array_update_73439[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_73446 = smul32b_32b_x_32b(array_index_73375[add_73438 > 32'h0000_0009 ? 4'h9 : add_73438[3:0]], array_index_73441[literal_73371 > 32'h0000_0009 ? 4'h9 : literal_73371[3:0]]);
  assign add_73448 = array_index_73442[literal_73371 > 32'h0000_0009 ? 4'h9 : literal_73371[3:0]] + smul_73446;
  assign array_update_73450[0] = literal_73371 == 32'h0000_0000 ? add_73448 : array_index_73442[0];
  assign array_update_73450[1] = literal_73371 == 32'h0000_0001 ? add_73448 : array_index_73442[1];
  assign array_update_73450[2] = literal_73371 == 32'h0000_0002 ? add_73448 : array_index_73442[2];
  assign array_update_73450[3] = literal_73371 == 32'h0000_0003 ? add_73448 : array_index_73442[3];
  assign array_update_73450[4] = literal_73371 == 32'h0000_0004 ? add_73448 : array_index_73442[4];
  assign array_update_73450[5] = literal_73371 == 32'h0000_0005 ? add_73448 : array_index_73442[5];
  assign array_update_73450[6] = literal_73371 == 32'h0000_0006 ? add_73448 : array_index_73442[6];
  assign array_update_73450[7] = literal_73371 == 32'h0000_0007 ? add_73448 : array_index_73442[7];
  assign array_update_73450[8] = literal_73371 == 32'h0000_0008 ? add_73448 : array_index_73442[8];
  assign array_update_73450[9] = literal_73371 == 32'h0000_0009 ? add_73448 : array_index_73442[9];
  assign add_73451 = add_73438 + 32'h0000_0001;
  assign array_update_73452[0] = add_73368 == 32'h0000_0000 ? array_update_73450 : array_update_73439[0];
  assign array_update_73452[1] = add_73368 == 32'h0000_0001 ? array_update_73450 : array_update_73439[1];
  assign array_update_73452[2] = add_73368 == 32'h0000_0002 ? array_update_73450 : array_update_73439[2];
  assign array_update_73452[3] = add_73368 == 32'h0000_0003 ? array_update_73450 : array_update_73439[3];
  assign array_update_73452[4] = add_73368 == 32'h0000_0004 ? array_update_73450 : array_update_73439[4];
  assign array_update_73452[5] = add_73368 == 32'h0000_0005 ? array_update_73450 : array_update_73439[5];
  assign array_update_73452[6] = add_73368 == 32'h0000_0006 ? array_update_73450 : array_update_73439[6];
  assign array_update_73452[7] = add_73368 == 32'h0000_0007 ? array_update_73450 : array_update_73439[7];
  assign array_update_73452[8] = add_73368 == 32'h0000_0008 ? array_update_73450 : array_update_73439[8];
  assign array_update_73452[9] = add_73368 == 32'h0000_0009 ? array_update_73450 : array_update_73439[9];
  assign array_index_73454 = array_update_72021[add_73451 > 32'h0000_0009 ? 4'h9 : add_73451[3:0]];
  assign array_index_73455 = array_update_73452[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_73459 = smul32b_32b_x_32b(array_index_73375[add_73451 > 32'h0000_0009 ? 4'h9 : add_73451[3:0]], array_index_73454[literal_73371 > 32'h0000_0009 ? 4'h9 : literal_73371[3:0]]);
  assign add_73461 = array_index_73455[literal_73371 > 32'h0000_0009 ? 4'h9 : literal_73371[3:0]] + smul_73459;
  assign array_update_73463[0] = literal_73371 == 32'h0000_0000 ? add_73461 : array_index_73455[0];
  assign array_update_73463[1] = literal_73371 == 32'h0000_0001 ? add_73461 : array_index_73455[1];
  assign array_update_73463[2] = literal_73371 == 32'h0000_0002 ? add_73461 : array_index_73455[2];
  assign array_update_73463[3] = literal_73371 == 32'h0000_0003 ? add_73461 : array_index_73455[3];
  assign array_update_73463[4] = literal_73371 == 32'h0000_0004 ? add_73461 : array_index_73455[4];
  assign array_update_73463[5] = literal_73371 == 32'h0000_0005 ? add_73461 : array_index_73455[5];
  assign array_update_73463[6] = literal_73371 == 32'h0000_0006 ? add_73461 : array_index_73455[6];
  assign array_update_73463[7] = literal_73371 == 32'h0000_0007 ? add_73461 : array_index_73455[7];
  assign array_update_73463[8] = literal_73371 == 32'h0000_0008 ? add_73461 : array_index_73455[8];
  assign array_update_73463[9] = literal_73371 == 32'h0000_0009 ? add_73461 : array_index_73455[9];
  assign add_73464 = add_73451 + 32'h0000_0001;
  assign array_update_73465[0] = add_73368 == 32'h0000_0000 ? array_update_73463 : array_update_73452[0];
  assign array_update_73465[1] = add_73368 == 32'h0000_0001 ? array_update_73463 : array_update_73452[1];
  assign array_update_73465[2] = add_73368 == 32'h0000_0002 ? array_update_73463 : array_update_73452[2];
  assign array_update_73465[3] = add_73368 == 32'h0000_0003 ? array_update_73463 : array_update_73452[3];
  assign array_update_73465[4] = add_73368 == 32'h0000_0004 ? array_update_73463 : array_update_73452[4];
  assign array_update_73465[5] = add_73368 == 32'h0000_0005 ? array_update_73463 : array_update_73452[5];
  assign array_update_73465[6] = add_73368 == 32'h0000_0006 ? array_update_73463 : array_update_73452[6];
  assign array_update_73465[7] = add_73368 == 32'h0000_0007 ? array_update_73463 : array_update_73452[7];
  assign array_update_73465[8] = add_73368 == 32'h0000_0008 ? array_update_73463 : array_update_73452[8];
  assign array_update_73465[9] = add_73368 == 32'h0000_0009 ? array_update_73463 : array_update_73452[9];
  assign array_index_73467 = array_update_72021[add_73464 > 32'h0000_0009 ? 4'h9 : add_73464[3:0]];
  assign array_index_73468 = array_update_73465[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_73472 = smul32b_32b_x_32b(array_index_73375[add_73464 > 32'h0000_0009 ? 4'h9 : add_73464[3:0]], array_index_73467[literal_73371 > 32'h0000_0009 ? 4'h9 : literal_73371[3:0]]);
  assign add_73474 = array_index_73468[literal_73371 > 32'h0000_0009 ? 4'h9 : literal_73371[3:0]] + smul_73472;
  assign array_update_73476[0] = literal_73371 == 32'h0000_0000 ? add_73474 : array_index_73468[0];
  assign array_update_73476[1] = literal_73371 == 32'h0000_0001 ? add_73474 : array_index_73468[1];
  assign array_update_73476[2] = literal_73371 == 32'h0000_0002 ? add_73474 : array_index_73468[2];
  assign array_update_73476[3] = literal_73371 == 32'h0000_0003 ? add_73474 : array_index_73468[3];
  assign array_update_73476[4] = literal_73371 == 32'h0000_0004 ? add_73474 : array_index_73468[4];
  assign array_update_73476[5] = literal_73371 == 32'h0000_0005 ? add_73474 : array_index_73468[5];
  assign array_update_73476[6] = literal_73371 == 32'h0000_0006 ? add_73474 : array_index_73468[6];
  assign array_update_73476[7] = literal_73371 == 32'h0000_0007 ? add_73474 : array_index_73468[7];
  assign array_update_73476[8] = literal_73371 == 32'h0000_0008 ? add_73474 : array_index_73468[8];
  assign array_update_73476[9] = literal_73371 == 32'h0000_0009 ? add_73474 : array_index_73468[9];
  assign add_73477 = add_73464 + 32'h0000_0001;
  assign array_update_73478[0] = add_73368 == 32'h0000_0000 ? array_update_73476 : array_update_73465[0];
  assign array_update_73478[1] = add_73368 == 32'h0000_0001 ? array_update_73476 : array_update_73465[1];
  assign array_update_73478[2] = add_73368 == 32'h0000_0002 ? array_update_73476 : array_update_73465[2];
  assign array_update_73478[3] = add_73368 == 32'h0000_0003 ? array_update_73476 : array_update_73465[3];
  assign array_update_73478[4] = add_73368 == 32'h0000_0004 ? array_update_73476 : array_update_73465[4];
  assign array_update_73478[5] = add_73368 == 32'h0000_0005 ? array_update_73476 : array_update_73465[5];
  assign array_update_73478[6] = add_73368 == 32'h0000_0006 ? array_update_73476 : array_update_73465[6];
  assign array_update_73478[7] = add_73368 == 32'h0000_0007 ? array_update_73476 : array_update_73465[7];
  assign array_update_73478[8] = add_73368 == 32'h0000_0008 ? array_update_73476 : array_update_73465[8];
  assign array_update_73478[9] = add_73368 == 32'h0000_0009 ? array_update_73476 : array_update_73465[9];
  assign array_index_73480 = array_update_72021[add_73477 > 32'h0000_0009 ? 4'h9 : add_73477[3:0]];
  assign array_index_73481 = array_update_73478[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_73485 = smul32b_32b_x_32b(array_index_73375[add_73477 > 32'h0000_0009 ? 4'h9 : add_73477[3:0]], array_index_73480[literal_73371 > 32'h0000_0009 ? 4'h9 : literal_73371[3:0]]);
  assign add_73487 = array_index_73481[literal_73371 > 32'h0000_0009 ? 4'h9 : literal_73371[3:0]] + smul_73485;
  assign array_update_73489[0] = literal_73371 == 32'h0000_0000 ? add_73487 : array_index_73481[0];
  assign array_update_73489[1] = literal_73371 == 32'h0000_0001 ? add_73487 : array_index_73481[1];
  assign array_update_73489[2] = literal_73371 == 32'h0000_0002 ? add_73487 : array_index_73481[2];
  assign array_update_73489[3] = literal_73371 == 32'h0000_0003 ? add_73487 : array_index_73481[3];
  assign array_update_73489[4] = literal_73371 == 32'h0000_0004 ? add_73487 : array_index_73481[4];
  assign array_update_73489[5] = literal_73371 == 32'h0000_0005 ? add_73487 : array_index_73481[5];
  assign array_update_73489[6] = literal_73371 == 32'h0000_0006 ? add_73487 : array_index_73481[6];
  assign array_update_73489[7] = literal_73371 == 32'h0000_0007 ? add_73487 : array_index_73481[7];
  assign array_update_73489[8] = literal_73371 == 32'h0000_0008 ? add_73487 : array_index_73481[8];
  assign array_update_73489[9] = literal_73371 == 32'h0000_0009 ? add_73487 : array_index_73481[9];
  assign add_73490 = add_73477 + 32'h0000_0001;
  assign array_update_73491[0] = add_73368 == 32'h0000_0000 ? array_update_73489 : array_update_73478[0];
  assign array_update_73491[1] = add_73368 == 32'h0000_0001 ? array_update_73489 : array_update_73478[1];
  assign array_update_73491[2] = add_73368 == 32'h0000_0002 ? array_update_73489 : array_update_73478[2];
  assign array_update_73491[3] = add_73368 == 32'h0000_0003 ? array_update_73489 : array_update_73478[3];
  assign array_update_73491[4] = add_73368 == 32'h0000_0004 ? array_update_73489 : array_update_73478[4];
  assign array_update_73491[5] = add_73368 == 32'h0000_0005 ? array_update_73489 : array_update_73478[5];
  assign array_update_73491[6] = add_73368 == 32'h0000_0006 ? array_update_73489 : array_update_73478[6];
  assign array_update_73491[7] = add_73368 == 32'h0000_0007 ? array_update_73489 : array_update_73478[7];
  assign array_update_73491[8] = add_73368 == 32'h0000_0008 ? array_update_73489 : array_update_73478[8];
  assign array_update_73491[9] = add_73368 == 32'h0000_0009 ? array_update_73489 : array_update_73478[9];
  assign array_index_73493 = array_update_72021[add_73490 > 32'h0000_0009 ? 4'h9 : add_73490[3:0]];
  assign array_index_73494 = array_update_73491[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_73498 = smul32b_32b_x_32b(array_index_73375[add_73490 > 32'h0000_0009 ? 4'h9 : add_73490[3:0]], array_index_73493[literal_73371 > 32'h0000_0009 ? 4'h9 : literal_73371[3:0]]);
  assign add_73500 = array_index_73494[literal_73371 > 32'h0000_0009 ? 4'h9 : literal_73371[3:0]] + smul_73498;
  assign array_update_73501[0] = literal_73371 == 32'h0000_0000 ? add_73500 : array_index_73494[0];
  assign array_update_73501[1] = literal_73371 == 32'h0000_0001 ? add_73500 : array_index_73494[1];
  assign array_update_73501[2] = literal_73371 == 32'h0000_0002 ? add_73500 : array_index_73494[2];
  assign array_update_73501[3] = literal_73371 == 32'h0000_0003 ? add_73500 : array_index_73494[3];
  assign array_update_73501[4] = literal_73371 == 32'h0000_0004 ? add_73500 : array_index_73494[4];
  assign array_update_73501[5] = literal_73371 == 32'h0000_0005 ? add_73500 : array_index_73494[5];
  assign array_update_73501[6] = literal_73371 == 32'h0000_0006 ? add_73500 : array_index_73494[6];
  assign array_update_73501[7] = literal_73371 == 32'h0000_0007 ? add_73500 : array_index_73494[7];
  assign array_update_73501[8] = literal_73371 == 32'h0000_0008 ? add_73500 : array_index_73494[8];
  assign array_update_73501[9] = literal_73371 == 32'h0000_0009 ? add_73500 : array_index_73494[9];
  assign array_update_73502[0] = add_73368 == 32'h0000_0000 ? array_update_73501 : array_update_73491[0];
  assign array_update_73502[1] = add_73368 == 32'h0000_0001 ? array_update_73501 : array_update_73491[1];
  assign array_update_73502[2] = add_73368 == 32'h0000_0002 ? array_update_73501 : array_update_73491[2];
  assign array_update_73502[3] = add_73368 == 32'h0000_0003 ? array_update_73501 : array_update_73491[3];
  assign array_update_73502[4] = add_73368 == 32'h0000_0004 ? array_update_73501 : array_update_73491[4];
  assign array_update_73502[5] = add_73368 == 32'h0000_0005 ? array_update_73501 : array_update_73491[5];
  assign array_update_73502[6] = add_73368 == 32'h0000_0006 ? array_update_73501 : array_update_73491[6];
  assign array_update_73502[7] = add_73368 == 32'h0000_0007 ? array_update_73501 : array_update_73491[7];
  assign array_update_73502[8] = add_73368 == 32'h0000_0008 ? array_update_73501 : array_update_73491[8];
  assign array_update_73502[9] = add_73368 == 32'h0000_0009 ? array_update_73501 : array_update_73491[9];
  assign array_index_73504 = array_update_73502[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign add_73506 = literal_73371 + 32'h0000_0001;
  assign array_update_73507[0] = add_73506 == 32'h0000_0000 ? 32'h0000_0000 : array_index_73504[0];
  assign array_update_73507[1] = add_73506 == 32'h0000_0001 ? 32'h0000_0000 : array_index_73504[1];
  assign array_update_73507[2] = add_73506 == 32'h0000_0002 ? 32'h0000_0000 : array_index_73504[2];
  assign array_update_73507[3] = add_73506 == 32'h0000_0003 ? 32'h0000_0000 : array_index_73504[3];
  assign array_update_73507[4] = add_73506 == 32'h0000_0004 ? 32'h0000_0000 : array_index_73504[4];
  assign array_update_73507[5] = add_73506 == 32'h0000_0005 ? 32'h0000_0000 : array_index_73504[5];
  assign array_update_73507[6] = add_73506 == 32'h0000_0006 ? 32'h0000_0000 : array_index_73504[6];
  assign array_update_73507[7] = add_73506 == 32'h0000_0007 ? 32'h0000_0000 : array_index_73504[7];
  assign array_update_73507[8] = add_73506 == 32'h0000_0008 ? 32'h0000_0000 : array_index_73504[8];
  assign array_update_73507[9] = add_73506 == 32'h0000_0009 ? 32'h0000_0000 : array_index_73504[9];
  assign literal_73508 = 32'h0000_0000;
  assign array_update_73509[0] = add_73368 == 32'h0000_0000 ? array_update_73507 : array_update_73502[0];
  assign array_update_73509[1] = add_73368 == 32'h0000_0001 ? array_update_73507 : array_update_73502[1];
  assign array_update_73509[2] = add_73368 == 32'h0000_0002 ? array_update_73507 : array_update_73502[2];
  assign array_update_73509[3] = add_73368 == 32'h0000_0003 ? array_update_73507 : array_update_73502[3];
  assign array_update_73509[4] = add_73368 == 32'h0000_0004 ? array_update_73507 : array_update_73502[4];
  assign array_update_73509[5] = add_73368 == 32'h0000_0005 ? array_update_73507 : array_update_73502[5];
  assign array_update_73509[6] = add_73368 == 32'h0000_0006 ? array_update_73507 : array_update_73502[6];
  assign array_update_73509[7] = add_73368 == 32'h0000_0007 ? array_update_73507 : array_update_73502[7];
  assign array_update_73509[8] = add_73368 == 32'h0000_0008 ? array_update_73507 : array_update_73502[8];
  assign array_update_73509[9] = add_73368 == 32'h0000_0009 ? array_update_73507 : array_update_73502[9];
  assign array_index_73511 = array_update_72021[literal_73508 > 32'h0000_0009 ? 4'h9 : literal_73508[3:0]];
  assign array_index_73512 = array_update_73509[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_73516 = smul32b_32b_x_32b(array_index_73375[literal_73508 > 32'h0000_0009 ? 4'h9 : literal_73508[3:0]], array_index_73511[add_73506 > 32'h0000_0009 ? 4'h9 : add_73506[3:0]]);
  assign add_73518 = array_index_73512[add_73506 > 32'h0000_0009 ? 4'h9 : add_73506[3:0]] + smul_73516;
  assign array_update_73520[0] = add_73506 == 32'h0000_0000 ? add_73518 : array_index_73512[0];
  assign array_update_73520[1] = add_73506 == 32'h0000_0001 ? add_73518 : array_index_73512[1];
  assign array_update_73520[2] = add_73506 == 32'h0000_0002 ? add_73518 : array_index_73512[2];
  assign array_update_73520[3] = add_73506 == 32'h0000_0003 ? add_73518 : array_index_73512[3];
  assign array_update_73520[4] = add_73506 == 32'h0000_0004 ? add_73518 : array_index_73512[4];
  assign array_update_73520[5] = add_73506 == 32'h0000_0005 ? add_73518 : array_index_73512[5];
  assign array_update_73520[6] = add_73506 == 32'h0000_0006 ? add_73518 : array_index_73512[6];
  assign array_update_73520[7] = add_73506 == 32'h0000_0007 ? add_73518 : array_index_73512[7];
  assign array_update_73520[8] = add_73506 == 32'h0000_0008 ? add_73518 : array_index_73512[8];
  assign array_update_73520[9] = add_73506 == 32'h0000_0009 ? add_73518 : array_index_73512[9];
  assign add_73521 = literal_73508 + 32'h0000_0001;
  assign array_update_73522[0] = add_73368 == 32'h0000_0000 ? array_update_73520 : array_update_73509[0];
  assign array_update_73522[1] = add_73368 == 32'h0000_0001 ? array_update_73520 : array_update_73509[1];
  assign array_update_73522[2] = add_73368 == 32'h0000_0002 ? array_update_73520 : array_update_73509[2];
  assign array_update_73522[3] = add_73368 == 32'h0000_0003 ? array_update_73520 : array_update_73509[3];
  assign array_update_73522[4] = add_73368 == 32'h0000_0004 ? array_update_73520 : array_update_73509[4];
  assign array_update_73522[5] = add_73368 == 32'h0000_0005 ? array_update_73520 : array_update_73509[5];
  assign array_update_73522[6] = add_73368 == 32'h0000_0006 ? array_update_73520 : array_update_73509[6];
  assign array_update_73522[7] = add_73368 == 32'h0000_0007 ? array_update_73520 : array_update_73509[7];
  assign array_update_73522[8] = add_73368 == 32'h0000_0008 ? array_update_73520 : array_update_73509[8];
  assign array_update_73522[9] = add_73368 == 32'h0000_0009 ? array_update_73520 : array_update_73509[9];
  assign array_index_73524 = array_update_72021[add_73521 > 32'h0000_0009 ? 4'h9 : add_73521[3:0]];
  assign array_index_73525 = array_update_73522[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_73529 = smul32b_32b_x_32b(array_index_73375[add_73521 > 32'h0000_0009 ? 4'h9 : add_73521[3:0]], array_index_73524[add_73506 > 32'h0000_0009 ? 4'h9 : add_73506[3:0]]);
  assign add_73531 = array_index_73525[add_73506 > 32'h0000_0009 ? 4'h9 : add_73506[3:0]] + smul_73529;
  assign array_update_73533[0] = add_73506 == 32'h0000_0000 ? add_73531 : array_index_73525[0];
  assign array_update_73533[1] = add_73506 == 32'h0000_0001 ? add_73531 : array_index_73525[1];
  assign array_update_73533[2] = add_73506 == 32'h0000_0002 ? add_73531 : array_index_73525[2];
  assign array_update_73533[3] = add_73506 == 32'h0000_0003 ? add_73531 : array_index_73525[3];
  assign array_update_73533[4] = add_73506 == 32'h0000_0004 ? add_73531 : array_index_73525[4];
  assign array_update_73533[5] = add_73506 == 32'h0000_0005 ? add_73531 : array_index_73525[5];
  assign array_update_73533[6] = add_73506 == 32'h0000_0006 ? add_73531 : array_index_73525[6];
  assign array_update_73533[7] = add_73506 == 32'h0000_0007 ? add_73531 : array_index_73525[7];
  assign array_update_73533[8] = add_73506 == 32'h0000_0008 ? add_73531 : array_index_73525[8];
  assign array_update_73533[9] = add_73506 == 32'h0000_0009 ? add_73531 : array_index_73525[9];
  assign add_73534 = add_73521 + 32'h0000_0001;
  assign array_update_73535[0] = add_73368 == 32'h0000_0000 ? array_update_73533 : array_update_73522[0];
  assign array_update_73535[1] = add_73368 == 32'h0000_0001 ? array_update_73533 : array_update_73522[1];
  assign array_update_73535[2] = add_73368 == 32'h0000_0002 ? array_update_73533 : array_update_73522[2];
  assign array_update_73535[3] = add_73368 == 32'h0000_0003 ? array_update_73533 : array_update_73522[3];
  assign array_update_73535[4] = add_73368 == 32'h0000_0004 ? array_update_73533 : array_update_73522[4];
  assign array_update_73535[5] = add_73368 == 32'h0000_0005 ? array_update_73533 : array_update_73522[5];
  assign array_update_73535[6] = add_73368 == 32'h0000_0006 ? array_update_73533 : array_update_73522[6];
  assign array_update_73535[7] = add_73368 == 32'h0000_0007 ? array_update_73533 : array_update_73522[7];
  assign array_update_73535[8] = add_73368 == 32'h0000_0008 ? array_update_73533 : array_update_73522[8];
  assign array_update_73535[9] = add_73368 == 32'h0000_0009 ? array_update_73533 : array_update_73522[9];
  assign array_index_73537 = array_update_72021[add_73534 > 32'h0000_0009 ? 4'h9 : add_73534[3:0]];
  assign array_index_73538 = array_update_73535[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_73542 = smul32b_32b_x_32b(array_index_73375[add_73534 > 32'h0000_0009 ? 4'h9 : add_73534[3:0]], array_index_73537[add_73506 > 32'h0000_0009 ? 4'h9 : add_73506[3:0]]);
  assign add_73544 = array_index_73538[add_73506 > 32'h0000_0009 ? 4'h9 : add_73506[3:0]] + smul_73542;
  assign array_update_73546[0] = add_73506 == 32'h0000_0000 ? add_73544 : array_index_73538[0];
  assign array_update_73546[1] = add_73506 == 32'h0000_0001 ? add_73544 : array_index_73538[1];
  assign array_update_73546[2] = add_73506 == 32'h0000_0002 ? add_73544 : array_index_73538[2];
  assign array_update_73546[3] = add_73506 == 32'h0000_0003 ? add_73544 : array_index_73538[3];
  assign array_update_73546[4] = add_73506 == 32'h0000_0004 ? add_73544 : array_index_73538[4];
  assign array_update_73546[5] = add_73506 == 32'h0000_0005 ? add_73544 : array_index_73538[5];
  assign array_update_73546[6] = add_73506 == 32'h0000_0006 ? add_73544 : array_index_73538[6];
  assign array_update_73546[7] = add_73506 == 32'h0000_0007 ? add_73544 : array_index_73538[7];
  assign array_update_73546[8] = add_73506 == 32'h0000_0008 ? add_73544 : array_index_73538[8];
  assign array_update_73546[9] = add_73506 == 32'h0000_0009 ? add_73544 : array_index_73538[9];
  assign add_73547 = add_73534 + 32'h0000_0001;
  assign array_update_73548[0] = add_73368 == 32'h0000_0000 ? array_update_73546 : array_update_73535[0];
  assign array_update_73548[1] = add_73368 == 32'h0000_0001 ? array_update_73546 : array_update_73535[1];
  assign array_update_73548[2] = add_73368 == 32'h0000_0002 ? array_update_73546 : array_update_73535[2];
  assign array_update_73548[3] = add_73368 == 32'h0000_0003 ? array_update_73546 : array_update_73535[3];
  assign array_update_73548[4] = add_73368 == 32'h0000_0004 ? array_update_73546 : array_update_73535[4];
  assign array_update_73548[5] = add_73368 == 32'h0000_0005 ? array_update_73546 : array_update_73535[5];
  assign array_update_73548[6] = add_73368 == 32'h0000_0006 ? array_update_73546 : array_update_73535[6];
  assign array_update_73548[7] = add_73368 == 32'h0000_0007 ? array_update_73546 : array_update_73535[7];
  assign array_update_73548[8] = add_73368 == 32'h0000_0008 ? array_update_73546 : array_update_73535[8];
  assign array_update_73548[9] = add_73368 == 32'h0000_0009 ? array_update_73546 : array_update_73535[9];
  assign array_index_73550 = array_update_72021[add_73547 > 32'h0000_0009 ? 4'h9 : add_73547[3:0]];
  assign array_index_73551 = array_update_73548[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_73555 = smul32b_32b_x_32b(array_index_73375[add_73547 > 32'h0000_0009 ? 4'h9 : add_73547[3:0]], array_index_73550[add_73506 > 32'h0000_0009 ? 4'h9 : add_73506[3:0]]);
  assign add_73557 = array_index_73551[add_73506 > 32'h0000_0009 ? 4'h9 : add_73506[3:0]] + smul_73555;
  assign array_update_73559[0] = add_73506 == 32'h0000_0000 ? add_73557 : array_index_73551[0];
  assign array_update_73559[1] = add_73506 == 32'h0000_0001 ? add_73557 : array_index_73551[1];
  assign array_update_73559[2] = add_73506 == 32'h0000_0002 ? add_73557 : array_index_73551[2];
  assign array_update_73559[3] = add_73506 == 32'h0000_0003 ? add_73557 : array_index_73551[3];
  assign array_update_73559[4] = add_73506 == 32'h0000_0004 ? add_73557 : array_index_73551[4];
  assign array_update_73559[5] = add_73506 == 32'h0000_0005 ? add_73557 : array_index_73551[5];
  assign array_update_73559[6] = add_73506 == 32'h0000_0006 ? add_73557 : array_index_73551[6];
  assign array_update_73559[7] = add_73506 == 32'h0000_0007 ? add_73557 : array_index_73551[7];
  assign array_update_73559[8] = add_73506 == 32'h0000_0008 ? add_73557 : array_index_73551[8];
  assign array_update_73559[9] = add_73506 == 32'h0000_0009 ? add_73557 : array_index_73551[9];
  assign add_73560 = add_73547 + 32'h0000_0001;
  assign array_update_73561[0] = add_73368 == 32'h0000_0000 ? array_update_73559 : array_update_73548[0];
  assign array_update_73561[1] = add_73368 == 32'h0000_0001 ? array_update_73559 : array_update_73548[1];
  assign array_update_73561[2] = add_73368 == 32'h0000_0002 ? array_update_73559 : array_update_73548[2];
  assign array_update_73561[3] = add_73368 == 32'h0000_0003 ? array_update_73559 : array_update_73548[3];
  assign array_update_73561[4] = add_73368 == 32'h0000_0004 ? array_update_73559 : array_update_73548[4];
  assign array_update_73561[5] = add_73368 == 32'h0000_0005 ? array_update_73559 : array_update_73548[5];
  assign array_update_73561[6] = add_73368 == 32'h0000_0006 ? array_update_73559 : array_update_73548[6];
  assign array_update_73561[7] = add_73368 == 32'h0000_0007 ? array_update_73559 : array_update_73548[7];
  assign array_update_73561[8] = add_73368 == 32'h0000_0008 ? array_update_73559 : array_update_73548[8];
  assign array_update_73561[9] = add_73368 == 32'h0000_0009 ? array_update_73559 : array_update_73548[9];
  assign array_index_73563 = array_update_72021[add_73560 > 32'h0000_0009 ? 4'h9 : add_73560[3:0]];
  assign array_index_73564 = array_update_73561[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_73568 = smul32b_32b_x_32b(array_index_73375[add_73560 > 32'h0000_0009 ? 4'h9 : add_73560[3:0]], array_index_73563[add_73506 > 32'h0000_0009 ? 4'h9 : add_73506[3:0]]);
  assign add_73570 = array_index_73564[add_73506 > 32'h0000_0009 ? 4'h9 : add_73506[3:0]] + smul_73568;
  assign array_update_73572[0] = add_73506 == 32'h0000_0000 ? add_73570 : array_index_73564[0];
  assign array_update_73572[1] = add_73506 == 32'h0000_0001 ? add_73570 : array_index_73564[1];
  assign array_update_73572[2] = add_73506 == 32'h0000_0002 ? add_73570 : array_index_73564[2];
  assign array_update_73572[3] = add_73506 == 32'h0000_0003 ? add_73570 : array_index_73564[3];
  assign array_update_73572[4] = add_73506 == 32'h0000_0004 ? add_73570 : array_index_73564[4];
  assign array_update_73572[5] = add_73506 == 32'h0000_0005 ? add_73570 : array_index_73564[5];
  assign array_update_73572[6] = add_73506 == 32'h0000_0006 ? add_73570 : array_index_73564[6];
  assign array_update_73572[7] = add_73506 == 32'h0000_0007 ? add_73570 : array_index_73564[7];
  assign array_update_73572[8] = add_73506 == 32'h0000_0008 ? add_73570 : array_index_73564[8];
  assign array_update_73572[9] = add_73506 == 32'h0000_0009 ? add_73570 : array_index_73564[9];
  assign add_73573 = add_73560 + 32'h0000_0001;
  assign array_update_73574[0] = add_73368 == 32'h0000_0000 ? array_update_73572 : array_update_73561[0];
  assign array_update_73574[1] = add_73368 == 32'h0000_0001 ? array_update_73572 : array_update_73561[1];
  assign array_update_73574[2] = add_73368 == 32'h0000_0002 ? array_update_73572 : array_update_73561[2];
  assign array_update_73574[3] = add_73368 == 32'h0000_0003 ? array_update_73572 : array_update_73561[3];
  assign array_update_73574[4] = add_73368 == 32'h0000_0004 ? array_update_73572 : array_update_73561[4];
  assign array_update_73574[5] = add_73368 == 32'h0000_0005 ? array_update_73572 : array_update_73561[5];
  assign array_update_73574[6] = add_73368 == 32'h0000_0006 ? array_update_73572 : array_update_73561[6];
  assign array_update_73574[7] = add_73368 == 32'h0000_0007 ? array_update_73572 : array_update_73561[7];
  assign array_update_73574[8] = add_73368 == 32'h0000_0008 ? array_update_73572 : array_update_73561[8];
  assign array_update_73574[9] = add_73368 == 32'h0000_0009 ? array_update_73572 : array_update_73561[9];
  assign array_index_73576 = array_update_72021[add_73573 > 32'h0000_0009 ? 4'h9 : add_73573[3:0]];
  assign array_index_73577 = array_update_73574[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_73581 = smul32b_32b_x_32b(array_index_73375[add_73573 > 32'h0000_0009 ? 4'h9 : add_73573[3:0]], array_index_73576[add_73506 > 32'h0000_0009 ? 4'h9 : add_73506[3:0]]);
  assign add_73583 = array_index_73577[add_73506 > 32'h0000_0009 ? 4'h9 : add_73506[3:0]] + smul_73581;
  assign array_update_73585[0] = add_73506 == 32'h0000_0000 ? add_73583 : array_index_73577[0];
  assign array_update_73585[1] = add_73506 == 32'h0000_0001 ? add_73583 : array_index_73577[1];
  assign array_update_73585[2] = add_73506 == 32'h0000_0002 ? add_73583 : array_index_73577[2];
  assign array_update_73585[3] = add_73506 == 32'h0000_0003 ? add_73583 : array_index_73577[3];
  assign array_update_73585[4] = add_73506 == 32'h0000_0004 ? add_73583 : array_index_73577[4];
  assign array_update_73585[5] = add_73506 == 32'h0000_0005 ? add_73583 : array_index_73577[5];
  assign array_update_73585[6] = add_73506 == 32'h0000_0006 ? add_73583 : array_index_73577[6];
  assign array_update_73585[7] = add_73506 == 32'h0000_0007 ? add_73583 : array_index_73577[7];
  assign array_update_73585[8] = add_73506 == 32'h0000_0008 ? add_73583 : array_index_73577[8];
  assign array_update_73585[9] = add_73506 == 32'h0000_0009 ? add_73583 : array_index_73577[9];
  assign add_73586 = add_73573 + 32'h0000_0001;
  assign array_update_73587[0] = add_73368 == 32'h0000_0000 ? array_update_73585 : array_update_73574[0];
  assign array_update_73587[1] = add_73368 == 32'h0000_0001 ? array_update_73585 : array_update_73574[1];
  assign array_update_73587[2] = add_73368 == 32'h0000_0002 ? array_update_73585 : array_update_73574[2];
  assign array_update_73587[3] = add_73368 == 32'h0000_0003 ? array_update_73585 : array_update_73574[3];
  assign array_update_73587[4] = add_73368 == 32'h0000_0004 ? array_update_73585 : array_update_73574[4];
  assign array_update_73587[5] = add_73368 == 32'h0000_0005 ? array_update_73585 : array_update_73574[5];
  assign array_update_73587[6] = add_73368 == 32'h0000_0006 ? array_update_73585 : array_update_73574[6];
  assign array_update_73587[7] = add_73368 == 32'h0000_0007 ? array_update_73585 : array_update_73574[7];
  assign array_update_73587[8] = add_73368 == 32'h0000_0008 ? array_update_73585 : array_update_73574[8];
  assign array_update_73587[9] = add_73368 == 32'h0000_0009 ? array_update_73585 : array_update_73574[9];
  assign array_index_73589 = array_update_72021[add_73586 > 32'h0000_0009 ? 4'h9 : add_73586[3:0]];
  assign array_index_73590 = array_update_73587[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_73594 = smul32b_32b_x_32b(array_index_73375[add_73586 > 32'h0000_0009 ? 4'h9 : add_73586[3:0]], array_index_73589[add_73506 > 32'h0000_0009 ? 4'h9 : add_73506[3:0]]);
  assign add_73596 = array_index_73590[add_73506 > 32'h0000_0009 ? 4'h9 : add_73506[3:0]] + smul_73594;
  assign array_update_73598[0] = add_73506 == 32'h0000_0000 ? add_73596 : array_index_73590[0];
  assign array_update_73598[1] = add_73506 == 32'h0000_0001 ? add_73596 : array_index_73590[1];
  assign array_update_73598[2] = add_73506 == 32'h0000_0002 ? add_73596 : array_index_73590[2];
  assign array_update_73598[3] = add_73506 == 32'h0000_0003 ? add_73596 : array_index_73590[3];
  assign array_update_73598[4] = add_73506 == 32'h0000_0004 ? add_73596 : array_index_73590[4];
  assign array_update_73598[5] = add_73506 == 32'h0000_0005 ? add_73596 : array_index_73590[5];
  assign array_update_73598[6] = add_73506 == 32'h0000_0006 ? add_73596 : array_index_73590[6];
  assign array_update_73598[7] = add_73506 == 32'h0000_0007 ? add_73596 : array_index_73590[7];
  assign array_update_73598[8] = add_73506 == 32'h0000_0008 ? add_73596 : array_index_73590[8];
  assign array_update_73598[9] = add_73506 == 32'h0000_0009 ? add_73596 : array_index_73590[9];
  assign add_73599 = add_73586 + 32'h0000_0001;
  assign array_update_73600[0] = add_73368 == 32'h0000_0000 ? array_update_73598 : array_update_73587[0];
  assign array_update_73600[1] = add_73368 == 32'h0000_0001 ? array_update_73598 : array_update_73587[1];
  assign array_update_73600[2] = add_73368 == 32'h0000_0002 ? array_update_73598 : array_update_73587[2];
  assign array_update_73600[3] = add_73368 == 32'h0000_0003 ? array_update_73598 : array_update_73587[3];
  assign array_update_73600[4] = add_73368 == 32'h0000_0004 ? array_update_73598 : array_update_73587[4];
  assign array_update_73600[5] = add_73368 == 32'h0000_0005 ? array_update_73598 : array_update_73587[5];
  assign array_update_73600[6] = add_73368 == 32'h0000_0006 ? array_update_73598 : array_update_73587[6];
  assign array_update_73600[7] = add_73368 == 32'h0000_0007 ? array_update_73598 : array_update_73587[7];
  assign array_update_73600[8] = add_73368 == 32'h0000_0008 ? array_update_73598 : array_update_73587[8];
  assign array_update_73600[9] = add_73368 == 32'h0000_0009 ? array_update_73598 : array_update_73587[9];
  assign array_index_73602 = array_update_72021[add_73599 > 32'h0000_0009 ? 4'h9 : add_73599[3:0]];
  assign array_index_73603 = array_update_73600[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_73607 = smul32b_32b_x_32b(array_index_73375[add_73599 > 32'h0000_0009 ? 4'h9 : add_73599[3:0]], array_index_73602[add_73506 > 32'h0000_0009 ? 4'h9 : add_73506[3:0]]);
  assign add_73609 = array_index_73603[add_73506 > 32'h0000_0009 ? 4'h9 : add_73506[3:0]] + smul_73607;
  assign array_update_73611[0] = add_73506 == 32'h0000_0000 ? add_73609 : array_index_73603[0];
  assign array_update_73611[1] = add_73506 == 32'h0000_0001 ? add_73609 : array_index_73603[1];
  assign array_update_73611[2] = add_73506 == 32'h0000_0002 ? add_73609 : array_index_73603[2];
  assign array_update_73611[3] = add_73506 == 32'h0000_0003 ? add_73609 : array_index_73603[3];
  assign array_update_73611[4] = add_73506 == 32'h0000_0004 ? add_73609 : array_index_73603[4];
  assign array_update_73611[5] = add_73506 == 32'h0000_0005 ? add_73609 : array_index_73603[5];
  assign array_update_73611[6] = add_73506 == 32'h0000_0006 ? add_73609 : array_index_73603[6];
  assign array_update_73611[7] = add_73506 == 32'h0000_0007 ? add_73609 : array_index_73603[7];
  assign array_update_73611[8] = add_73506 == 32'h0000_0008 ? add_73609 : array_index_73603[8];
  assign array_update_73611[9] = add_73506 == 32'h0000_0009 ? add_73609 : array_index_73603[9];
  assign add_73612 = add_73599 + 32'h0000_0001;
  assign array_update_73613[0] = add_73368 == 32'h0000_0000 ? array_update_73611 : array_update_73600[0];
  assign array_update_73613[1] = add_73368 == 32'h0000_0001 ? array_update_73611 : array_update_73600[1];
  assign array_update_73613[2] = add_73368 == 32'h0000_0002 ? array_update_73611 : array_update_73600[2];
  assign array_update_73613[3] = add_73368 == 32'h0000_0003 ? array_update_73611 : array_update_73600[3];
  assign array_update_73613[4] = add_73368 == 32'h0000_0004 ? array_update_73611 : array_update_73600[4];
  assign array_update_73613[5] = add_73368 == 32'h0000_0005 ? array_update_73611 : array_update_73600[5];
  assign array_update_73613[6] = add_73368 == 32'h0000_0006 ? array_update_73611 : array_update_73600[6];
  assign array_update_73613[7] = add_73368 == 32'h0000_0007 ? array_update_73611 : array_update_73600[7];
  assign array_update_73613[8] = add_73368 == 32'h0000_0008 ? array_update_73611 : array_update_73600[8];
  assign array_update_73613[9] = add_73368 == 32'h0000_0009 ? array_update_73611 : array_update_73600[9];
  assign array_index_73615 = array_update_72021[add_73612 > 32'h0000_0009 ? 4'h9 : add_73612[3:0]];
  assign array_index_73616 = array_update_73613[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_73620 = smul32b_32b_x_32b(array_index_73375[add_73612 > 32'h0000_0009 ? 4'h9 : add_73612[3:0]], array_index_73615[add_73506 > 32'h0000_0009 ? 4'h9 : add_73506[3:0]]);
  assign add_73622 = array_index_73616[add_73506 > 32'h0000_0009 ? 4'h9 : add_73506[3:0]] + smul_73620;
  assign array_update_73624[0] = add_73506 == 32'h0000_0000 ? add_73622 : array_index_73616[0];
  assign array_update_73624[1] = add_73506 == 32'h0000_0001 ? add_73622 : array_index_73616[1];
  assign array_update_73624[2] = add_73506 == 32'h0000_0002 ? add_73622 : array_index_73616[2];
  assign array_update_73624[3] = add_73506 == 32'h0000_0003 ? add_73622 : array_index_73616[3];
  assign array_update_73624[4] = add_73506 == 32'h0000_0004 ? add_73622 : array_index_73616[4];
  assign array_update_73624[5] = add_73506 == 32'h0000_0005 ? add_73622 : array_index_73616[5];
  assign array_update_73624[6] = add_73506 == 32'h0000_0006 ? add_73622 : array_index_73616[6];
  assign array_update_73624[7] = add_73506 == 32'h0000_0007 ? add_73622 : array_index_73616[7];
  assign array_update_73624[8] = add_73506 == 32'h0000_0008 ? add_73622 : array_index_73616[8];
  assign array_update_73624[9] = add_73506 == 32'h0000_0009 ? add_73622 : array_index_73616[9];
  assign add_73625 = add_73612 + 32'h0000_0001;
  assign array_update_73626[0] = add_73368 == 32'h0000_0000 ? array_update_73624 : array_update_73613[0];
  assign array_update_73626[1] = add_73368 == 32'h0000_0001 ? array_update_73624 : array_update_73613[1];
  assign array_update_73626[2] = add_73368 == 32'h0000_0002 ? array_update_73624 : array_update_73613[2];
  assign array_update_73626[3] = add_73368 == 32'h0000_0003 ? array_update_73624 : array_update_73613[3];
  assign array_update_73626[4] = add_73368 == 32'h0000_0004 ? array_update_73624 : array_update_73613[4];
  assign array_update_73626[5] = add_73368 == 32'h0000_0005 ? array_update_73624 : array_update_73613[5];
  assign array_update_73626[6] = add_73368 == 32'h0000_0006 ? array_update_73624 : array_update_73613[6];
  assign array_update_73626[7] = add_73368 == 32'h0000_0007 ? array_update_73624 : array_update_73613[7];
  assign array_update_73626[8] = add_73368 == 32'h0000_0008 ? array_update_73624 : array_update_73613[8];
  assign array_update_73626[9] = add_73368 == 32'h0000_0009 ? array_update_73624 : array_update_73613[9];
  assign array_index_73628 = array_update_72021[add_73625 > 32'h0000_0009 ? 4'h9 : add_73625[3:0]];
  assign array_index_73629 = array_update_73626[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_73633 = smul32b_32b_x_32b(array_index_73375[add_73625 > 32'h0000_0009 ? 4'h9 : add_73625[3:0]], array_index_73628[add_73506 > 32'h0000_0009 ? 4'h9 : add_73506[3:0]]);
  assign add_73635 = array_index_73629[add_73506 > 32'h0000_0009 ? 4'h9 : add_73506[3:0]] + smul_73633;
  assign array_update_73636[0] = add_73506 == 32'h0000_0000 ? add_73635 : array_index_73629[0];
  assign array_update_73636[1] = add_73506 == 32'h0000_0001 ? add_73635 : array_index_73629[1];
  assign array_update_73636[2] = add_73506 == 32'h0000_0002 ? add_73635 : array_index_73629[2];
  assign array_update_73636[3] = add_73506 == 32'h0000_0003 ? add_73635 : array_index_73629[3];
  assign array_update_73636[4] = add_73506 == 32'h0000_0004 ? add_73635 : array_index_73629[4];
  assign array_update_73636[5] = add_73506 == 32'h0000_0005 ? add_73635 : array_index_73629[5];
  assign array_update_73636[6] = add_73506 == 32'h0000_0006 ? add_73635 : array_index_73629[6];
  assign array_update_73636[7] = add_73506 == 32'h0000_0007 ? add_73635 : array_index_73629[7];
  assign array_update_73636[8] = add_73506 == 32'h0000_0008 ? add_73635 : array_index_73629[8];
  assign array_update_73636[9] = add_73506 == 32'h0000_0009 ? add_73635 : array_index_73629[9];
  assign array_update_73637[0] = add_73368 == 32'h0000_0000 ? array_update_73636 : array_update_73626[0];
  assign array_update_73637[1] = add_73368 == 32'h0000_0001 ? array_update_73636 : array_update_73626[1];
  assign array_update_73637[2] = add_73368 == 32'h0000_0002 ? array_update_73636 : array_update_73626[2];
  assign array_update_73637[3] = add_73368 == 32'h0000_0003 ? array_update_73636 : array_update_73626[3];
  assign array_update_73637[4] = add_73368 == 32'h0000_0004 ? array_update_73636 : array_update_73626[4];
  assign array_update_73637[5] = add_73368 == 32'h0000_0005 ? array_update_73636 : array_update_73626[5];
  assign array_update_73637[6] = add_73368 == 32'h0000_0006 ? array_update_73636 : array_update_73626[6];
  assign array_update_73637[7] = add_73368 == 32'h0000_0007 ? array_update_73636 : array_update_73626[7];
  assign array_update_73637[8] = add_73368 == 32'h0000_0008 ? array_update_73636 : array_update_73626[8];
  assign array_update_73637[9] = add_73368 == 32'h0000_0009 ? array_update_73636 : array_update_73626[9];
  assign array_index_73639 = array_update_73637[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign add_73641 = add_73506 + 32'h0000_0001;
  assign array_update_73642[0] = add_73641 == 32'h0000_0000 ? 32'h0000_0000 : array_index_73639[0];
  assign array_update_73642[1] = add_73641 == 32'h0000_0001 ? 32'h0000_0000 : array_index_73639[1];
  assign array_update_73642[2] = add_73641 == 32'h0000_0002 ? 32'h0000_0000 : array_index_73639[2];
  assign array_update_73642[3] = add_73641 == 32'h0000_0003 ? 32'h0000_0000 : array_index_73639[3];
  assign array_update_73642[4] = add_73641 == 32'h0000_0004 ? 32'h0000_0000 : array_index_73639[4];
  assign array_update_73642[5] = add_73641 == 32'h0000_0005 ? 32'h0000_0000 : array_index_73639[5];
  assign array_update_73642[6] = add_73641 == 32'h0000_0006 ? 32'h0000_0000 : array_index_73639[6];
  assign array_update_73642[7] = add_73641 == 32'h0000_0007 ? 32'h0000_0000 : array_index_73639[7];
  assign array_update_73642[8] = add_73641 == 32'h0000_0008 ? 32'h0000_0000 : array_index_73639[8];
  assign array_update_73642[9] = add_73641 == 32'h0000_0009 ? 32'h0000_0000 : array_index_73639[9];
  assign literal_73643 = 32'h0000_0000;
  assign array_update_73644[0] = add_73368 == 32'h0000_0000 ? array_update_73642 : array_update_73637[0];
  assign array_update_73644[1] = add_73368 == 32'h0000_0001 ? array_update_73642 : array_update_73637[1];
  assign array_update_73644[2] = add_73368 == 32'h0000_0002 ? array_update_73642 : array_update_73637[2];
  assign array_update_73644[3] = add_73368 == 32'h0000_0003 ? array_update_73642 : array_update_73637[3];
  assign array_update_73644[4] = add_73368 == 32'h0000_0004 ? array_update_73642 : array_update_73637[4];
  assign array_update_73644[5] = add_73368 == 32'h0000_0005 ? array_update_73642 : array_update_73637[5];
  assign array_update_73644[6] = add_73368 == 32'h0000_0006 ? array_update_73642 : array_update_73637[6];
  assign array_update_73644[7] = add_73368 == 32'h0000_0007 ? array_update_73642 : array_update_73637[7];
  assign array_update_73644[8] = add_73368 == 32'h0000_0008 ? array_update_73642 : array_update_73637[8];
  assign array_update_73644[9] = add_73368 == 32'h0000_0009 ? array_update_73642 : array_update_73637[9];
  assign array_index_73646 = array_update_72021[literal_73643 > 32'h0000_0009 ? 4'h9 : literal_73643[3:0]];
  assign array_index_73647 = array_update_73644[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_73651 = smul32b_32b_x_32b(array_index_73375[literal_73643 > 32'h0000_0009 ? 4'h9 : literal_73643[3:0]], array_index_73646[add_73641 > 32'h0000_0009 ? 4'h9 : add_73641[3:0]]);
  assign add_73653 = array_index_73647[add_73641 > 32'h0000_0009 ? 4'h9 : add_73641[3:0]] + smul_73651;
  assign array_update_73655[0] = add_73641 == 32'h0000_0000 ? add_73653 : array_index_73647[0];
  assign array_update_73655[1] = add_73641 == 32'h0000_0001 ? add_73653 : array_index_73647[1];
  assign array_update_73655[2] = add_73641 == 32'h0000_0002 ? add_73653 : array_index_73647[2];
  assign array_update_73655[3] = add_73641 == 32'h0000_0003 ? add_73653 : array_index_73647[3];
  assign array_update_73655[4] = add_73641 == 32'h0000_0004 ? add_73653 : array_index_73647[4];
  assign array_update_73655[5] = add_73641 == 32'h0000_0005 ? add_73653 : array_index_73647[5];
  assign array_update_73655[6] = add_73641 == 32'h0000_0006 ? add_73653 : array_index_73647[6];
  assign array_update_73655[7] = add_73641 == 32'h0000_0007 ? add_73653 : array_index_73647[7];
  assign array_update_73655[8] = add_73641 == 32'h0000_0008 ? add_73653 : array_index_73647[8];
  assign array_update_73655[9] = add_73641 == 32'h0000_0009 ? add_73653 : array_index_73647[9];
  assign add_73656 = literal_73643 + 32'h0000_0001;
  assign array_update_73657[0] = add_73368 == 32'h0000_0000 ? array_update_73655 : array_update_73644[0];
  assign array_update_73657[1] = add_73368 == 32'h0000_0001 ? array_update_73655 : array_update_73644[1];
  assign array_update_73657[2] = add_73368 == 32'h0000_0002 ? array_update_73655 : array_update_73644[2];
  assign array_update_73657[3] = add_73368 == 32'h0000_0003 ? array_update_73655 : array_update_73644[3];
  assign array_update_73657[4] = add_73368 == 32'h0000_0004 ? array_update_73655 : array_update_73644[4];
  assign array_update_73657[5] = add_73368 == 32'h0000_0005 ? array_update_73655 : array_update_73644[5];
  assign array_update_73657[6] = add_73368 == 32'h0000_0006 ? array_update_73655 : array_update_73644[6];
  assign array_update_73657[7] = add_73368 == 32'h0000_0007 ? array_update_73655 : array_update_73644[7];
  assign array_update_73657[8] = add_73368 == 32'h0000_0008 ? array_update_73655 : array_update_73644[8];
  assign array_update_73657[9] = add_73368 == 32'h0000_0009 ? array_update_73655 : array_update_73644[9];
  assign array_index_73659 = array_update_72021[add_73656 > 32'h0000_0009 ? 4'h9 : add_73656[3:0]];
  assign array_index_73660 = array_update_73657[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_73664 = smul32b_32b_x_32b(array_index_73375[add_73656 > 32'h0000_0009 ? 4'h9 : add_73656[3:0]], array_index_73659[add_73641 > 32'h0000_0009 ? 4'h9 : add_73641[3:0]]);
  assign add_73666 = array_index_73660[add_73641 > 32'h0000_0009 ? 4'h9 : add_73641[3:0]] + smul_73664;
  assign array_update_73668[0] = add_73641 == 32'h0000_0000 ? add_73666 : array_index_73660[0];
  assign array_update_73668[1] = add_73641 == 32'h0000_0001 ? add_73666 : array_index_73660[1];
  assign array_update_73668[2] = add_73641 == 32'h0000_0002 ? add_73666 : array_index_73660[2];
  assign array_update_73668[3] = add_73641 == 32'h0000_0003 ? add_73666 : array_index_73660[3];
  assign array_update_73668[4] = add_73641 == 32'h0000_0004 ? add_73666 : array_index_73660[4];
  assign array_update_73668[5] = add_73641 == 32'h0000_0005 ? add_73666 : array_index_73660[5];
  assign array_update_73668[6] = add_73641 == 32'h0000_0006 ? add_73666 : array_index_73660[6];
  assign array_update_73668[7] = add_73641 == 32'h0000_0007 ? add_73666 : array_index_73660[7];
  assign array_update_73668[8] = add_73641 == 32'h0000_0008 ? add_73666 : array_index_73660[8];
  assign array_update_73668[9] = add_73641 == 32'h0000_0009 ? add_73666 : array_index_73660[9];
  assign add_73669 = add_73656 + 32'h0000_0001;
  assign array_update_73670[0] = add_73368 == 32'h0000_0000 ? array_update_73668 : array_update_73657[0];
  assign array_update_73670[1] = add_73368 == 32'h0000_0001 ? array_update_73668 : array_update_73657[1];
  assign array_update_73670[2] = add_73368 == 32'h0000_0002 ? array_update_73668 : array_update_73657[2];
  assign array_update_73670[3] = add_73368 == 32'h0000_0003 ? array_update_73668 : array_update_73657[3];
  assign array_update_73670[4] = add_73368 == 32'h0000_0004 ? array_update_73668 : array_update_73657[4];
  assign array_update_73670[5] = add_73368 == 32'h0000_0005 ? array_update_73668 : array_update_73657[5];
  assign array_update_73670[6] = add_73368 == 32'h0000_0006 ? array_update_73668 : array_update_73657[6];
  assign array_update_73670[7] = add_73368 == 32'h0000_0007 ? array_update_73668 : array_update_73657[7];
  assign array_update_73670[8] = add_73368 == 32'h0000_0008 ? array_update_73668 : array_update_73657[8];
  assign array_update_73670[9] = add_73368 == 32'h0000_0009 ? array_update_73668 : array_update_73657[9];
  assign array_index_73672 = array_update_72021[add_73669 > 32'h0000_0009 ? 4'h9 : add_73669[3:0]];
  assign array_index_73673 = array_update_73670[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_73677 = smul32b_32b_x_32b(array_index_73375[add_73669 > 32'h0000_0009 ? 4'h9 : add_73669[3:0]], array_index_73672[add_73641 > 32'h0000_0009 ? 4'h9 : add_73641[3:0]]);
  assign add_73679 = array_index_73673[add_73641 > 32'h0000_0009 ? 4'h9 : add_73641[3:0]] + smul_73677;
  assign array_update_73681[0] = add_73641 == 32'h0000_0000 ? add_73679 : array_index_73673[0];
  assign array_update_73681[1] = add_73641 == 32'h0000_0001 ? add_73679 : array_index_73673[1];
  assign array_update_73681[2] = add_73641 == 32'h0000_0002 ? add_73679 : array_index_73673[2];
  assign array_update_73681[3] = add_73641 == 32'h0000_0003 ? add_73679 : array_index_73673[3];
  assign array_update_73681[4] = add_73641 == 32'h0000_0004 ? add_73679 : array_index_73673[4];
  assign array_update_73681[5] = add_73641 == 32'h0000_0005 ? add_73679 : array_index_73673[5];
  assign array_update_73681[6] = add_73641 == 32'h0000_0006 ? add_73679 : array_index_73673[6];
  assign array_update_73681[7] = add_73641 == 32'h0000_0007 ? add_73679 : array_index_73673[7];
  assign array_update_73681[8] = add_73641 == 32'h0000_0008 ? add_73679 : array_index_73673[8];
  assign array_update_73681[9] = add_73641 == 32'h0000_0009 ? add_73679 : array_index_73673[9];
  assign add_73682 = add_73669 + 32'h0000_0001;
  assign array_update_73683[0] = add_73368 == 32'h0000_0000 ? array_update_73681 : array_update_73670[0];
  assign array_update_73683[1] = add_73368 == 32'h0000_0001 ? array_update_73681 : array_update_73670[1];
  assign array_update_73683[2] = add_73368 == 32'h0000_0002 ? array_update_73681 : array_update_73670[2];
  assign array_update_73683[3] = add_73368 == 32'h0000_0003 ? array_update_73681 : array_update_73670[3];
  assign array_update_73683[4] = add_73368 == 32'h0000_0004 ? array_update_73681 : array_update_73670[4];
  assign array_update_73683[5] = add_73368 == 32'h0000_0005 ? array_update_73681 : array_update_73670[5];
  assign array_update_73683[6] = add_73368 == 32'h0000_0006 ? array_update_73681 : array_update_73670[6];
  assign array_update_73683[7] = add_73368 == 32'h0000_0007 ? array_update_73681 : array_update_73670[7];
  assign array_update_73683[8] = add_73368 == 32'h0000_0008 ? array_update_73681 : array_update_73670[8];
  assign array_update_73683[9] = add_73368 == 32'h0000_0009 ? array_update_73681 : array_update_73670[9];
  assign array_index_73685 = array_update_72021[add_73682 > 32'h0000_0009 ? 4'h9 : add_73682[3:0]];
  assign array_index_73686 = array_update_73683[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_73690 = smul32b_32b_x_32b(array_index_73375[add_73682 > 32'h0000_0009 ? 4'h9 : add_73682[3:0]], array_index_73685[add_73641 > 32'h0000_0009 ? 4'h9 : add_73641[3:0]]);
  assign add_73692 = array_index_73686[add_73641 > 32'h0000_0009 ? 4'h9 : add_73641[3:0]] + smul_73690;
  assign array_update_73694[0] = add_73641 == 32'h0000_0000 ? add_73692 : array_index_73686[0];
  assign array_update_73694[1] = add_73641 == 32'h0000_0001 ? add_73692 : array_index_73686[1];
  assign array_update_73694[2] = add_73641 == 32'h0000_0002 ? add_73692 : array_index_73686[2];
  assign array_update_73694[3] = add_73641 == 32'h0000_0003 ? add_73692 : array_index_73686[3];
  assign array_update_73694[4] = add_73641 == 32'h0000_0004 ? add_73692 : array_index_73686[4];
  assign array_update_73694[5] = add_73641 == 32'h0000_0005 ? add_73692 : array_index_73686[5];
  assign array_update_73694[6] = add_73641 == 32'h0000_0006 ? add_73692 : array_index_73686[6];
  assign array_update_73694[7] = add_73641 == 32'h0000_0007 ? add_73692 : array_index_73686[7];
  assign array_update_73694[8] = add_73641 == 32'h0000_0008 ? add_73692 : array_index_73686[8];
  assign array_update_73694[9] = add_73641 == 32'h0000_0009 ? add_73692 : array_index_73686[9];
  assign add_73695 = add_73682 + 32'h0000_0001;
  assign array_update_73696[0] = add_73368 == 32'h0000_0000 ? array_update_73694 : array_update_73683[0];
  assign array_update_73696[1] = add_73368 == 32'h0000_0001 ? array_update_73694 : array_update_73683[1];
  assign array_update_73696[2] = add_73368 == 32'h0000_0002 ? array_update_73694 : array_update_73683[2];
  assign array_update_73696[3] = add_73368 == 32'h0000_0003 ? array_update_73694 : array_update_73683[3];
  assign array_update_73696[4] = add_73368 == 32'h0000_0004 ? array_update_73694 : array_update_73683[4];
  assign array_update_73696[5] = add_73368 == 32'h0000_0005 ? array_update_73694 : array_update_73683[5];
  assign array_update_73696[6] = add_73368 == 32'h0000_0006 ? array_update_73694 : array_update_73683[6];
  assign array_update_73696[7] = add_73368 == 32'h0000_0007 ? array_update_73694 : array_update_73683[7];
  assign array_update_73696[8] = add_73368 == 32'h0000_0008 ? array_update_73694 : array_update_73683[8];
  assign array_update_73696[9] = add_73368 == 32'h0000_0009 ? array_update_73694 : array_update_73683[9];
  assign array_index_73698 = array_update_72021[add_73695 > 32'h0000_0009 ? 4'h9 : add_73695[3:0]];
  assign array_index_73699 = array_update_73696[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_73703 = smul32b_32b_x_32b(array_index_73375[add_73695 > 32'h0000_0009 ? 4'h9 : add_73695[3:0]], array_index_73698[add_73641 > 32'h0000_0009 ? 4'h9 : add_73641[3:0]]);
  assign add_73705 = array_index_73699[add_73641 > 32'h0000_0009 ? 4'h9 : add_73641[3:0]] + smul_73703;
  assign array_update_73707[0] = add_73641 == 32'h0000_0000 ? add_73705 : array_index_73699[0];
  assign array_update_73707[1] = add_73641 == 32'h0000_0001 ? add_73705 : array_index_73699[1];
  assign array_update_73707[2] = add_73641 == 32'h0000_0002 ? add_73705 : array_index_73699[2];
  assign array_update_73707[3] = add_73641 == 32'h0000_0003 ? add_73705 : array_index_73699[3];
  assign array_update_73707[4] = add_73641 == 32'h0000_0004 ? add_73705 : array_index_73699[4];
  assign array_update_73707[5] = add_73641 == 32'h0000_0005 ? add_73705 : array_index_73699[5];
  assign array_update_73707[6] = add_73641 == 32'h0000_0006 ? add_73705 : array_index_73699[6];
  assign array_update_73707[7] = add_73641 == 32'h0000_0007 ? add_73705 : array_index_73699[7];
  assign array_update_73707[8] = add_73641 == 32'h0000_0008 ? add_73705 : array_index_73699[8];
  assign array_update_73707[9] = add_73641 == 32'h0000_0009 ? add_73705 : array_index_73699[9];
  assign add_73708 = add_73695 + 32'h0000_0001;
  assign array_update_73709[0] = add_73368 == 32'h0000_0000 ? array_update_73707 : array_update_73696[0];
  assign array_update_73709[1] = add_73368 == 32'h0000_0001 ? array_update_73707 : array_update_73696[1];
  assign array_update_73709[2] = add_73368 == 32'h0000_0002 ? array_update_73707 : array_update_73696[2];
  assign array_update_73709[3] = add_73368 == 32'h0000_0003 ? array_update_73707 : array_update_73696[3];
  assign array_update_73709[4] = add_73368 == 32'h0000_0004 ? array_update_73707 : array_update_73696[4];
  assign array_update_73709[5] = add_73368 == 32'h0000_0005 ? array_update_73707 : array_update_73696[5];
  assign array_update_73709[6] = add_73368 == 32'h0000_0006 ? array_update_73707 : array_update_73696[6];
  assign array_update_73709[7] = add_73368 == 32'h0000_0007 ? array_update_73707 : array_update_73696[7];
  assign array_update_73709[8] = add_73368 == 32'h0000_0008 ? array_update_73707 : array_update_73696[8];
  assign array_update_73709[9] = add_73368 == 32'h0000_0009 ? array_update_73707 : array_update_73696[9];
  assign array_index_73711 = array_update_72021[add_73708 > 32'h0000_0009 ? 4'h9 : add_73708[3:0]];
  assign array_index_73712 = array_update_73709[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_73716 = smul32b_32b_x_32b(array_index_73375[add_73708 > 32'h0000_0009 ? 4'h9 : add_73708[3:0]], array_index_73711[add_73641 > 32'h0000_0009 ? 4'h9 : add_73641[3:0]]);
  assign add_73718 = array_index_73712[add_73641 > 32'h0000_0009 ? 4'h9 : add_73641[3:0]] + smul_73716;
  assign array_update_73720[0] = add_73641 == 32'h0000_0000 ? add_73718 : array_index_73712[0];
  assign array_update_73720[1] = add_73641 == 32'h0000_0001 ? add_73718 : array_index_73712[1];
  assign array_update_73720[2] = add_73641 == 32'h0000_0002 ? add_73718 : array_index_73712[2];
  assign array_update_73720[3] = add_73641 == 32'h0000_0003 ? add_73718 : array_index_73712[3];
  assign array_update_73720[4] = add_73641 == 32'h0000_0004 ? add_73718 : array_index_73712[4];
  assign array_update_73720[5] = add_73641 == 32'h0000_0005 ? add_73718 : array_index_73712[5];
  assign array_update_73720[6] = add_73641 == 32'h0000_0006 ? add_73718 : array_index_73712[6];
  assign array_update_73720[7] = add_73641 == 32'h0000_0007 ? add_73718 : array_index_73712[7];
  assign array_update_73720[8] = add_73641 == 32'h0000_0008 ? add_73718 : array_index_73712[8];
  assign array_update_73720[9] = add_73641 == 32'h0000_0009 ? add_73718 : array_index_73712[9];
  assign add_73721 = add_73708 + 32'h0000_0001;
  assign array_update_73722[0] = add_73368 == 32'h0000_0000 ? array_update_73720 : array_update_73709[0];
  assign array_update_73722[1] = add_73368 == 32'h0000_0001 ? array_update_73720 : array_update_73709[1];
  assign array_update_73722[2] = add_73368 == 32'h0000_0002 ? array_update_73720 : array_update_73709[2];
  assign array_update_73722[3] = add_73368 == 32'h0000_0003 ? array_update_73720 : array_update_73709[3];
  assign array_update_73722[4] = add_73368 == 32'h0000_0004 ? array_update_73720 : array_update_73709[4];
  assign array_update_73722[5] = add_73368 == 32'h0000_0005 ? array_update_73720 : array_update_73709[5];
  assign array_update_73722[6] = add_73368 == 32'h0000_0006 ? array_update_73720 : array_update_73709[6];
  assign array_update_73722[7] = add_73368 == 32'h0000_0007 ? array_update_73720 : array_update_73709[7];
  assign array_update_73722[8] = add_73368 == 32'h0000_0008 ? array_update_73720 : array_update_73709[8];
  assign array_update_73722[9] = add_73368 == 32'h0000_0009 ? array_update_73720 : array_update_73709[9];
  assign array_index_73724 = array_update_72021[add_73721 > 32'h0000_0009 ? 4'h9 : add_73721[3:0]];
  assign array_index_73725 = array_update_73722[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_73729 = smul32b_32b_x_32b(array_index_73375[add_73721 > 32'h0000_0009 ? 4'h9 : add_73721[3:0]], array_index_73724[add_73641 > 32'h0000_0009 ? 4'h9 : add_73641[3:0]]);
  assign add_73731 = array_index_73725[add_73641 > 32'h0000_0009 ? 4'h9 : add_73641[3:0]] + smul_73729;
  assign array_update_73733[0] = add_73641 == 32'h0000_0000 ? add_73731 : array_index_73725[0];
  assign array_update_73733[1] = add_73641 == 32'h0000_0001 ? add_73731 : array_index_73725[1];
  assign array_update_73733[2] = add_73641 == 32'h0000_0002 ? add_73731 : array_index_73725[2];
  assign array_update_73733[3] = add_73641 == 32'h0000_0003 ? add_73731 : array_index_73725[3];
  assign array_update_73733[4] = add_73641 == 32'h0000_0004 ? add_73731 : array_index_73725[4];
  assign array_update_73733[5] = add_73641 == 32'h0000_0005 ? add_73731 : array_index_73725[5];
  assign array_update_73733[6] = add_73641 == 32'h0000_0006 ? add_73731 : array_index_73725[6];
  assign array_update_73733[7] = add_73641 == 32'h0000_0007 ? add_73731 : array_index_73725[7];
  assign array_update_73733[8] = add_73641 == 32'h0000_0008 ? add_73731 : array_index_73725[8];
  assign array_update_73733[9] = add_73641 == 32'h0000_0009 ? add_73731 : array_index_73725[9];
  assign add_73734 = add_73721 + 32'h0000_0001;
  assign array_update_73735[0] = add_73368 == 32'h0000_0000 ? array_update_73733 : array_update_73722[0];
  assign array_update_73735[1] = add_73368 == 32'h0000_0001 ? array_update_73733 : array_update_73722[1];
  assign array_update_73735[2] = add_73368 == 32'h0000_0002 ? array_update_73733 : array_update_73722[2];
  assign array_update_73735[3] = add_73368 == 32'h0000_0003 ? array_update_73733 : array_update_73722[3];
  assign array_update_73735[4] = add_73368 == 32'h0000_0004 ? array_update_73733 : array_update_73722[4];
  assign array_update_73735[5] = add_73368 == 32'h0000_0005 ? array_update_73733 : array_update_73722[5];
  assign array_update_73735[6] = add_73368 == 32'h0000_0006 ? array_update_73733 : array_update_73722[6];
  assign array_update_73735[7] = add_73368 == 32'h0000_0007 ? array_update_73733 : array_update_73722[7];
  assign array_update_73735[8] = add_73368 == 32'h0000_0008 ? array_update_73733 : array_update_73722[8];
  assign array_update_73735[9] = add_73368 == 32'h0000_0009 ? array_update_73733 : array_update_73722[9];
  assign array_index_73737 = array_update_72021[add_73734 > 32'h0000_0009 ? 4'h9 : add_73734[3:0]];
  assign array_index_73738 = array_update_73735[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_73742 = smul32b_32b_x_32b(array_index_73375[add_73734 > 32'h0000_0009 ? 4'h9 : add_73734[3:0]], array_index_73737[add_73641 > 32'h0000_0009 ? 4'h9 : add_73641[3:0]]);
  assign add_73744 = array_index_73738[add_73641 > 32'h0000_0009 ? 4'h9 : add_73641[3:0]] + smul_73742;
  assign array_update_73746[0] = add_73641 == 32'h0000_0000 ? add_73744 : array_index_73738[0];
  assign array_update_73746[1] = add_73641 == 32'h0000_0001 ? add_73744 : array_index_73738[1];
  assign array_update_73746[2] = add_73641 == 32'h0000_0002 ? add_73744 : array_index_73738[2];
  assign array_update_73746[3] = add_73641 == 32'h0000_0003 ? add_73744 : array_index_73738[3];
  assign array_update_73746[4] = add_73641 == 32'h0000_0004 ? add_73744 : array_index_73738[4];
  assign array_update_73746[5] = add_73641 == 32'h0000_0005 ? add_73744 : array_index_73738[5];
  assign array_update_73746[6] = add_73641 == 32'h0000_0006 ? add_73744 : array_index_73738[6];
  assign array_update_73746[7] = add_73641 == 32'h0000_0007 ? add_73744 : array_index_73738[7];
  assign array_update_73746[8] = add_73641 == 32'h0000_0008 ? add_73744 : array_index_73738[8];
  assign array_update_73746[9] = add_73641 == 32'h0000_0009 ? add_73744 : array_index_73738[9];
  assign add_73747 = add_73734 + 32'h0000_0001;
  assign array_update_73748[0] = add_73368 == 32'h0000_0000 ? array_update_73746 : array_update_73735[0];
  assign array_update_73748[1] = add_73368 == 32'h0000_0001 ? array_update_73746 : array_update_73735[1];
  assign array_update_73748[2] = add_73368 == 32'h0000_0002 ? array_update_73746 : array_update_73735[2];
  assign array_update_73748[3] = add_73368 == 32'h0000_0003 ? array_update_73746 : array_update_73735[3];
  assign array_update_73748[4] = add_73368 == 32'h0000_0004 ? array_update_73746 : array_update_73735[4];
  assign array_update_73748[5] = add_73368 == 32'h0000_0005 ? array_update_73746 : array_update_73735[5];
  assign array_update_73748[6] = add_73368 == 32'h0000_0006 ? array_update_73746 : array_update_73735[6];
  assign array_update_73748[7] = add_73368 == 32'h0000_0007 ? array_update_73746 : array_update_73735[7];
  assign array_update_73748[8] = add_73368 == 32'h0000_0008 ? array_update_73746 : array_update_73735[8];
  assign array_update_73748[9] = add_73368 == 32'h0000_0009 ? array_update_73746 : array_update_73735[9];
  assign array_index_73750 = array_update_72021[add_73747 > 32'h0000_0009 ? 4'h9 : add_73747[3:0]];
  assign array_index_73751 = array_update_73748[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_73755 = smul32b_32b_x_32b(array_index_73375[add_73747 > 32'h0000_0009 ? 4'h9 : add_73747[3:0]], array_index_73750[add_73641 > 32'h0000_0009 ? 4'h9 : add_73641[3:0]]);
  assign add_73757 = array_index_73751[add_73641 > 32'h0000_0009 ? 4'h9 : add_73641[3:0]] + smul_73755;
  assign array_update_73759[0] = add_73641 == 32'h0000_0000 ? add_73757 : array_index_73751[0];
  assign array_update_73759[1] = add_73641 == 32'h0000_0001 ? add_73757 : array_index_73751[1];
  assign array_update_73759[2] = add_73641 == 32'h0000_0002 ? add_73757 : array_index_73751[2];
  assign array_update_73759[3] = add_73641 == 32'h0000_0003 ? add_73757 : array_index_73751[3];
  assign array_update_73759[4] = add_73641 == 32'h0000_0004 ? add_73757 : array_index_73751[4];
  assign array_update_73759[5] = add_73641 == 32'h0000_0005 ? add_73757 : array_index_73751[5];
  assign array_update_73759[6] = add_73641 == 32'h0000_0006 ? add_73757 : array_index_73751[6];
  assign array_update_73759[7] = add_73641 == 32'h0000_0007 ? add_73757 : array_index_73751[7];
  assign array_update_73759[8] = add_73641 == 32'h0000_0008 ? add_73757 : array_index_73751[8];
  assign array_update_73759[9] = add_73641 == 32'h0000_0009 ? add_73757 : array_index_73751[9];
  assign add_73760 = add_73747 + 32'h0000_0001;
  assign array_update_73761[0] = add_73368 == 32'h0000_0000 ? array_update_73759 : array_update_73748[0];
  assign array_update_73761[1] = add_73368 == 32'h0000_0001 ? array_update_73759 : array_update_73748[1];
  assign array_update_73761[2] = add_73368 == 32'h0000_0002 ? array_update_73759 : array_update_73748[2];
  assign array_update_73761[3] = add_73368 == 32'h0000_0003 ? array_update_73759 : array_update_73748[3];
  assign array_update_73761[4] = add_73368 == 32'h0000_0004 ? array_update_73759 : array_update_73748[4];
  assign array_update_73761[5] = add_73368 == 32'h0000_0005 ? array_update_73759 : array_update_73748[5];
  assign array_update_73761[6] = add_73368 == 32'h0000_0006 ? array_update_73759 : array_update_73748[6];
  assign array_update_73761[7] = add_73368 == 32'h0000_0007 ? array_update_73759 : array_update_73748[7];
  assign array_update_73761[8] = add_73368 == 32'h0000_0008 ? array_update_73759 : array_update_73748[8];
  assign array_update_73761[9] = add_73368 == 32'h0000_0009 ? array_update_73759 : array_update_73748[9];
  assign array_index_73763 = array_update_72021[add_73760 > 32'h0000_0009 ? 4'h9 : add_73760[3:0]];
  assign array_index_73764 = array_update_73761[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_73768 = smul32b_32b_x_32b(array_index_73375[add_73760 > 32'h0000_0009 ? 4'h9 : add_73760[3:0]], array_index_73763[add_73641 > 32'h0000_0009 ? 4'h9 : add_73641[3:0]]);
  assign add_73770 = array_index_73764[add_73641 > 32'h0000_0009 ? 4'h9 : add_73641[3:0]] + smul_73768;
  assign array_update_73771[0] = add_73641 == 32'h0000_0000 ? add_73770 : array_index_73764[0];
  assign array_update_73771[1] = add_73641 == 32'h0000_0001 ? add_73770 : array_index_73764[1];
  assign array_update_73771[2] = add_73641 == 32'h0000_0002 ? add_73770 : array_index_73764[2];
  assign array_update_73771[3] = add_73641 == 32'h0000_0003 ? add_73770 : array_index_73764[3];
  assign array_update_73771[4] = add_73641 == 32'h0000_0004 ? add_73770 : array_index_73764[4];
  assign array_update_73771[5] = add_73641 == 32'h0000_0005 ? add_73770 : array_index_73764[5];
  assign array_update_73771[6] = add_73641 == 32'h0000_0006 ? add_73770 : array_index_73764[6];
  assign array_update_73771[7] = add_73641 == 32'h0000_0007 ? add_73770 : array_index_73764[7];
  assign array_update_73771[8] = add_73641 == 32'h0000_0008 ? add_73770 : array_index_73764[8];
  assign array_update_73771[9] = add_73641 == 32'h0000_0009 ? add_73770 : array_index_73764[9];
  assign array_update_73772[0] = add_73368 == 32'h0000_0000 ? array_update_73771 : array_update_73761[0];
  assign array_update_73772[1] = add_73368 == 32'h0000_0001 ? array_update_73771 : array_update_73761[1];
  assign array_update_73772[2] = add_73368 == 32'h0000_0002 ? array_update_73771 : array_update_73761[2];
  assign array_update_73772[3] = add_73368 == 32'h0000_0003 ? array_update_73771 : array_update_73761[3];
  assign array_update_73772[4] = add_73368 == 32'h0000_0004 ? array_update_73771 : array_update_73761[4];
  assign array_update_73772[5] = add_73368 == 32'h0000_0005 ? array_update_73771 : array_update_73761[5];
  assign array_update_73772[6] = add_73368 == 32'h0000_0006 ? array_update_73771 : array_update_73761[6];
  assign array_update_73772[7] = add_73368 == 32'h0000_0007 ? array_update_73771 : array_update_73761[7];
  assign array_update_73772[8] = add_73368 == 32'h0000_0008 ? array_update_73771 : array_update_73761[8];
  assign array_update_73772[9] = add_73368 == 32'h0000_0009 ? array_update_73771 : array_update_73761[9];
  assign array_index_73774 = array_update_73772[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign add_73776 = add_73641 + 32'h0000_0001;
  assign array_update_73777[0] = add_73776 == 32'h0000_0000 ? 32'h0000_0000 : array_index_73774[0];
  assign array_update_73777[1] = add_73776 == 32'h0000_0001 ? 32'h0000_0000 : array_index_73774[1];
  assign array_update_73777[2] = add_73776 == 32'h0000_0002 ? 32'h0000_0000 : array_index_73774[2];
  assign array_update_73777[3] = add_73776 == 32'h0000_0003 ? 32'h0000_0000 : array_index_73774[3];
  assign array_update_73777[4] = add_73776 == 32'h0000_0004 ? 32'h0000_0000 : array_index_73774[4];
  assign array_update_73777[5] = add_73776 == 32'h0000_0005 ? 32'h0000_0000 : array_index_73774[5];
  assign array_update_73777[6] = add_73776 == 32'h0000_0006 ? 32'h0000_0000 : array_index_73774[6];
  assign array_update_73777[7] = add_73776 == 32'h0000_0007 ? 32'h0000_0000 : array_index_73774[7];
  assign array_update_73777[8] = add_73776 == 32'h0000_0008 ? 32'h0000_0000 : array_index_73774[8];
  assign array_update_73777[9] = add_73776 == 32'h0000_0009 ? 32'h0000_0000 : array_index_73774[9];
  assign literal_73778 = 32'h0000_0000;
  assign array_update_73779[0] = add_73368 == 32'h0000_0000 ? array_update_73777 : array_update_73772[0];
  assign array_update_73779[1] = add_73368 == 32'h0000_0001 ? array_update_73777 : array_update_73772[1];
  assign array_update_73779[2] = add_73368 == 32'h0000_0002 ? array_update_73777 : array_update_73772[2];
  assign array_update_73779[3] = add_73368 == 32'h0000_0003 ? array_update_73777 : array_update_73772[3];
  assign array_update_73779[4] = add_73368 == 32'h0000_0004 ? array_update_73777 : array_update_73772[4];
  assign array_update_73779[5] = add_73368 == 32'h0000_0005 ? array_update_73777 : array_update_73772[5];
  assign array_update_73779[6] = add_73368 == 32'h0000_0006 ? array_update_73777 : array_update_73772[6];
  assign array_update_73779[7] = add_73368 == 32'h0000_0007 ? array_update_73777 : array_update_73772[7];
  assign array_update_73779[8] = add_73368 == 32'h0000_0008 ? array_update_73777 : array_update_73772[8];
  assign array_update_73779[9] = add_73368 == 32'h0000_0009 ? array_update_73777 : array_update_73772[9];
  assign array_index_73781 = array_update_72021[literal_73778 > 32'h0000_0009 ? 4'h9 : literal_73778[3:0]];
  assign array_index_73782 = array_update_73779[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_73786 = smul32b_32b_x_32b(array_index_73375[literal_73778 > 32'h0000_0009 ? 4'h9 : literal_73778[3:0]], array_index_73781[add_73776 > 32'h0000_0009 ? 4'h9 : add_73776[3:0]]);
  assign add_73788 = array_index_73782[add_73776 > 32'h0000_0009 ? 4'h9 : add_73776[3:0]] + smul_73786;
  assign array_update_73790[0] = add_73776 == 32'h0000_0000 ? add_73788 : array_index_73782[0];
  assign array_update_73790[1] = add_73776 == 32'h0000_0001 ? add_73788 : array_index_73782[1];
  assign array_update_73790[2] = add_73776 == 32'h0000_0002 ? add_73788 : array_index_73782[2];
  assign array_update_73790[3] = add_73776 == 32'h0000_0003 ? add_73788 : array_index_73782[3];
  assign array_update_73790[4] = add_73776 == 32'h0000_0004 ? add_73788 : array_index_73782[4];
  assign array_update_73790[5] = add_73776 == 32'h0000_0005 ? add_73788 : array_index_73782[5];
  assign array_update_73790[6] = add_73776 == 32'h0000_0006 ? add_73788 : array_index_73782[6];
  assign array_update_73790[7] = add_73776 == 32'h0000_0007 ? add_73788 : array_index_73782[7];
  assign array_update_73790[8] = add_73776 == 32'h0000_0008 ? add_73788 : array_index_73782[8];
  assign array_update_73790[9] = add_73776 == 32'h0000_0009 ? add_73788 : array_index_73782[9];
  assign add_73791 = literal_73778 + 32'h0000_0001;
  assign array_update_73792[0] = add_73368 == 32'h0000_0000 ? array_update_73790 : array_update_73779[0];
  assign array_update_73792[1] = add_73368 == 32'h0000_0001 ? array_update_73790 : array_update_73779[1];
  assign array_update_73792[2] = add_73368 == 32'h0000_0002 ? array_update_73790 : array_update_73779[2];
  assign array_update_73792[3] = add_73368 == 32'h0000_0003 ? array_update_73790 : array_update_73779[3];
  assign array_update_73792[4] = add_73368 == 32'h0000_0004 ? array_update_73790 : array_update_73779[4];
  assign array_update_73792[5] = add_73368 == 32'h0000_0005 ? array_update_73790 : array_update_73779[5];
  assign array_update_73792[6] = add_73368 == 32'h0000_0006 ? array_update_73790 : array_update_73779[6];
  assign array_update_73792[7] = add_73368 == 32'h0000_0007 ? array_update_73790 : array_update_73779[7];
  assign array_update_73792[8] = add_73368 == 32'h0000_0008 ? array_update_73790 : array_update_73779[8];
  assign array_update_73792[9] = add_73368 == 32'h0000_0009 ? array_update_73790 : array_update_73779[9];
  assign array_index_73794 = array_update_72021[add_73791 > 32'h0000_0009 ? 4'h9 : add_73791[3:0]];
  assign array_index_73795 = array_update_73792[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_73799 = smul32b_32b_x_32b(array_index_73375[add_73791 > 32'h0000_0009 ? 4'h9 : add_73791[3:0]], array_index_73794[add_73776 > 32'h0000_0009 ? 4'h9 : add_73776[3:0]]);
  assign add_73801 = array_index_73795[add_73776 > 32'h0000_0009 ? 4'h9 : add_73776[3:0]] + smul_73799;
  assign array_update_73803[0] = add_73776 == 32'h0000_0000 ? add_73801 : array_index_73795[0];
  assign array_update_73803[1] = add_73776 == 32'h0000_0001 ? add_73801 : array_index_73795[1];
  assign array_update_73803[2] = add_73776 == 32'h0000_0002 ? add_73801 : array_index_73795[2];
  assign array_update_73803[3] = add_73776 == 32'h0000_0003 ? add_73801 : array_index_73795[3];
  assign array_update_73803[4] = add_73776 == 32'h0000_0004 ? add_73801 : array_index_73795[4];
  assign array_update_73803[5] = add_73776 == 32'h0000_0005 ? add_73801 : array_index_73795[5];
  assign array_update_73803[6] = add_73776 == 32'h0000_0006 ? add_73801 : array_index_73795[6];
  assign array_update_73803[7] = add_73776 == 32'h0000_0007 ? add_73801 : array_index_73795[7];
  assign array_update_73803[8] = add_73776 == 32'h0000_0008 ? add_73801 : array_index_73795[8];
  assign array_update_73803[9] = add_73776 == 32'h0000_0009 ? add_73801 : array_index_73795[9];
  assign add_73804 = add_73791 + 32'h0000_0001;
  assign array_update_73805[0] = add_73368 == 32'h0000_0000 ? array_update_73803 : array_update_73792[0];
  assign array_update_73805[1] = add_73368 == 32'h0000_0001 ? array_update_73803 : array_update_73792[1];
  assign array_update_73805[2] = add_73368 == 32'h0000_0002 ? array_update_73803 : array_update_73792[2];
  assign array_update_73805[3] = add_73368 == 32'h0000_0003 ? array_update_73803 : array_update_73792[3];
  assign array_update_73805[4] = add_73368 == 32'h0000_0004 ? array_update_73803 : array_update_73792[4];
  assign array_update_73805[5] = add_73368 == 32'h0000_0005 ? array_update_73803 : array_update_73792[5];
  assign array_update_73805[6] = add_73368 == 32'h0000_0006 ? array_update_73803 : array_update_73792[6];
  assign array_update_73805[7] = add_73368 == 32'h0000_0007 ? array_update_73803 : array_update_73792[7];
  assign array_update_73805[8] = add_73368 == 32'h0000_0008 ? array_update_73803 : array_update_73792[8];
  assign array_update_73805[9] = add_73368 == 32'h0000_0009 ? array_update_73803 : array_update_73792[9];
  assign array_index_73807 = array_update_72021[add_73804 > 32'h0000_0009 ? 4'h9 : add_73804[3:0]];
  assign array_index_73808 = array_update_73805[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_73812 = smul32b_32b_x_32b(array_index_73375[add_73804 > 32'h0000_0009 ? 4'h9 : add_73804[3:0]], array_index_73807[add_73776 > 32'h0000_0009 ? 4'h9 : add_73776[3:0]]);
  assign add_73814 = array_index_73808[add_73776 > 32'h0000_0009 ? 4'h9 : add_73776[3:0]] + smul_73812;
  assign array_update_73816[0] = add_73776 == 32'h0000_0000 ? add_73814 : array_index_73808[0];
  assign array_update_73816[1] = add_73776 == 32'h0000_0001 ? add_73814 : array_index_73808[1];
  assign array_update_73816[2] = add_73776 == 32'h0000_0002 ? add_73814 : array_index_73808[2];
  assign array_update_73816[3] = add_73776 == 32'h0000_0003 ? add_73814 : array_index_73808[3];
  assign array_update_73816[4] = add_73776 == 32'h0000_0004 ? add_73814 : array_index_73808[4];
  assign array_update_73816[5] = add_73776 == 32'h0000_0005 ? add_73814 : array_index_73808[5];
  assign array_update_73816[6] = add_73776 == 32'h0000_0006 ? add_73814 : array_index_73808[6];
  assign array_update_73816[7] = add_73776 == 32'h0000_0007 ? add_73814 : array_index_73808[7];
  assign array_update_73816[8] = add_73776 == 32'h0000_0008 ? add_73814 : array_index_73808[8];
  assign array_update_73816[9] = add_73776 == 32'h0000_0009 ? add_73814 : array_index_73808[9];
  assign add_73817 = add_73804 + 32'h0000_0001;
  assign array_update_73818[0] = add_73368 == 32'h0000_0000 ? array_update_73816 : array_update_73805[0];
  assign array_update_73818[1] = add_73368 == 32'h0000_0001 ? array_update_73816 : array_update_73805[1];
  assign array_update_73818[2] = add_73368 == 32'h0000_0002 ? array_update_73816 : array_update_73805[2];
  assign array_update_73818[3] = add_73368 == 32'h0000_0003 ? array_update_73816 : array_update_73805[3];
  assign array_update_73818[4] = add_73368 == 32'h0000_0004 ? array_update_73816 : array_update_73805[4];
  assign array_update_73818[5] = add_73368 == 32'h0000_0005 ? array_update_73816 : array_update_73805[5];
  assign array_update_73818[6] = add_73368 == 32'h0000_0006 ? array_update_73816 : array_update_73805[6];
  assign array_update_73818[7] = add_73368 == 32'h0000_0007 ? array_update_73816 : array_update_73805[7];
  assign array_update_73818[8] = add_73368 == 32'h0000_0008 ? array_update_73816 : array_update_73805[8];
  assign array_update_73818[9] = add_73368 == 32'h0000_0009 ? array_update_73816 : array_update_73805[9];
  assign array_index_73820 = array_update_72021[add_73817 > 32'h0000_0009 ? 4'h9 : add_73817[3:0]];
  assign array_index_73821 = array_update_73818[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_73825 = smul32b_32b_x_32b(array_index_73375[add_73817 > 32'h0000_0009 ? 4'h9 : add_73817[3:0]], array_index_73820[add_73776 > 32'h0000_0009 ? 4'h9 : add_73776[3:0]]);
  assign add_73827 = array_index_73821[add_73776 > 32'h0000_0009 ? 4'h9 : add_73776[3:0]] + smul_73825;
  assign array_update_73829[0] = add_73776 == 32'h0000_0000 ? add_73827 : array_index_73821[0];
  assign array_update_73829[1] = add_73776 == 32'h0000_0001 ? add_73827 : array_index_73821[1];
  assign array_update_73829[2] = add_73776 == 32'h0000_0002 ? add_73827 : array_index_73821[2];
  assign array_update_73829[3] = add_73776 == 32'h0000_0003 ? add_73827 : array_index_73821[3];
  assign array_update_73829[4] = add_73776 == 32'h0000_0004 ? add_73827 : array_index_73821[4];
  assign array_update_73829[5] = add_73776 == 32'h0000_0005 ? add_73827 : array_index_73821[5];
  assign array_update_73829[6] = add_73776 == 32'h0000_0006 ? add_73827 : array_index_73821[6];
  assign array_update_73829[7] = add_73776 == 32'h0000_0007 ? add_73827 : array_index_73821[7];
  assign array_update_73829[8] = add_73776 == 32'h0000_0008 ? add_73827 : array_index_73821[8];
  assign array_update_73829[9] = add_73776 == 32'h0000_0009 ? add_73827 : array_index_73821[9];
  assign add_73830 = add_73817 + 32'h0000_0001;
  assign array_update_73831[0] = add_73368 == 32'h0000_0000 ? array_update_73829 : array_update_73818[0];
  assign array_update_73831[1] = add_73368 == 32'h0000_0001 ? array_update_73829 : array_update_73818[1];
  assign array_update_73831[2] = add_73368 == 32'h0000_0002 ? array_update_73829 : array_update_73818[2];
  assign array_update_73831[3] = add_73368 == 32'h0000_0003 ? array_update_73829 : array_update_73818[3];
  assign array_update_73831[4] = add_73368 == 32'h0000_0004 ? array_update_73829 : array_update_73818[4];
  assign array_update_73831[5] = add_73368 == 32'h0000_0005 ? array_update_73829 : array_update_73818[5];
  assign array_update_73831[6] = add_73368 == 32'h0000_0006 ? array_update_73829 : array_update_73818[6];
  assign array_update_73831[7] = add_73368 == 32'h0000_0007 ? array_update_73829 : array_update_73818[7];
  assign array_update_73831[8] = add_73368 == 32'h0000_0008 ? array_update_73829 : array_update_73818[8];
  assign array_update_73831[9] = add_73368 == 32'h0000_0009 ? array_update_73829 : array_update_73818[9];
  assign array_index_73833 = array_update_72021[add_73830 > 32'h0000_0009 ? 4'h9 : add_73830[3:0]];
  assign array_index_73834 = array_update_73831[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_73838 = smul32b_32b_x_32b(array_index_73375[add_73830 > 32'h0000_0009 ? 4'h9 : add_73830[3:0]], array_index_73833[add_73776 > 32'h0000_0009 ? 4'h9 : add_73776[3:0]]);
  assign add_73840 = array_index_73834[add_73776 > 32'h0000_0009 ? 4'h9 : add_73776[3:0]] + smul_73838;
  assign array_update_73842[0] = add_73776 == 32'h0000_0000 ? add_73840 : array_index_73834[0];
  assign array_update_73842[1] = add_73776 == 32'h0000_0001 ? add_73840 : array_index_73834[1];
  assign array_update_73842[2] = add_73776 == 32'h0000_0002 ? add_73840 : array_index_73834[2];
  assign array_update_73842[3] = add_73776 == 32'h0000_0003 ? add_73840 : array_index_73834[3];
  assign array_update_73842[4] = add_73776 == 32'h0000_0004 ? add_73840 : array_index_73834[4];
  assign array_update_73842[5] = add_73776 == 32'h0000_0005 ? add_73840 : array_index_73834[5];
  assign array_update_73842[6] = add_73776 == 32'h0000_0006 ? add_73840 : array_index_73834[6];
  assign array_update_73842[7] = add_73776 == 32'h0000_0007 ? add_73840 : array_index_73834[7];
  assign array_update_73842[8] = add_73776 == 32'h0000_0008 ? add_73840 : array_index_73834[8];
  assign array_update_73842[9] = add_73776 == 32'h0000_0009 ? add_73840 : array_index_73834[9];
  assign add_73843 = add_73830 + 32'h0000_0001;
  assign array_update_73844[0] = add_73368 == 32'h0000_0000 ? array_update_73842 : array_update_73831[0];
  assign array_update_73844[1] = add_73368 == 32'h0000_0001 ? array_update_73842 : array_update_73831[1];
  assign array_update_73844[2] = add_73368 == 32'h0000_0002 ? array_update_73842 : array_update_73831[2];
  assign array_update_73844[3] = add_73368 == 32'h0000_0003 ? array_update_73842 : array_update_73831[3];
  assign array_update_73844[4] = add_73368 == 32'h0000_0004 ? array_update_73842 : array_update_73831[4];
  assign array_update_73844[5] = add_73368 == 32'h0000_0005 ? array_update_73842 : array_update_73831[5];
  assign array_update_73844[6] = add_73368 == 32'h0000_0006 ? array_update_73842 : array_update_73831[6];
  assign array_update_73844[7] = add_73368 == 32'h0000_0007 ? array_update_73842 : array_update_73831[7];
  assign array_update_73844[8] = add_73368 == 32'h0000_0008 ? array_update_73842 : array_update_73831[8];
  assign array_update_73844[9] = add_73368 == 32'h0000_0009 ? array_update_73842 : array_update_73831[9];
  assign array_index_73846 = array_update_72021[add_73843 > 32'h0000_0009 ? 4'h9 : add_73843[3:0]];
  assign array_index_73847 = array_update_73844[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_73851 = smul32b_32b_x_32b(array_index_73375[add_73843 > 32'h0000_0009 ? 4'h9 : add_73843[3:0]], array_index_73846[add_73776 > 32'h0000_0009 ? 4'h9 : add_73776[3:0]]);
  assign add_73853 = array_index_73847[add_73776 > 32'h0000_0009 ? 4'h9 : add_73776[3:0]] + smul_73851;
  assign array_update_73855[0] = add_73776 == 32'h0000_0000 ? add_73853 : array_index_73847[0];
  assign array_update_73855[1] = add_73776 == 32'h0000_0001 ? add_73853 : array_index_73847[1];
  assign array_update_73855[2] = add_73776 == 32'h0000_0002 ? add_73853 : array_index_73847[2];
  assign array_update_73855[3] = add_73776 == 32'h0000_0003 ? add_73853 : array_index_73847[3];
  assign array_update_73855[4] = add_73776 == 32'h0000_0004 ? add_73853 : array_index_73847[4];
  assign array_update_73855[5] = add_73776 == 32'h0000_0005 ? add_73853 : array_index_73847[5];
  assign array_update_73855[6] = add_73776 == 32'h0000_0006 ? add_73853 : array_index_73847[6];
  assign array_update_73855[7] = add_73776 == 32'h0000_0007 ? add_73853 : array_index_73847[7];
  assign array_update_73855[8] = add_73776 == 32'h0000_0008 ? add_73853 : array_index_73847[8];
  assign array_update_73855[9] = add_73776 == 32'h0000_0009 ? add_73853 : array_index_73847[9];
  assign add_73856 = add_73843 + 32'h0000_0001;
  assign array_update_73857[0] = add_73368 == 32'h0000_0000 ? array_update_73855 : array_update_73844[0];
  assign array_update_73857[1] = add_73368 == 32'h0000_0001 ? array_update_73855 : array_update_73844[1];
  assign array_update_73857[2] = add_73368 == 32'h0000_0002 ? array_update_73855 : array_update_73844[2];
  assign array_update_73857[3] = add_73368 == 32'h0000_0003 ? array_update_73855 : array_update_73844[3];
  assign array_update_73857[4] = add_73368 == 32'h0000_0004 ? array_update_73855 : array_update_73844[4];
  assign array_update_73857[5] = add_73368 == 32'h0000_0005 ? array_update_73855 : array_update_73844[5];
  assign array_update_73857[6] = add_73368 == 32'h0000_0006 ? array_update_73855 : array_update_73844[6];
  assign array_update_73857[7] = add_73368 == 32'h0000_0007 ? array_update_73855 : array_update_73844[7];
  assign array_update_73857[8] = add_73368 == 32'h0000_0008 ? array_update_73855 : array_update_73844[8];
  assign array_update_73857[9] = add_73368 == 32'h0000_0009 ? array_update_73855 : array_update_73844[9];
  assign array_index_73859 = array_update_72021[add_73856 > 32'h0000_0009 ? 4'h9 : add_73856[3:0]];
  assign array_index_73860 = array_update_73857[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_73864 = smul32b_32b_x_32b(array_index_73375[add_73856 > 32'h0000_0009 ? 4'h9 : add_73856[3:0]], array_index_73859[add_73776 > 32'h0000_0009 ? 4'h9 : add_73776[3:0]]);
  assign add_73866 = array_index_73860[add_73776 > 32'h0000_0009 ? 4'h9 : add_73776[3:0]] + smul_73864;
  assign array_update_73868[0] = add_73776 == 32'h0000_0000 ? add_73866 : array_index_73860[0];
  assign array_update_73868[1] = add_73776 == 32'h0000_0001 ? add_73866 : array_index_73860[1];
  assign array_update_73868[2] = add_73776 == 32'h0000_0002 ? add_73866 : array_index_73860[2];
  assign array_update_73868[3] = add_73776 == 32'h0000_0003 ? add_73866 : array_index_73860[3];
  assign array_update_73868[4] = add_73776 == 32'h0000_0004 ? add_73866 : array_index_73860[4];
  assign array_update_73868[5] = add_73776 == 32'h0000_0005 ? add_73866 : array_index_73860[5];
  assign array_update_73868[6] = add_73776 == 32'h0000_0006 ? add_73866 : array_index_73860[6];
  assign array_update_73868[7] = add_73776 == 32'h0000_0007 ? add_73866 : array_index_73860[7];
  assign array_update_73868[8] = add_73776 == 32'h0000_0008 ? add_73866 : array_index_73860[8];
  assign array_update_73868[9] = add_73776 == 32'h0000_0009 ? add_73866 : array_index_73860[9];
  assign add_73869 = add_73856 + 32'h0000_0001;
  assign array_update_73870[0] = add_73368 == 32'h0000_0000 ? array_update_73868 : array_update_73857[0];
  assign array_update_73870[1] = add_73368 == 32'h0000_0001 ? array_update_73868 : array_update_73857[1];
  assign array_update_73870[2] = add_73368 == 32'h0000_0002 ? array_update_73868 : array_update_73857[2];
  assign array_update_73870[3] = add_73368 == 32'h0000_0003 ? array_update_73868 : array_update_73857[3];
  assign array_update_73870[4] = add_73368 == 32'h0000_0004 ? array_update_73868 : array_update_73857[4];
  assign array_update_73870[5] = add_73368 == 32'h0000_0005 ? array_update_73868 : array_update_73857[5];
  assign array_update_73870[6] = add_73368 == 32'h0000_0006 ? array_update_73868 : array_update_73857[6];
  assign array_update_73870[7] = add_73368 == 32'h0000_0007 ? array_update_73868 : array_update_73857[7];
  assign array_update_73870[8] = add_73368 == 32'h0000_0008 ? array_update_73868 : array_update_73857[8];
  assign array_update_73870[9] = add_73368 == 32'h0000_0009 ? array_update_73868 : array_update_73857[9];
  assign array_index_73872 = array_update_72021[add_73869 > 32'h0000_0009 ? 4'h9 : add_73869[3:0]];
  assign array_index_73873 = array_update_73870[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_73877 = smul32b_32b_x_32b(array_index_73375[add_73869 > 32'h0000_0009 ? 4'h9 : add_73869[3:0]], array_index_73872[add_73776 > 32'h0000_0009 ? 4'h9 : add_73776[3:0]]);
  assign add_73879 = array_index_73873[add_73776 > 32'h0000_0009 ? 4'h9 : add_73776[3:0]] + smul_73877;
  assign array_update_73881[0] = add_73776 == 32'h0000_0000 ? add_73879 : array_index_73873[0];
  assign array_update_73881[1] = add_73776 == 32'h0000_0001 ? add_73879 : array_index_73873[1];
  assign array_update_73881[2] = add_73776 == 32'h0000_0002 ? add_73879 : array_index_73873[2];
  assign array_update_73881[3] = add_73776 == 32'h0000_0003 ? add_73879 : array_index_73873[3];
  assign array_update_73881[4] = add_73776 == 32'h0000_0004 ? add_73879 : array_index_73873[4];
  assign array_update_73881[5] = add_73776 == 32'h0000_0005 ? add_73879 : array_index_73873[5];
  assign array_update_73881[6] = add_73776 == 32'h0000_0006 ? add_73879 : array_index_73873[6];
  assign array_update_73881[7] = add_73776 == 32'h0000_0007 ? add_73879 : array_index_73873[7];
  assign array_update_73881[8] = add_73776 == 32'h0000_0008 ? add_73879 : array_index_73873[8];
  assign array_update_73881[9] = add_73776 == 32'h0000_0009 ? add_73879 : array_index_73873[9];
  assign add_73882 = add_73869 + 32'h0000_0001;
  assign array_update_73883[0] = add_73368 == 32'h0000_0000 ? array_update_73881 : array_update_73870[0];
  assign array_update_73883[1] = add_73368 == 32'h0000_0001 ? array_update_73881 : array_update_73870[1];
  assign array_update_73883[2] = add_73368 == 32'h0000_0002 ? array_update_73881 : array_update_73870[2];
  assign array_update_73883[3] = add_73368 == 32'h0000_0003 ? array_update_73881 : array_update_73870[3];
  assign array_update_73883[4] = add_73368 == 32'h0000_0004 ? array_update_73881 : array_update_73870[4];
  assign array_update_73883[5] = add_73368 == 32'h0000_0005 ? array_update_73881 : array_update_73870[5];
  assign array_update_73883[6] = add_73368 == 32'h0000_0006 ? array_update_73881 : array_update_73870[6];
  assign array_update_73883[7] = add_73368 == 32'h0000_0007 ? array_update_73881 : array_update_73870[7];
  assign array_update_73883[8] = add_73368 == 32'h0000_0008 ? array_update_73881 : array_update_73870[8];
  assign array_update_73883[9] = add_73368 == 32'h0000_0009 ? array_update_73881 : array_update_73870[9];
  assign array_index_73885 = array_update_72021[add_73882 > 32'h0000_0009 ? 4'h9 : add_73882[3:0]];
  assign array_index_73886 = array_update_73883[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_73890 = smul32b_32b_x_32b(array_index_73375[add_73882 > 32'h0000_0009 ? 4'h9 : add_73882[3:0]], array_index_73885[add_73776 > 32'h0000_0009 ? 4'h9 : add_73776[3:0]]);
  assign add_73892 = array_index_73886[add_73776 > 32'h0000_0009 ? 4'h9 : add_73776[3:0]] + smul_73890;
  assign array_update_73894[0] = add_73776 == 32'h0000_0000 ? add_73892 : array_index_73886[0];
  assign array_update_73894[1] = add_73776 == 32'h0000_0001 ? add_73892 : array_index_73886[1];
  assign array_update_73894[2] = add_73776 == 32'h0000_0002 ? add_73892 : array_index_73886[2];
  assign array_update_73894[3] = add_73776 == 32'h0000_0003 ? add_73892 : array_index_73886[3];
  assign array_update_73894[4] = add_73776 == 32'h0000_0004 ? add_73892 : array_index_73886[4];
  assign array_update_73894[5] = add_73776 == 32'h0000_0005 ? add_73892 : array_index_73886[5];
  assign array_update_73894[6] = add_73776 == 32'h0000_0006 ? add_73892 : array_index_73886[6];
  assign array_update_73894[7] = add_73776 == 32'h0000_0007 ? add_73892 : array_index_73886[7];
  assign array_update_73894[8] = add_73776 == 32'h0000_0008 ? add_73892 : array_index_73886[8];
  assign array_update_73894[9] = add_73776 == 32'h0000_0009 ? add_73892 : array_index_73886[9];
  assign add_73895 = add_73882 + 32'h0000_0001;
  assign array_update_73896[0] = add_73368 == 32'h0000_0000 ? array_update_73894 : array_update_73883[0];
  assign array_update_73896[1] = add_73368 == 32'h0000_0001 ? array_update_73894 : array_update_73883[1];
  assign array_update_73896[2] = add_73368 == 32'h0000_0002 ? array_update_73894 : array_update_73883[2];
  assign array_update_73896[3] = add_73368 == 32'h0000_0003 ? array_update_73894 : array_update_73883[3];
  assign array_update_73896[4] = add_73368 == 32'h0000_0004 ? array_update_73894 : array_update_73883[4];
  assign array_update_73896[5] = add_73368 == 32'h0000_0005 ? array_update_73894 : array_update_73883[5];
  assign array_update_73896[6] = add_73368 == 32'h0000_0006 ? array_update_73894 : array_update_73883[6];
  assign array_update_73896[7] = add_73368 == 32'h0000_0007 ? array_update_73894 : array_update_73883[7];
  assign array_update_73896[8] = add_73368 == 32'h0000_0008 ? array_update_73894 : array_update_73883[8];
  assign array_update_73896[9] = add_73368 == 32'h0000_0009 ? array_update_73894 : array_update_73883[9];
  assign array_index_73898 = array_update_72021[add_73895 > 32'h0000_0009 ? 4'h9 : add_73895[3:0]];
  assign array_index_73899 = array_update_73896[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_73903 = smul32b_32b_x_32b(array_index_73375[add_73895 > 32'h0000_0009 ? 4'h9 : add_73895[3:0]], array_index_73898[add_73776 > 32'h0000_0009 ? 4'h9 : add_73776[3:0]]);
  assign add_73905 = array_index_73899[add_73776 > 32'h0000_0009 ? 4'h9 : add_73776[3:0]] + smul_73903;
  assign array_update_73906[0] = add_73776 == 32'h0000_0000 ? add_73905 : array_index_73899[0];
  assign array_update_73906[1] = add_73776 == 32'h0000_0001 ? add_73905 : array_index_73899[1];
  assign array_update_73906[2] = add_73776 == 32'h0000_0002 ? add_73905 : array_index_73899[2];
  assign array_update_73906[3] = add_73776 == 32'h0000_0003 ? add_73905 : array_index_73899[3];
  assign array_update_73906[4] = add_73776 == 32'h0000_0004 ? add_73905 : array_index_73899[4];
  assign array_update_73906[5] = add_73776 == 32'h0000_0005 ? add_73905 : array_index_73899[5];
  assign array_update_73906[6] = add_73776 == 32'h0000_0006 ? add_73905 : array_index_73899[6];
  assign array_update_73906[7] = add_73776 == 32'h0000_0007 ? add_73905 : array_index_73899[7];
  assign array_update_73906[8] = add_73776 == 32'h0000_0008 ? add_73905 : array_index_73899[8];
  assign array_update_73906[9] = add_73776 == 32'h0000_0009 ? add_73905 : array_index_73899[9];
  assign array_update_73907[0] = add_73368 == 32'h0000_0000 ? array_update_73906 : array_update_73896[0];
  assign array_update_73907[1] = add_73368 == 32'h0000_0001 ? array_update_73906 : array_update_73896[1];
  assign array_update_73907[2] = add_73368 == 32'h0000_0002 ? array_update_73906 : array_update_73896[2];
  assign array_update_73907[3] = add_73368 == 32'h0000_0003 ? array_update_73906 : array_update_73896[3];
  assign array_update_73907[4] = add_73368 == 32'h0000_0004 ? array_update_73906 : array_update_73896[4];
  assign array_update_73907[5] = add_73368 == 32'h0000_0005 ? array_update_73906 : array_update_73896[5];
  assign array_update_73907[6] = add_73368 == 32'h0000_0006 ? array_update_73906 : array_update_73896[6];
  assign array_update_73907[7] = add_73368 == 32'h0000_0007 ? array_update_73906 : array_update_73896[7];
  assign array_update_73907[8] = add_73368 == 32'h0000_0008 ? array_update_73906 : array_update_73896[8];
  assign array_update_73907[9] = add_73368 == 32'h0000_0009 ? array_update_73906 : array_update_73896[9];
  assign array_index_73909 = array_update_73907[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign add_73911 = add_73776 + 32'h0000_0001;
  assign array_update_73912[0] = add_73911 == 32'h0000_0000 ? 32'h0000_0000 : array_index_73909[0];
  assign array_update_73912[1] = add_73911 == 32'h0000_0001 ? 32'h0000_0000 : array_index_73909[1];
  assign array_update_73912[2] = add_73911 == 32'h0000_0002 ? 32'h0000_0000 : array_index_73909[2];
  assign array_update_73912[3] = add_73911 == 32'h0000_0003 ? 32'h0000_0000 : array_index_73909[3];
  assign array_update_73912[4] = add_73911 == 32'h0000_0004 ? 32'h0000_0000 : array_index_73909[4];
  assign array_update_73912[5] = add_73911 == 32'h0000_0005 ? 32'h0000_0000 : array_index_73909[5];
  assign array_update_73912[6] = add_73911 == 32'h0000_0006 ? 32'h0000_0000 : array_index_73909[6];
  assign array_update_73912[7] = add_73911 == 32'h0000_0007 ? 32'h0000_0000 : array_index_73909[7];
  assign array_update_73912[8] = add_73911 == 32'h0000_0008 ? 32'h0000_0000 : array_index_73909[8];
  assign array_update_73912[9] = add_73911 == 32'h0000_0009 ? 32'h0000_0000 : array_index_73909[9];
  assign literal_73913 = 32'h0000_0000;
  assign array_update_73914[0] = add_73368 == 32'h0000_0000 ? array_update_73912 : array_update_73907[0];
  assign array_update_73914[1] = add_73368 == 32'h0000_0001 ? array_update_73912 : array_update_73907[1];
  assign array_update_73914[2] = add_73368 == 32'h0000_0002 ? array_update_73912 : array_update_73907[2];
  assign array_update_73914[3] = add_73368 == 32'h0000_0003 ? array_update_73912 : array_update_73907[3];
  assign array_update_73914[4] = add_73368 == 32'h0000_0004 ? array_update_73912 : array_update_73907[4];
  assign array_update_73914[5] = add_73368 == 32'h0000_0005 ? array_update_73912 : array_update_73907[5];
  assign array_update_73914[6] = add_73368 == 32'h0000_0006 ? array_update_73912 : array_update_73907[6];
  assign array_update_73914[7] = add_73368 == 32'h0000_0007 ? array_update_73912 : array_update_73907[7];
  assign array_update_73914[8] = add_73368 == 32'h0000_0008 ? array_update_73912 : array_update_73907[8];
  assign array_update_73914[9] = add_73368 == 32'h0000_0009 ? array_update_73912 : array_update_73907[9];
  assign array_index_73916 = array_update_72021[literal_73913 > 32'h0000_0009 ? 4'h9 : literal_73913[3:0]];
  assign array_index_73917 = array_update_73914[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_73921 = smul32b_32b_x_32b(array_index_73375[literal_73913 > 32'h0000_0009 ? 4'h9 : literal_73913[3:0]], array_index_73916[add_73911 > 32'h0000_0009 ? 4'h9 : add_73911[3:0]]);
  assign add_73923 = array_index_73917[add_73911 > 32'h0000_0009 ? 4'h9 : add_73911[3:0]] + smul_73921;
  assign array_update_73925[0] = add_73911 == 32'h0000_0000 ? add_73923 : array_index_73917[0];
  assign array_update_73925[1] = add_73911 == 32'h0000_0001 ? add_73923 : array_index_73917[1];
  assign array_update_73925[2] = add_73911 == 32'h0000_0002 ? add_73923 : array_index_73917[2];
  assign array_update_73925[3] = add_73911 == 32'h0000_0003 ? add_73923 : array_index_73917[3];
  assign array_update_73925[4] = add_73911 == 32'h0000_0004 ? add_73923 : array_index_73917[4];
  assign array_update_73925[5] = add_73911 == 32'h0000_0005 ? add_73923 : array_index_73917[5];
  assign array_update_73925[6] = add_73911 == 32'h0000_0006 ? add_73923 : array_index_73917[6];
  assign array_update_73925[7] = add_73911 == 32'h0000_0007 ? add_73923 : array_index_73917[7];
  assign array_update_73925[8] = add_73911 == 32'h0000_0008 ? add_73923 : array_index_73917[8];
  assign array_update_73925[9] = add_73911 == 32'h0000_0009 ? add_73923 : array_index_73917[9];
  assign add_73926 = literal_73913 + 32'h0000_0001;
  assign array_update_73927[0] = add_73368 == 32'h0000_0000 ? array_update_73925 : array_update_73914[0];
  assign array_update_73927[1] = add_73368 == 32'h0000_0001 ? array_update_73925 : array_update_73914[1];
  assign array_update_73927[2] = add_73368 == 32'h0000_0002 ? array_update_73925 : array_update_73914[2];
  assign array_update_73927[3] = add_73368 == 32'h0000_0003 ? array_update_73925 : array_update_73914[3];
  assign array_update_73927[4] = add_73368 == 32'h0000_0004 ? array_update_73925 : array_update_73914[4];
  assign array_update_73927[5] = add_73368 == 32'h0000_0005 ? array_update_73925 : array_update_73914[5];
  assign array_update_73927[6] = add_73368 == 32'h0000_0006 ? array_update_73925 : array_update_73914[6];
  assign array_update_73927[7] = add_73368 == 32'h0000_0007 ? array_update_73925 : array_update_73914[7];
  assign array_update_73927[8] = add_73368 == 32'h0000_0008 ? array_update_73925 : array_update_73914[8];
  assign array_update_73927[9] = add_73368 == 32'h0000_0009 ? array_update_73925 : array_update_73914[9];
  assign array_index_73929 = array_update_72021[add_73926 > 32'h0000_0009 ? 4'h9 : add_73926[3:0]];
  assign array_index_73930 = array_update_73927[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_73934 = smul32b_32b_x_32b(array_index_73375[add_73926 > 32'h0000_0009 ? 4'h9 : add_73926[3:0]], array_index_73929[add_73911 > 32'h0000_0009 ? 4'h9 : add_73911[3:0]]);
  assign add_73936 = array_index_73930[add_73911 > 32'h0000_0009 ? 4'h9 : add_73911[3:0]] + smul_73934;
  assign array_update_73938[0] = add_73911 == 32'h0000_0000 ? add_73936 : array_index_73930[0];
  assign array_update_73938[1] = add_73911 == 32'h0000_0001 ? add_73936 : array_index_73930[1];
  assign array_update_73938[2] = add_73911 == 32'h0000_0002 ? add_73936 : array_index_73930[2];
  assign array_update_73938[3] = add_73911 == 32'h0000_0003 ? add_73936 : array_index_73930[3];
  assign array_update_73938[4] = add_73911 == 32'h0000_0004 ? add_73936 : array_index_73930[4];
  assign array_update_73938[5] = add_73911 == 32'h0000_0005 ? add_73936 : array_index_73930[5];
  assign array_update_73938[6] = add_73911 == 32'h0000_0006 ? add_73936 : array_index_73930[6];
  assign array_update_73938[7] = add_73911 == 32'h0000_0007 ? add_73936 : array_index_73930[7];
  assign array_update_73938[8] = add_73911 == 32'h0000_0008 ? add_73936 : array_index_73930[8];
  assign array_update_73938[9] = add_73911 == 32'h0000_0009 ? add_73936 : array_index_73930[9];
  assign add_73939 = add_73926 + 32'h0000_0001;
  assign array_update_73940[0] = add_73368 == 32'h0000_0000 ? array_update_73938 : array_update_73927[0];
  assign array_update_73940[1] = add_73368 == 32'h0000_0001 ? array_update_73938 : array_update_73927[1];
  assign array_update_73940[2] = add_73368 == 32'h0000_0002 ? array_update_73938 : array_update_73927[2];
  assign array_update_73940[3] = add_73368 == 32'h0000_0003 ? array_update_73938 : array_update_73927[3];
  assign array_update_73940[4] = add_73368 == 32'h0000_0004 ? array_update_73938 : array_update_73927[4];
  assign array_update_73940[5] = add_73368 == 32'h0000_0005 ? array_update_73938 : array_update_73927[5];
  assign array_update_73940[6] = add_73368 == 32'h0000_0006 ? array_update_73938 : array_update_73927[6];
  assign array_update_73940[7] = add_73368 == 32'h0000_0007 ? array_update_73938 : array_update_73927[7];
  assign array_update_73940[8] = add_73368 == 32'h0000_0008 ? array_update_73938 : array_update_73927[8];
  assign array_update_73940[9] = add_73368 == 32'h0000_0009 ? array_update_73938 : array_update_73927[9];
  assign array_index_73942 = array_update_72021[add_73939 > 32'h0000_0009 ? 4'h9 : add_73939[3:0]];
  assign array_index_73943 = array_update_73940[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_73947 = smul32b_32b_x_32b(array_index_73375[add_73939 > 32'h0000_0009 ? 4'h9 : add_73939[3:0]], array_index_73942[add_73911 > 32'h0000_0009 ? 4'h9 : add_73911[3:0]]);
  assign add_73949 = array_index_73943[add_73911 > 32'h0000_0009 ? 4'h9 : add_73911[3:0]] + smul_73947;
  assign array_update_73951[0] = add_73911 == 32'h0000_0000 ? add_73949 : array_index_73943[0];
  assign array_update_73951[1] = add_73911 == 32'h0000_0001 ? add_73949 : array_index_73943[1];
  assign array_update_73951[2] = add_73911 == 32'h0000_0002 ? add_73949 : array_index_73943[2];
  assign array_update_73951[3] = add_73911 == 32'h0000_0003 ? add_73949 : array_index_73943[3];
  assign array_update_73951[4] = add_73911 == 32'h0000_0004 ? add_73949 : array_index_73943[4];
  assign array_update_73951[5] = add_73911 == 32'h0000_0005 ? add_73949 : array_index_73943[5];
  assign array_update_73951[6] = add_73911 == 32'h0000_0006 ? add_73949 : array_index_73943[6];
  assign array_update_73951[7] = add_73911 == 32'h0000_0007 ? add_73949 : array_index_73943[7];
  assign array_update_73951[8] = add_73911 == 32'h0000_0008 ? add_73949 : array_index_73943[8];
  assign array_update_73951[9] = add_73911 == 32'h0000_0009 ? add_73949 : array_index_73943[9];
  assign add_73952 = add_73939 + 32'h0000_0001;
  assign array_update_73953[0] = add_73368 == 32'h0000_0000 ? array_update_73951 : array_update_73940[0];
  assign array_update_73953[1] = add_73368 == 32'h0000_0001 ? array_update_73951 : array_update_73940[1];
  assign array_update_73953[2] = add_73368 == 32'h0000_0002 ? array_update_73951 : array_update_73940[2];
  assign array_update_73953[3] = add_73368 == 32'h0000_0003 ? array_update_73951 : array_update_73940[3];
  assign array_update_73953[4] = add_73368 == 32'h0000_0004 ? array_update_73951 : array_update_73940[4];
  assign array_update_73953[5] = add_73368 == 32'h0000_0005 ? array_update_73951 : array_update_73940[5];
  assign array_update_73953[6] = add_73368 == 32'h0000_0006 ? array_update_73951 : array_update_73940[6];
  assign array_update_73953[7] = add_73368 == 32'h0000_0007 ? array_update_73951 : array_update_73940[7];
  assign array_update_73953[8] = add_73368 == 32'h0000_0008 ? array_update_73951 : array_update_73940[8];
  assign array_update_73953[9] = add_73368 == 32'h0000_0009 ? array_update_73951 : array_update_73940[9];
  assign array_index_73955 = array_update_72021[add_73952 > 32'h0000_0009 ? 4'h9 : add_73952[3:0]];
  assign array_index_73956 = array_update_73953[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_73960 = smul32b_32b_x_32b(array_index_73375[add_73952 > 32'h0000_0009 ? 4'h9 : add_73952[3:0]], array_index_73955[add_73911 > 32'h0000_0009 ? 4'h9 : add_73911[3:0]]);
  assign add_73962 = array_index_73956[add_73911 > 32'h0000_0009 ? 4'h9 : add_73911[3:0]] + smul_73960;
  assign array_update_73964[0] = add_73911 == 32'h0000_0000 ? add_73962 : array_index_73956[0];
  assign array_update_73964[1] = add_73911 == 32'h0000_0001 ? add_73962 : array_index_73956[1];
  assign array_update_73964[2] = add_73911 == 32'h0000_0002 ? add_73962 : array_index_73956[2];
  assign array_update_73964[3] = add_73911 == 32'h0000_0003 ? add_73962 : array_index_73956[3];
  assign array_update_73964[4] = add_73911 == 32'h0000_0004 ? add_73962 : array_index_73956[4];
  assign array_update_73964[5] = add_73911 == 32'h0000_0005 ? add_73962 : array_index_73956[5];
  assign array_update_73964[6] = add_73911 == 32'h0000_0006 ? add_73962 : array_index_73956[6];
  assign array_update_73964[7] = add_73911 == 32'h0000_0007 ? add_73962 : array_index_73956[7];
  assign array_update_73964[8] = add_73911 == 32'h0000_0008 ? add_73962 : array_index_73956[8];
  assign array_update_73964[9] = add_73911 == 32'h0000_0009 ? add_73962 : array_index_73956[9];
  assign add_73965 = add_73952 + 32'h0000_0001;
  assign array_update_73966[0] = add_73368 == 32'h0000_0000 ? array_update_73964 : array_update_73953[0];
  assign array_update_73966[1] = add_73368 == 32'h0000_0001 ? array_update_73964 : array_update_73953[1];
  assign array_update_73966[2] = add_73368 == 32'h0000_0002 ? array_update_73964 : array_update_73953[2];
  assign array_update_73966[3] = add_73368 == 32'h0000_0003 ? array_update_73964 : array_update_73953[3];
  assign array_update_73966[4] = add_73368 == 32'h0000_0004 ? array_update_73964 : array_update_73953[4];
  assign array_update_73966[5] = add_73368 == 32'h0000_0005 ? array_update_73964 : array_update_73953[5];
  assign array_update_73966[6] = add_73368 == 32'h0000_0006 ? array_update_73964 : array_update_73953[6];
  assign array_update_73966[7] = add_73368 == 32'h0000_0007 ? array_update_73964 : array_update_73953[7];
  assign array_update_73966[8] = add_73368 == 32'h0000_0008 ? array_update_73964 : array_update_73953[8];
  assign array_update_73966[9] = add_73368 == 32'h0000_0009 ? array_update_73964 : array_update_73953[9];
  assign array_index_73968 = array_update_72021[add_73965 > 32'h0000_0009 ? 4'h9 : add_73965[3:0]];
  assign array_index_73969 = array_update_73966[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_73973 = smul32b_32b_x_32b(array_index_73375[add_73965 > 32'h0000_0009 ? 4'h9 : add_73965[3:0]], array_index_73968[add_73911 > 32'h0000_0009 ? 4'h9 : add_73911[3:0]]);
  assign add_73975 = array_index_73969[add_73911 > 32'h0000_0009 ? 4'h9 : add_73911[3:0]] + smul_73973;
  assign array_update_73977[0] = add_73911 == 32'h0000_0000 ? add_73975 : array_index_73969[0];
  assign array_update_73977[1] = add_73911 == 32'h0000_0001 ? add_73975 : array_index_73969[1];
  assign array_update_73977[2] = add_73911 == 32'h0000_0002 ? add_73975 : array_index_73969[2];
  assign array_update_73977[3] = add_73911 == 32'h0000_0003 ? add_73975 : array_index_73969[3];
  assign array_update_73977[4] = add_73911 == 32'h0000_0004 ? add_73975 : array_index_73969[4];
  assign array_update_73977[5] = add_73911 == 32'h0000_0005 ? add_73975 : array_index_73969[5];
  assign array_update_73977[6] = add_73911 == 32'h0000_0006 ? add_73975 : array_index_73969[6];
  assign array_update_73977[7] = add_73911 == 32'h0000_0007 ? add_73975 : array_index_73969[7];
  assign array_update_73977[8] = add_73911 == 32'h0000_0008 ? add_73975 : array_index_73969[8];
  assign array_update_73977[9] = add_73911 == 32'h0000_0009 ? add_73975 : array_index_73969[9];
  assign add_73978 = add_73965 + 32'h0000_0001;
  assign array_update_73979[0] = add_73368 == 32'h0000_0000 ? array_update_73977 : array_update_73966[0];
  assign array_update_73979[1] = add_73368 == 32'h0000_0001 ? array_update_73977 : array_update_73966[1];
  assign array_update_73979[2] = add_73368 == 32'h0000_0002 ? array_update_73977 : array_update_73966[2];
  assign array_update_73979[3] = add_73368 == 32'h0000_0003 ? array_update_73977 : array_update_73966[3];
  assign array_update_73979[4] = add_73368 == 32'h0000_0004 ? array_update_73977 : array_update_73966[4];
  assign array_update_73979[5] = add_73368 == 32'h0000_0005 ? array_update_73977 : array_update_73966[5];
  assign array_update_73979[6] = add_73368 == 32'h0000_0006 ? array_update_73977 : array_update_73966[6];
  assign array_update_73979[7] = add_73368 == 32'h0000_0007 ? array_update_73977 : array_update_73966[7];
  assign array_update_73979[8] = add_73368 == 32'h0000_0008 ? array_update_73977 : array_update_73966[8];
  assign array_update_73979[9] = add_73368 == 32'h0000_0009 ? array_update_73977 : array_update_73966[9];
  assign array_index_73981 = array_update_72021[add_73978 > 32'h0000_0009 ? 4'h9 : add_73978[3:0]];
  assign array_index_73982 = array_update_73979[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_73986 = smul32b_32b_x_32b(array_index_73375[add_73978 > 32'h0000_0009 ? 4'h9 : add_73978[3:0]], array_index_73981[add_73911 > 32'h0000_0009 ? 4'h9 : add_73911[3:0]]);
  assign add_73988 = array_index_73982[add_73911 > 32'h0000_0009 ? 4'h9 : add_73911[3:0]] + smul_73986;
  assign array_update_73990[0] = add_73911 == 32'h0000_0000 ? add_73988 : array_index_73982[0];
  assign array_update_73990[1] = add_73911 == 32'h0000_0001 ? add_73988 : array_index_73982[1];
  assign array_update_73990[2] = add_73911 == 32'h0000_0002 ? add_73988 : array_index_73982[2];
  assign array_update_73990[3] = add_73911 == 32'h0000_0003 ? add_73988 : array_index_73982[3];
  assign array_update_73990[4] = add_73911 == 32'h0000_0004 ? add_73988 : array_index_73982[4];
  assign array_update_73990[5] = add_73911 == 32'h0000_0005 ? add_73988 : array_index_73982[5];
  assign array_update_73990[6] = add_73911 == 32'h0000_0006 ? add_73988 : array_index_73982[6];
  assign array_update_73990[7] = add_73911 == 32'h0000_0007 ? add_73988 : array_index_73982[7];
  assign array_update_73990[8] = add_73911 == 32'h0000_0008 ? add_73988 : array_index_73982[8];
  assign array_update_73990[9] = add_73911 == 32'h0000_0009 ? add_73988 : array_index_73982[9];
  assign add_73991 = add_73978 + 32'h0000_0001;
  assign array_update_73992[0] = add_73368 == 32'h0000_0000 ? array_update_73990 : array_update_73979[0];
  assign array_update_73992[1] = add_73368 == 32'h0000_0001 ? array_update_73990 : array_update_73979[1];
  assign array_update_73992[2] = add_73368 == 32'h0000_0002 ? array_update_73990 : array_update_73979[2];
  assign array_update_73992[3] = add_73368 == 32'h0000_0003 ? array_update_73990 : array_update_73979[3];
  assign array_update_73992[4] = add_73368 == 32'h0000_0004 ? array_update_73990 : array_update_73979[4];
  assign array_update_73992[5] = add_73368 == 32'h0000_0005 ? array_update_73990 : array_update_73979[5];
  assign array_update_73992[6] = add_73368 == 32'h0000_0006 ? array_update_73990 : array_update_73979[6];
  assign array_update_73992[7] = add_73368 == 32'h0000_0007 ? array_update_73990 : array_update_73979[7];
  assign array_update_73992[8] = add_73368 == 32'h0000_0008 ? array_update_73990 : array_update_73979[8];
  assign array_update_73992[9] = add_73368 == 32'h0000_0009 ? array_update_73990 : array_update_73979[9];
  assign array_index_73994 = array_update_72021[add_73991 > 32'h0000_0009 ? 4'h9 : add_73991[3:0]];
  assign array_index_73995 = array_update_73992[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_73999 = smul32b_32b_x_32b(array_index_73375[add_73991 > 32'h0000_0009 ? 4'h9 : add_73991[3:0]], array_index_73994[add_73911 > 32'h0000_0009 ? 4'h9 : add_73911[3:0]]);
  assign add_74001 = array_index_73995[add_73911 > 32'h0000_0009 ? 4'h9 : add_73911[3:0]] + smul_73999;
  assign array_update_74003[0] = add_73911 == 32'h0000_0000 ? add_74001 : array_index_73995[0];
  assign array_update_74003[1] = add_73911 == 32'h0000_0001 ? add_74001 : array_index_73995[1];
  assign array_update_74003[2] = add_73911 == 32'h0000_0002 ? add_74001 : array_index_73995[2];
  assign array_update_74003[3] = add_73911 == 32'h0000_0003 ? add_74001 : array_index_73995[3];
  assign array_update_74003[4] = add_73911 == 32'h0000_0004 ? add_74001 : array_index_73995[4];
  assign array_update_74003[5] = add_73911 == 32'h0000_0005 ? add_74001 : array_index_73995[5];
  assign array_update_74003[6] = add_73911 == 32'h0000_0006 ? add_74001 : array_index_73995[6];
  assign array_update_74003[7] = add_73911 == 32'h0000_0007 ? add_74001 : array_index_73995[7];
  assign array_update_74003[8] = add_73911 == 32'h0000_0008 ? add_74001 : array_index_73995[8];
  assign array_update_74003[9] = add_73911 == 32'h0000_0009 ? add_74001 : array_index_73995[9];
  assign add_74004 = add_73991 + 32'h0000_0001;
  assign array_update_74005[0] = add_73368 == 32'h0000_0000 ? array_update_74003 : array_update_73992[0];
  assign array_update_74005[1] = add_73368 == 32'h0000_0001 ? array_update_74003 : array_update_73992[1];
  assign array_update_74005[2] = add_73368 == 32'h0000_0002 ? array_update_74003 : array_update_73992[2];
  assign array_update_74005[3] = add_73368 == 32'h0000_0003 ? array_update_74003 : array_update_73992[3];
  assign array_update_74005[4] = add_73368 == 32'h0000_0004 ? array_update_74003 : array_update_73992[4];
  assign array_update_74005[5] = add_73368 == 32'h0000_0005 ? array_update_74003 : array_update_73992[5];
  assign array_update_74005[6] = add_73368 == 32'h0000_0006 ? array_update_74003 : array_update_73992[6];
  assign array_update_74005[7] = add_73368 == 32'h0000_0007 ? array_update_74003 : array_update_73992[7];
  assign array_update_74005[8] = add_73368 == 32'h0000_0008 ? array_update_74003 : array_update_73992[8];
  assign array_update_74005[9] = add_73368 == 32'h0000_0009 ? array_update_74003 : array_update_73992[9];
  assign array_index_74007 = array_update_72021[add_74004 > 32'h0000_0009 ? 4'h9 : add_74004[3:0]];
  assign array_index_74008 = array_update_74005[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_74012 = smul32b_32b_x_32b(array_index_73375[add_74004 > 32'h0000_0009 ? 4'h9 : add_74004[3:0]], array_index_74007[add_73911 > 32'h0000_0009 ? 4'h9 : add_73911[3:0]]);
  assign add_74014 = array_index_74008[add_73911 > 32'h0000_0009 ? 4'h9 : add_73911[3:0]] + smul_74012;
  assign array_update_74016[0] = add_73911 == 32'h0000_0000 ? add_74014 : array_index_74008[0];
  assign array_update_74016[1] = add_73911 == 32'h0000_0001 ? add_74014 : array_index_74008[1];
  assign array_update_74016[2] = add_73911 == 32'h0000_0002 ? add_74014 : array_index_74008[2];
  assign array_update_74016[3] = add_73911 == 32'h0000_0003 ? add_74014 : array_index_74008[3];
  assign array_update_74016[4] = add_73911 == 32'h0000_0004 ? add_74014 : array_index_74008[4];
  assign array_update_74016[5] = add_73911 == 32'h0000_0005 ? add_74014 : array_index_74008[5];
  assign array_update_74016[6] = add_73911 == 32'h0000_0006 ? add_74014 : array_index_74008[6];
  assign array_update_74016[7] = add_73911 == 32'h0000_0007 ? add_74014 : array_index_74008[7];
  assign array_update_74016[8] = add_73911 == 32'h0000_0008 ? add_74014 : array_index_74008[8];
  assign array_update_74016[9] = add_73911 == 32'h0000_0009 ? add_74014 : array_index_74008[9];
  assign add_74017 = add_74004 + 32'h0000_0001;
  assign array_update_74018[0] = add_73368 == 32'h0000_0000 ? array_update_74016 : array_update_74005[0];
  assign array_update_74018[1] = add_73368 == 32'h0000_0001 ? array_update_74016 : array_update_74005[1];
  assign array_update_74018[2] = add_73368 == 32'h0000_0002 ? array_update_74016 : array_update_74005[2];
  assign array_update_74018[3] = add_73368 == 32'h0000_0003 ? array_update_74016 : array_update_74005[3];
  assign array_update_74018[4] = add_73368 == 32'h0000_0004 ? array_update_74016 : array_update_74005[4];
  assign array_update_74018[5] = add_73368 == 32'h0000_0005 ? array_update_74016 : array_update_74005[5];
  assign array_update_74018[6] = add_73368 == 32'h0000_0006 ? array_update_74016 : array_update_74005[6];
  assign array_update_74018[7] = add_73368 == 32'h0000_0007 ? array_update_74016 : array_update_74005[7];
  assign array_update_74018[8] = add_73368 == 32'h0000_0008 ? array_update_74016 : array_update_74005[8];
  assign array_update_74018[9] = add_73368 == 32'h0000_0009 ? array_update_74016 : array_update_74005[9];
  assign array_index_74020 = array_update_72021[add_74017 > 32'h0000_0009 ? 4'h9 : add_74017[3:0]];
  assign array_index_74021 = array_update_74018[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_74025 = smul32b_32b_x_32b(array_index_73375[add_74017 > 32'h0000_0009 ? 4'h9 : add_74017[3:0]], array_index_74020[add_73911 > 32'h0000_0009 ? 4'h9 : add_73911[3:0]]);
  assign add_74027 = array_index_74021[add_73911 > 32'h0000_0009 ? 4'h9 : add_73911[3:0]] + smul_74025;
  assign array_update_74029[0] = add_73911 == 32'h0000_0000 ? add_74027 : array_index_74021[0];
  assign array_update_74029[1] = add_73911 == 32'h0000_0001 ? add_74027 : array_index_74021[1];
  assign array_update_74029[2] = add_73911 == 32'h0000_0002 ? add_74027 : array_index_74021[2];
  assign array_update_74029[3] = add_73911 == 32'h0000_0003 ? add_74027 : array_index_74021[3];
  assign array_update_74029[4] = add_73911 == 32'h0000_0004 ? add_74027 : array_index_74021[4];
  assign array_update_74029[5] = add_73911 == 32'h0000_0005 ? add_74027 : array_index_74021[5];
  assign array_update_74029[6] = add_73911 == 32'h0000_0006 ? add_74027 : array_index_74021[6];
  assign array_update_74029[7] = add_73911 == 32'h0000_0007 ? add_74027 : array_index_74021[7];
  assign array_update_74029[8] = add_73911 == 32'h0000_0008 ? add_74027 : array_index_74021[8];
  assign array_update_74029[9] = add_73911 == 32'h0000_0009 ? add_74027 : array_index_74021[9];
  assign add_74030 = add_74017 + 32'h0000_0001;
  assign array_update_74031[0] = add_73368 == 32'h0000_0000 ? array_update_74029 : array_update_74018[0];
  assign array_update_74031[1] = add_73368 == 32'h0000_0001 ? array_update_74029 : array_update_74018[1];
  assign array_update_74031[2] = add_73368 == 32'h0000_0002 ? array_update_74029 : array_update_74018[2];
  assign array_update_74031[3] = add_73368 == 32'h0000_0003 ? array_update_74029 : array_update_74018[3];
  assign array_update_74031[4] = add_73368 == 32'h0000_0004 ? array_update_74029 : array_update_74018[4];
  assign array_update_74031[5] = add_73368 == 32'h0000_0005 ? array_update_74029 : array_update_74018[5];
  assign array_update_74031[6] = add_73368 == 32'h0000_0006 ? array_update_74029 : array_update_74018[6];
  assign array_update_74031[7] = add_73368 == 32'h0000_0007 ? array_update_74029 : array_update_74018[7];
  assign array_update_74031[8] = add_73368 == 32'h0000_0008 ? array_update_74029 : array_update_74018[8];
  assign array_update_74031[9] = add_73368 == 32'h0000_0009 ? array_update_74029 : array_update_74018[9];
  assign array_index_74033 = array_update_72021[add_74030 > 32'h0000_0009 ? 4'h9 : add_74030[3:0]];
  assign array_index_74034 = array_update_74031[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_74038 = smul32b_32b_x_32b(array_index_73375[add_74030 > 32'h0000_0009 ? 4'h9 : add_74030[3:0]], array_index_74033[add_73911 > 32'h0000_0009 ? 4'h9 : add_73911[3:0]]);
  assign add_74040 = array_index_74034[add_73911 > 32'h0000_0009 ? 4'h9 : add_73911[3:0]] + smul_74038;
  assign array_update_74041[0] = add_73911 == 32'h0000_0000 ? add_74040 : array_index_74034[0];
  assign array_update_74041[1] = add_73911 == 32'h0000_0001 ? add_74040 : array_index_74034[1];
  assign array_update_74041[2] = add_73911 == 32'h0000_0002 ? add_74040 : array_index_74034[2];
  assign array_update_74041[3] = add_73911 == 32'h0000_0003 ? add_74040 : array_index_74034[3];
  assign array_update_74041[4] = add_73911 == 32'h0000_0004 ? add_74040 : array_index_74034[4];
  assign array_update_74041[5] = add_73911 == 32'h0000_0005 ? add_74040 : array_index_74034[5];
  assign array_update_74041[6] = add_73911 == 32'h0000_0006 ? add_74040 : array_index_74034[6];
  assign array_update_74041[7] = add_73911 == 32'h0000_0007 ? add_74040 : array_index_74034[7];
  assign array_update_74041[8] = add_73911 == 32'h0000_0008 ? add_74040 : array_index_74034[8];
  assign array_update_74041[9] = add_73911 == 32'h0000_0009 ? add_74040 : array_index_74034[9];
  assign array_update_74042[0] = add_73368 == 32'h0000_0000 ? array_update_74041 : array_update_74031[0];
  assign array_update_74042[1] = add_73368 == 32'h0000_0001 ? array_update_74041 : array_update_74031[1];
  assign array_update_74042[2] = add_73368 == 32'h0000_0002 ? array_update_74041 : array_update_74031[2];
  assign array_update_74042[3] = add_73368 == 32'h0000_0003 ? array_update_74041 : array_update_74031[3];
  assign array_update_74042[4] = add_73368 == 32'h0000_0004 ? array_update_74041 : array_update_74031[4];
  assign array_update_74042[5] = add_73368 == 32'h0000_0005 ? array_update_74041 : array_update_74031[5];
  assign array_update_74042[6] = add_73368 == 32'h0000_0006 ? array_update_74041 : array_update_74031[6];
  assign array_update_74042[7] = add_73368 == 32'h0000_0007 ? array_update_74041 : array_update_74031[7];
  assign array_update_74042[8] = add_73368 == 32'h0000_0008 ? array_update_74041 : array_update_74031[8];
  assign array_update_74042[9] = add_73368 == 32'h0000_0009 ? array_update_74041 : array_update_74031[9];
  assign array_index_74044 = array_update_74042[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign add_74046 = add_73911 + 32'h0000_0001;
  assign array_update_74047[0] = add_74046 == 32'h0000_0000 ? 32'h0000_0000 : array_index_74044[0];
  assign array_update_74047[1] = add_74046 == 32'h0000_0001 ? 32'h0000_0000 : array_index_74044[1];
  assign array_update_74047[2] = add_74046 == 32'h0000_0002 ? 32'h0000_0000 : array_index_74044[2];
  assign array_update_74047[3] = add_74046 == 32'h0000_0003 ? 32'h0000_0000 : array_index_74044[3];
  assign array_update_74047[4] = add_74046 == 32'h0000_0004 ? 32'h0000_0000 : array_index_74044[4];
  assign array_update_74047[5] = add_74046 == 32'h0000_0005 ? 32'h0000_0000 : array_index_74044[5];
  assign array_update_74047[6] = add_74046 == 32'h0000_0006 ? 32'h0000_0000 : array_index_74044[6];
  assign array_update_74047[7] = add_74046 == 32'h0000_0007 ? 32'h0000_0000 : array_index_74044[7];
  assign array_update_74047[8] = add_74046 == 32'h0000_0008 ? 32'h0000_0000 : array_index_74044[8];
  assign array_update_74047[9] = add_74046 == 32'h0000_0009 ? 32'h0000_0000 : array_index_74044[9];
  assign literal_74048 = 32'h0000_0000;
  assign array_update_74049[0] = add_73368 == 32'h0000_0000 ? array_update_74047 : array_update_74042[0];
  assign array_update_74049[1] = add_73368 == 32'h0000_0001 ? array_update_74047 : array_update_74042[1];
  assign array_update_74049[2] = add_73368 == 32'h0000_0002 ? array_update_74047 : array_update_74042[2];
  assign array_update_74049[3] = add_73368 == 32'h0000_0003 ? array_update_74047 : array_update_74042[3];
  assign array_update_74049[4] = add_73368 == 32'h0000_0004 ? array_update_74047 : array_update_74042[4];
  assign array_update_74049[5] = add_73368 == 32'h0000_0005 ? array_update_74047 : array_update_74042[5];
  assign array_update_74049[6] = add_73368 == 32'h0000_0006 ? array_update_74047 : array_update_74042[6];
  assign array_update_74049[7] = add_73368 == 32'h0000_0007 ? array_update_74047 : array_update_74042[7];
  assign array_update_74049[8] = add_73368 == 32'h0000_0008 ? array_update_74047 : array_update_74042[8];
  assign array_update_74049[9] = add_73368 == 32'h0000_0009 ? array_update_74047 : array_update_74042[9];
  assign array_index_74051 = array_update_72021[literal_74048 > 32'h0000_0009 ? 4'h9 : literal_74048[3:0]];
  assign array_index_74052 = array_update_74049[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_74056 = smul32b_32b_x_32b(array_index_73375[literal_74048 > 32'h0000_0009 ? 4'h9 : literal_74048[3:0]], array_index_74051[add_74046 > 32'h0000_0009 ? 4'h9 : add_74046[3:0]]);
  assign add_74058 = array_index_74052[add_74046 > 32'h0000_0009 ? 4'h9 : add_74046[3:0]] + smul_74056;
  assign array_update_74060[0] = add_74046 == 32'h0000_0000 ? add_74058 : array_index_74052[0];
  assign array_update_74060[1] = add_74046 == 32'h0000_0001 ? add_74058 : array_index_74052[1];
  assign array_update_74060[2] = add_74046 == 32'h0000_0002 ? add_74058 : array_index_74052[2];
  assign array_update_74060[3] = add_74046 == 32'h0000_0003 ? add_74058 : array_index_74052[3];
  assign array_update_74060[4] = add_74046 == 32'h0000_0004 ? add_74058 : array_index_74052[4];
  assign array_update_74060[5] = add_74046 == 32'h0000_0005 ? add_74058 : array_index_74052[5];
  assign array_update_74060[6] = add_74046 == 32'h0000_0006 ? add_74058 : array_index_74052[6];
  assign array_update_74060[7] = add_74046 == 32'h0000_0007 ? add_74058 : array_index_74052[7];
  assign array_update_74060[8] = add_74046 == 32'h0000_0008 ? add_74058 : array_index_74052[8];
  assign array_update_74060[9] = add_74046 == 32'h0000_0009 ? add_74058 : array_index_74052[9];
  assign add_74061 = literal_74048 + 32'h0000_0001;
  assign array_update_74062[0] = add_73368 == 32'h0000_0000 ? array_update_74060 : array_update_74049[0];
  assign array_update_74062[1] = add_73368 == 32'h0000_0001 ? array_update_74060 : array_update_74049[1];
  assign array_update_74062[2] = add_73368 == 32'h0000_0002 ? array_update_74060 : array_update_74049[2];
  assign array_update_74062[3] = add_73368 == 32'h0000_0003 ? array_update_74060 : array_update_74049[3];
  assign array_update_74062[4] = add_73368 == 32'h0000_0004 ? array_update_74060 : array_update_74049[4];
  assign array_update_74062[5] = add_73368 == 32'h0000_0005 ? array_update_74060 : array_update_74049[5];
  assign array_update_74062[6] = add_73368 == 32'h0000_0006 ? array_update_74060 : array_update_74049[6];
  assign array_update_74062[7] = add_73368 == 32'h0000_0007 ? array_update_74060 : array_update_74049[7];
  assign array_update_74062[8] = add_73368 == 32'h0000_0008 ? array_update_74060 : array_update_74049[8];
  assign array_update_74062[9] = add_73368 == 32'h0000_0009 ? array_update_74060 : array_update_74049[9];
  assign array_index_74064 = array_update_72021[add_74061 > 32'h0000_0009 ? 4'h9 : add_74061[3:0]];
  assign array_index_74065 = array_update_74062[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_74069 = smul32b_32b_x_32b(array_index_73375[add_74061 > 32'h0000_0009 ? 4'h9 : add_74061[3:0]], array_index_74064[add_74046 > 32'h0000_0009 ? 4'h9 : add_74046[3:0]]);
  assign add_74071 = array_index_74065[add_74046 > 32'h0000_0009 ? 4'h9 : add_74046[3:0]] + smul_74069;
  assign array_update_74073[0] = add_74046 == 32'h0000_0000 ? add_74071 : array_index_74065[0];
  assign array_update_74073[1] = add_74046 == 32'h0000_0001 ? add_74071 : array_index_74065[1];
  assign array_update_74073[2] = add_74046 == 32'h0000_0002 ? add_74071 : array_index_74065[2];
  assign array_update_74073[3] = add_74046 == 32'h0000_0003 ? add_74071 : array_index_74065[3];
  assign array_update_74073[4] = add_74046 == 32'h0000_0004 ? add_74071 : array_index_74065[4];
  assign array_update_74073[5] = add_74046 == 32'h0000_0005 ? add_74071 : array_index_74065[5];
  assign array_update_74073[6] = add_74046 == 32'h0000_0006 ? add_74071 : array_index_74065[6];
  assign array_update_74073[7] = add_74046 == 32'h0000_0007 ? add_74071 : array_index_74065[7];
  assign array_update_74073[8] = add_74046 == 32'h0000_0008 ? add_74071 : array_index_74065[8];
  assign array_update_74073[9] = add_74046 == 32'h0000_0009 ? add_74071 : array_index_74065[9];
  assign add_74074 = add_74061 + 32'h0000_0001;
  assign array_update_74075[0] = add_73368 == 32'h0000_0000 ? array_update_74073 : array_update_74062[0];
  assign array_update_74075[1] = add_73368 == 32'h0000_0001 ? array_update_74073 : array_update_74062[1];
  assign array_update_74075[2] = add_73368 == 32'h0000_0002 ? array_update_74073 : array_update_74062[2];
  assign array_update_74075[3] = add_73368 == 32'h0000_0003 ? array_update_74073 : array_update_74062[3];
  assign array_update_74075[4] = add_73368 == 32'h0000_0004 ? array_update_74073 : array_update_74062[4];
  assign array_update_74075[5] = add_73368 == 32'h0000_0005 ? array_update_74073 : array_update_74062[5];
  assign array_update_74075[6] = add_73368 == 32'h0000_0006 ? array_update_74073 : array_update_74062[6];
  assign array_update_74075[7] = add_73368 == 32'h0000_0007 ? array_update_74073 : array_update_74062[7];
  assign array_update_74075[8] = add_73368 == 32'h0000_0008 ? array_update_74073 : array_update_74062[8];
  assign array_update_74075[9] = add_73368 == 32'h0000_0009 ? array_update_74073 : array_update_74062[9];
  assign array_index_74077 = array_update_72021[add_74074 > 32'h0000_0009 ? 4'h9 : add_74074[3:0]];
  assign array_index_74078 = array_update_74075[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_74082 = smul32b_32b_x_32b(array_index_73375[add_74074 > 32'h0000_0009 ? 4'h9 : add_74074[3:0]], array_index_74077[add_74046 > 32'h0000_0009 ? 4'h9 : add_74046[3:0]]);
  assign add_74084 = array_index_74078[add_74046 > 32'h0000_0009 ? 4'h9 : add_74046[3:0]] + smul_74082;
  assign array_update_74086[0] = add_74046 == 32'h0000_0000 ? add_74084 : array_index_74078[0];
  assign array_update_74086[1] = add_74046 == 32'h0000_0001 ? add_74084 : array_index_74078[1];
  assign array_update_74086[2] = add_74046 == 32'h0000_0002 ? add_74084 : array_index_74078[2];
  assign array_update_74086[3] = add_74046 == 32'h0000_0003 ? add_74084 : array_index_74078[3];
  assign array_update_74086[4] = add_74046 == 32'h0000_0004 ? add_74084 : array_index_74078[4];
  assign array_update_74086[5] = add_74046 == 32'h0000_0005 ? add_74084 : array_index_74078[5];
  assign array_update_74086[6] = add_74046 == 32'h0000_0006 ? add_74084 : array_index_74078[6];
  assign array_update_74086[7] = add_74046 == 32'h0000_0007 ? add_74084 : array_index_74078[7];
  assign array_update_74086[8] = add_74046 == 32'h0000_0008 ? add_74084 : array_index_74078[8];
  assign array_update_74086[9] = add_74046 == 32'h0000_0009 ? add_74084 : array_index_74078[9];
  assign add_74087 = add_74074 + 32'h0000_0001;
  assign array_update_74088[0] = add_73368 == 32'h0000_0000 ? array_update_74086 : array_update_74075[0];
  assign array_update_74088[1] = add_73368 == 32'h0000_0001 ? array_update_74086 : array_update_74075[1];
  assign array_update_74088[2] = add_73368 == 32'h0000_0002 ? array_update_74086 : array_update_74075[2];
  assign array_update_74088[3] = add_73368 == 32'h0000_0003 ? array_update_74086 : array_update_74075[3];
  assign array_update_74088[4] = add_73368 == 32'h0000_0004 ? array_update_74086 : array_update_74075[4];
  assign array_update_74088[5] = add_73368 == 32'h0000_0005 ? array_update_74086 : array_update_74075[5];
  assign array_update_74088[6] = add_73368 == 32'h0000_0006 ? array_update_74086 : array_update_74075[6];
  assign array_update_74088[7] = add_73368 == 32'h0000_0007 ? array_update_74086 : array_update_74075[7];
  assign array_update_74088[8] = add_73368 == 32'h0000_0008 ? array_update_74086 : array_update_74075[8];
  assign array_update_74088[9] = add_73368 == 32'h0000_0009 ? array_update_74086 : array_update_74075[9];
  assign array_index_74090 = array_update_72021[add_74087 > 32'h0000_0009 ? 4'h9 : add_74087[3:0]];
  assign array_index_74091 = array_update_74088[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_74095 = smul32b_32b_x_32b(array_index_73375[add_74087 > 32'h0000_0009 ? 4'h9 : add_74087[3:0]], array_index_74090[add_74046 > 32'h0000_0009 ? 4'h9 : add_74046[3:0]]);
  assign add_74097 = array_index_74091[add_74046 > 32'h0000_0009 ? 4'h9 : add_74046[3:0]] + smul_74095;
  assign array_update_74099[0] = add_74046 == 32'h0000_0000 ? add_74097 : array_index_74091[0];
  assign array_update_74099[1] = add_74046 == 32'h0000_0001 ? add_74097 : array_index_74091[1];
  assign array_update_74099[2] = add_74046 == 32'h0000_0002 ? add_74097 : array_index_74091[2];
  assign array_update_74099[3] = add_74046 == 32'h0000_0003 ? add_74097 : array_index_74091[3];
  assign array_update_74099[4] = add_74046 == 32'h0000_0004 ? add_74097 : array_index_74091[4];
  assign array_update_74099[5] = add_74046 == 32'h0000_0005 ? add_74097 : array_index_74091[5];
  assign array_update_74099[6] = add_74046 == 32'h0000_0006 ? add_74097 : array_index_74091[6];
  assign array_update_74099[7] = add_74046 == 32'h0000_0007 ? add_74097 : array_index_74091[7];
  assign array_update_74099[8] = add_74046 == 32'h0000_0008 ? add_74097 : array_index_74091[8];
  assign array_update_74099[9] = add_74046 == 32'h0000_0009 ? add_74097 : array_index_74091[9];
  assign add_74100 = add_74087 + 32'h0000_0001;
  assign array_update_74101[0] = add_73368 == 32'h0000_0000 ? array_update_74099 : array_update_74088[0];
  assign array_update_74101[1] = add_73368 == 32'h0000_0001 ? array_update_74099 : array_update_74088[1];
  assign array_update_74101[2] = add_73368 == 32'h0000_0002 ? array_update_74099 : array_update_74088[2];
  assign array_update_74101[3] = add_73368 == 32'h0000_0003 ? array_update_74099 : array_update_74088[3];
  assign array_update_74101[4] = add_73368 == 32'h0000_0004 ? array_update_74099 : array_update_74088[4];
  assign array_update_74101[5] = add_73368 == 32'h0000_0005 ? array_update_74099 : array_update_74088[5];
  assign array_update_74101[6] = add_73368 == 32'h0000_0006 ? array_update_74099 : array_update_74088[6];
  assign array_update_74101[7] = add_73368 == 32'h0000_0007 ? array_update_74099 : array_update_74088[7];
  assign array_update_74101[8] = add_73368 == 32'h0000_0008 ? array_update_74099 : array_update_74088[8];
  assign array_update_74101[9] = add_73368 == 32'h0000_0009 ? array_update_74099 : array_update_74088[9];
  assign array_index_74103 = array_update_72021[add_74100 > 32'h0000_0009 ? 4'h9 : add_74100[3:0]];
  assign array_index_74104 = array_update_74101[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_74108 = smul32b_32b_x_32b(array_index_73375[add_74100 > 32'h0000_0009 ? 4'h9 : add_74100[3:0]], array_index_74103[add_74046 > 32'h0000_0009 ? 4'h9 : add_74046[3:0]]);
  assign add_74110 = array_index_74104[add_74046 > 32'h0000_0009 ? 4'h9 : add_74046[3:0]] + smul_74108;
  assign array_update_74112[0] = add_74046 == 32'h0000_0000 ? add_74110 : array_index_74104[0];
  assign array_update_74112[1] = add_74046 == 32'h0000_0001 ? add_74110 : array_index_74104[1];
  assign array_update_74112[2] = add_74046 == 32'h0000_0002 ? add_74110 : array_index_74104[2];
  assign array_update_74112[3] = add_74046 == 32'h0000_0003 ? add_74110 : array_index_74104[3];
  assign array_update_74112[4] = add_74046 == 32'h0000_0004 ? add_74110 : array_index_74104[4];
  assign array_update_74112[5] = add_74046 == 32'h0000_0005 ? add_74110 : array_index_74104[5];
  assign array_update_74112[6] = add_74046 == 32'h0000_0006 ? add_74110 : array_index_74104[6];
  assign array_update_74112[7] = add_74046 == 32'h0000_0007 ? add_74110 : array_index_74104[7];
  assign array_update_74112[8] = add_74046 == 32'h0000_0008 ? add_74110 : array_index_74104[8];
  assign array_update_74112[9] = add_74046 == 32'h0000_0009 ? add_74110 : array_index_74104[9];
  assign add_74113 = add_74100 + 32'h0000_0001;
  assign array_update_74114[0] = add_73368 == 32'h0000_0000 ? array_update_74112 : array_update_74101[0];
  assign array_update_74114[1] = add_73368 == 32'h0000_0001 ? array_update_74112 : array_update_74101[1];
  assign array_update_74114[2] = add_73368 == 32'h0000_0002 ? array_update_74112 : array_update_74101[2];
  assign array_update_74114[3] = add_73368 == 32'h0000_0003 ? array_update_74112 : array_update_74101[3];
  assign array_update_74114[4] = add_73368 == 32'h0000_0004 ? array_update_74112 : array_update_74101[4];
  assign array_update_74114[5] = add_73368 == 32'h0000_0005 ? array_update_74112 : array_update_74101[5];
  assign array_update_74114[6] = add_73368 == 32'h0000_0006 ? array_update_74112 : array_update_74101[6];
  assign array_update_74114[7] = add_73368 == 32'h0000_0007 ? array_update_74112 : array_update_74101[7];
  assign array_update_74114[8] = add_73368 == 32'h0000_0008 ? array_update_74112 : array_update_74101[8];
  assign array_update_74114[9] = add_73368 == 32'h0000_0009 ? array_update_74112 : array_update_74101[9];
  assign array_index_74116 = array_update_72021[add_74113 > 32'h0000_0009 ? 4'h9 : add_74113[3:0]];
  assign array_index_74117 = array_update_74114[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_74121 = smul32b_32b_x_32b(array_index_73375[add_74113 > 32'h0000_0009 ? 4'h9 : add_74113[3:0]], array_index_74116[add_74046 > 32'h0000_0009 ? 4'h9 : add_74046[3:0]]);
  assign add_74123 = array_index_74117[add_74046 > 32'h0000_0009 ? 4'h9 : add_74046[3:0]] + smul_74121;
  assign array_update_74125[0] = add_74046 == 32'h0000_0000 ? add_74123 : array_index_74117[0];
  assign array_update_74125[1] = add_74046 == 32'h0000_0001 ? add_74123 : array_index_74117[1];
  assign array_update_74125[2] = add_74046 == 32'h0000_0002 ? add_74123 : array_index_74117[2];
  assign array_update_74125[3] = add_74046 == 32'h0000_0003 ? add_74123 : array_index_74117[3];
  assign array_update_74125[4] = add_74046 == 32'h0000_0004 ? add_74123 : array_index_74117[4];
  assign array_update_74125[5] = add_74046 == 32'h0000_0005 ? add_74123 : array_index_74117[5];
  assign array_update_74125[6] = add_74046 == 32'h0000_0006 ? add_74123 : array_index_74117[6];
  assign array_update_74125[7] = add_74046 == 32'h0000_0007 ? add_74123 : array_index_74117[7];
  assign array_update_74125[8] = add_74046 == 32'h0000_0008 ? add_74123 : array_index_74117[8];
  assign array_update_74125[9] = add_74046 == 32'h0000_0009 ? add_74123 : array_index_74117[9];
  assign add_74126 = add_74113 + 32'h0000_0001;
  assign array_update_74127[0] = add_73368 == 32'h0000_0000 ? array_update_74125 : array_update_74114[0];
  assign array_update_74127[1] = add_73368 == 32'h0000_0001 ? array_update_74125 : array_update_74114[1];
  assign array_update_74127[2] = add_73368 == 32'h0000_0002 ? array_update_74125 : array_update_74114[2];
  assign array_update_74127[3] = add_73368 == 32'h0000_0003 ? array_update_74125 : array_update_74114[3];
  assign array_update_74127[4] = add_73368 == 32'h0000_0004 ? array_update_74125 : array_update_74114[4];
  assign array_update_74127[5] = add_73368 == 32'h0000_0005 ? array_update_74125 : array_update_74114[5];
  assign array_update_74127[6] = add_73368 == 32'h0000_0006 ? array_update_74125 : array_update_74114[6];
  assign array_update_74127[7] = add_73368 == 32'h0000_0007 ? array_update_74125 : array_update_74114[7];
  assign array_update_74127[8] = add_73368 == 32'h0000_0008 ? array_update_74125 : array_update_74114[8];
  assign array_update_74127[9] = add_73368 == 32'h0000_0009 ? array_update_74125 : array_update_74114[9];
  assign array_index_74129 = array_update_72021[add_74126 > 32'h0000_0009 ? 4'h9 : add_74126[3:0]];
  assign array_index_74130 = array_update_74127[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_74134 = smul32b_32b_x_32b(array_index_73375[add_74126 > 32'h0000_0009 ? 4'h9 : add_74126[3:0]], array_index_74129[add_74046 > 32'h0000_0009 ? 4'h9 : add_74046[3:0]]);
  assign add_74136 = array_index_74130[add_74046 > 32'h0000_0009 ? 4'h9 : add_74046[3:0]] + smul_74134;
  assign array_update_74138[0] = add_74046 == 32'h0000_0000 ? add_74136 : array_index_74130[0];
  assign array_update_74138[1] = add_74046 == 32'h0000_0001 ? add_74136 : array_index_74130[1];
  assign array_update_74138[2] = add_74046 == 32'h0000_0002 ? add_74136 : array_index_74130[2];
  assign array_update_74138[3] = add_74046 == 32'h0000_0003 ? add_74136 : array_index_74130[3];
  assign array_update_74138[4] = add_74046 == 32'h0000_0004 ? add_74136 : array_index_74130[4];
  assign array_update_74138[5] = add_74046 == 32'h0000_0005 ? add_74136 : array_index_74130[5];
  assign array_update_74138[6] = add_74046 == 32'h0000_0006 ? add_74136 : array_index_74130[6];
  assign array_update_74138[7] = add_74046 == 32'h0000_0007 ? add_74136 : array_index_74130[7];
  assign array_update_74138[8] = add_74046 == 32'h0000_0008 ? add_74136 : array_index_74130[8];
  assign array_update_74138[9] = add_74046 == 32'h0000_0009 ? add_74136 : array_index_74130[9];
  assign add_74139 = add_74126 + 32'h0000_0001;
  assign array_update_74140[0] = add_73368 == 32'h0000_0000 ? array_update_74138 : array_update_74127[0];
  assign array_update_74140[1] = add_73368 == 32'h0000_0001 ? array_update_74138 : array_update_74127[1];
  assign array_update_74140[2] = add_73368 == 32'h0000_0002 ? array_update_74138 : array_update_74127[2];
  assign array_update_74140[3] = add_73368 == 32'h0000_0003 ? array_update_74138 : array_update_74127[3];
  assign array_update_74140[4] = add_73368 == 32'h0000_0004 ? array_update_74138 : array_update_74127[4];
  assign array_update_74140[5] = add_73368 == 32'h0000_0005 ? array_update_74138 : array_update_74127[5];
  assign array_update_74140[6] = add_73368 == 32'h0000_0006 ? array_update_74138 : array_update_74127[6];
  assign array_update_74140[7] = add_73368 == 32'h0000_0007 ? array_update_74138 : array_update_74127[7];
  assign array_update_74140[8] = add_73368 == 32'h0000_0008 ? array_update_74138 : array_update_74127[8];
  assign array_update_74140[9] = add_73368 == 32'h0000_0009 ? array_update_74138 : array_update_74127[9];
  assign array_index_74142 = array_update_72021[add_74139 > 32'h0000_0009 ? 4'h9 : add_74139[3:0]];
  assign array_index_74143 = array_update_74140[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_74147 = smul32b_32b_x_32b(array_index_73375[add_74139 > 32'h0000_0009 ? 4'h9 : add_74139[3:0]], array_index_74142[add_74046 > 32'h0000_0009 ? 4'h9 : add_74046[3:0]]);
  assign add_74149 = array_index_74143[add_74046 > 32'h0000_0009 ? 4'h9 : add_74046[3:0]] + smul_74147;
  assign array_update_74151[0] = add_74046 == 32'h0000_0000 ? add_74149 : array_index_74143[0];
  assign array_update_74151[1] = add_74046 == 32'h0000_0001 ? add_74149 : array_index_74143[1];
  assign array_update_74151[2] = add_74046 == 32'h0000_0002 ? add_74149 : array_index_74143[2];
  assign array_update_74151[3] = add_74046 == 32'h0000_0003 ? add_74149 : array_index_74143[3];
  assign array_update_74151[4] = add_74046 == 32'h0000_0004 ? add_74149 : array_index_74143[4];
  assign array_update_74151[5] = add_74046 == 32'h0000_0005 ? add_74149 : array_index_74143[5];
  assign array_update_74151[6] = add_74046 == 32'h0000_0006 ? add_74149 : array_index_74143[6];
  assign array_update_74151[7] = add_74046 == 32'h0000_0007 ? add_74149 : array_index_74143[7];
  assign array_update_74151[8] = add_74046 == 32'h0000_0008 ? add_74149 : array_index_74143[8];
  assign array_update_74151[9] = add_74046 == 32'h0000_0009 ? add_74149 : array_index_74143[9];
  assign add_74152 = add_74139 + 32'h0000_0001;
  assign array_update_74153[0] = add_73368 == 32'h0000_0000 ? array_update_74151 : array_update_74140[0];
  assign array_update_74153[1] = add_73368 == 32'h0000_0001 ? array_update_74151 : array_update_74140[1];
  assign array_update_74153[2] = add_73368 == 32'h0000_0002 ? array_update_74151 : array_update_74140[2];
  assign array_update_74153[3] = add_73368 == 32'h0000_0003 ? array_update_74151 : array_update_74140[3];
  assign array_update_74153[4] = add_73368 == 32'h0000_0004 ? array_update_74151 : array_update_74140[4];
  assign array_update_74153[5] = add_73368 == 32'h0000_0005 ? array_update_74151 : array_update_74140[5];
  assign array_update_74153[6] = add_73368 == 32'h0000_0006 ? array_update_74151 : array_update_74140[6];
  assign array_update_74153[7] = add_73368 == 32'h0000_0007 ? array_update_74151 : array_update_74140[7];
  assign array_update_74153[8] = add_73368 == 32'h0000_0008 ? array_update_74151 : array_update_74140[8];
  assign array_update_74153[9] = add_73368 == 32'h0000_0009 ? array_update_74151 : array_update_74140[9];
  assign array_index_74155 = array_update_72021[add_74152 > 32'h0000_0009 ? 4'h9 : add_74152[3:0]];
  assign array_index_74156 = array_update_74153[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_74160 = smul32b_32b_x_32b(array_index_73375[add_74152 > 32'h0000_0009 ? 4'h9 : add_74152[3:0]], array_index_74155[add_74046 > 32'h0000_0009 ? 4'h9 : add_74046[3:0]]);
  assign add_74162 = array_index_74156[add_74046 > 32'h0000_0009 ? 4'h9 : add_74046[3:0]] + smul_74160;
  assign array_update_74164[0] = add_74046 == 32'h0000_0000 ? add_74162 : array_index_74156[0];
  assign array_update_74164[1] = add_74046 == 32'h0000_0001 ? add_74162 : array_index_74156[1];
  assign array_update_74164[2] = add_74046 == 32'h0000_0002 ? add_74162 : array_index_74156[2];
  assign array_update_74164[3] = add_74046 == 32'h0000_0003 ? add_74162 : array_index_74156[3];
  assign array_update_74164[4] = add_74046 == 32'h0000_0004 ? add_74162 : array_index_74156[4];
  assign array_update_74164[5] = add_74046 == 32'h0000_0005 ? add_74162 : array_index_74156[5];
  assign array_update_74164[6] = add_74046 == 32'h0000_0006 ? add_74162 : array_index_74156[6];
  assign array_update_74164[7] = add_74046 == 32'h0000_0007 ? add_74162 : array_index_74156[7];
  assign array_update_74164[8] = add_74046 == 32'h0000_0008 ? add_74162 : array_index_74156[8];
  assign array_update_74164[9] = add_74046 == 32'h0000_0009 ? add_74162 : array_index_74156[9];
  assign add_74165 = add_74152 + 32'h0000_0001;
  assign array_update_74166[0] = add_73368 == 32'h0000_0000 ? array_update_74164 : array_update_74153[0];
  assign array_update_74166[1] = add_73368 == 32'h0000_0001 ? array_update_74164 : array_update_74153[1];
  assign array_update_74166[2] = add_73368 == 32'h0000_0002 ? array_update_74164 : array_update_74153[2];
  assign array_update_74166[3] = add_73368 == 32'h0000_0003 ? array_update_74164 : array_update_74153[3];
  assign array_update_74166[4] = add_73368 == 32'h0000_0004 ? array_update_74164 : array_update_74153[4];
  assign array_update_74166[5] = add_73368 == 32'h0000_0005 ? array_update_74164 : array_update_74153[5];
  assign array_update_74166[6] = add_73368 == 32'h0000_0006 ? array_update_74164 : array_update_74153[6];
  assign array_update_74166[7] = add_73368 == 32'h0000_0007 ? array_update_74164 : array_update_74153[7];
  assign array_update_74166[8] = add_73368 == 32'h0000_0008 ? array_update_74164 : array_update_74153[8];
  assign array_update_74166[9] = add_73368 == 32'h0000_0009 ? array_update_74164 : array_update_74153[9];
  assign array_index_74168 = array_update_72021[add_74165 > 32'h0000_0009 ? 4'h9 : add_74165[3:0]];
  assign array_index_74169 = array_update_74166[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_74173 = smul32b_32b_x_32b(array_index_73375[add_74165 > 32'h0000_0009 ? 4'h9 : add_74165[3:0]], array_index_74168[add_74046 > 32'h0000_0009 ? 4'h9 : add_74046[3:0]]);
  assign add_74175 = array_index_74169[add_74046 > 32'h0000_0009 ? 4'h9 : add_74046[3:0]] + smul_74173;
  assign array_update_74176[0] = add_74046 == 32'h0000_0000 ? add_74175 : array_index_74169[0];
  assign array_update_74176[1] = add_74046 == 32'h0000_0001 ? add_74175 : array_index_74169[1];
  assign array_update_74176[2] = add_74046 == 32'h0000_0002 ? add_74175 : array_index_74169[2];
  assign array_update_74176[3] = add_74046 == 32'h0000_0003 ? add_74175 : array_index_74169[3];
  assign array_update_74176[4] = add_74046 == 32'h0000_0004 ? add_74175 : array_index_74169[4];
  assign array_update_74176[5] = add_74046 == 32'h0000_0005 ? add_74175 : array_index_74169[5];
  assign array_update_74176[6] = add_74046 == 32'h0000_0006 ? add_74175 : array_index_74169[6];
  assign array_update_74176[7] = add_74046 == 32'h0000_0007 ? add_74175 : array_index_74169[7];
  assign array_update_74176[8] = add_74046 == 32'h0000_0008 ? add_74175 : array_index_74169[8];
  assign array_update_74176[9] = add_74046 == 32'h0000_0009 ? add_74175 : array_index_74169[9];
  assign array_update_74177[0] = add_73368 == 32'h0000_0000 ? array_update_74176 : array_update_74166[0];
  assign array_update_74177[1] = add_73368 == 32'h0000_0001 ? array_update_74176 : array_update_74166[1];
  assign array_update_74177[2] = add_73368 == 32'h0000_0002 ? array_update_74176 : array_update_74166[2];
  assign array_update_74177[3] = add_73368 == 32'h0000_0003 ? array_update_74176 : array_update_74166[3];
  assign array_update_74177[4] = add_73368 == 32'h0000_0004 ? array_update_74176 : array_update_74166[4];
  assign array_update_74177[5] = add_73368 == 32'h0000_0005 ? array_update_74176 : array_update_74166[5];
  assign array_update_74177[6] = add_73368 == 32'h0000_0006 ? array_update_74176 : array_update_74166[6];
  assign array_update_74177[7] = add_73368 == 32'h0000_0007 ? array_update_74176 : array_update_74166[7];
  assign array_update_74177[8] = add_73368 == 32'h0000_0008 ? array_update_74176 : array_update_74166[8];
  assign array_update_74177[9] = add_73368 == 32'h0000_0009 ? array_update_74176 : array_update_74166[9];
  assign array_index_74179 = array_update_74177[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign add_74181 = add_74046 + 32'h0000_0001;
  assign array_update_74182[0] = add_74181 == 32'h0000_0000 ? 32'h0000_0000 : array_index_74179[0];
  assign array_update_74182[1] = add_74181 == 32'h0000_0001 ? 32'h0000_0000 : array_index_74179[1];
  assign array_update_74182[2] = add_74181 == 32'h0000_0002 ? 32'h0000_0000 : array_index_74179[2];
  assign array_update_74182[3] = add_74181 == 32'h0000_0003 ? 32'h0000_0000 : array_index_74179[3];
  assign array_update_74182[4] = add_74181 == 32'h0000_0004 ? 32'h0000_0000 : array_index_74179[4];
  assign array_update_74182[5] = add_74181 == 32'h0000_0005 ? 32'h0000_0000 : array_index_74179[5];
  assign array_update_74182[6] = add_74181 == 32'h0000_0006 ? 32'h0000_0000 : array_index_74179[6];
  assign array_update_74182[7] = add_74181 == 32'h0000_0007 ? 32'h0000_0000 : array_index_74179[7];
  assign array_update_74182[8] = add_74181 == 32'h0000_0008 ? 32'h0000_0000 : array_index_74179[8];
  assign array_update_74182[9] = add_74181 == 32'h0000_0009 ? 32'h0000_0000 : array_index_74179[9];
  assign literal_74183 = 32'h0000_0000;
  assign array_update_74184[0] = add_73368 == 32'h0000_0000 ? array_update_74182 : array_update_74177[0];
  assign array_update_74184[1] = add_73368 == 32'h0000_0001 ? array_update_74182 : array_update_74177[1];
  assign array_update_74184[2] = add_73368 == 32'h0000_0002 ? array_update_74182 : array_update_74177[2];
  assign array_update_74184[3] = add_73368 == 32'h0000_0003 ? array_update_74182 : array_update_74177[3];
  assign array_update_74184[4] = add_73368 == 32'h0000_0004 ? array_update_74182 : array_update_74177[4];
  assign array_update_74184[5] = add_73368 == 32'h0000_0005 ? array_update_74182 : array_update_74177[5];
  assign array_update_74184[6] = add_73368 == 32'h0000_0006 ? array_update_74182 : array_update_74177[6];
  assign array_update_74184[7] = add_73368 == 32'h0000_0007 ? array_update_74182 : array_update_74177[7];
  assign array_update_74184[8] = add_73368 == 32'h0000_0008 ? array_update_74182 : array_update_74177[8];
  assign array_update_74184[9] = add_73368 == 32'h0000_0009 ? array_update_74182 : array_update_74177[9];
  assign array_index_74186 = array_update_72021[literal_74183 > 32'h0000_0009 ? 4'h9 : literal_74183[3:0]];
  assign array_index_74187 = array_update_74184[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_74191 = smul32b_32b_x_32b(array_index_73375[literal_74183 > 32'h0000_0009 ? 4'h9 : literal_74183[3:0]], array_index_74186[add_74181 > 32'h0000_0009 ? 4'h9 : add_74181[3:0]]);
  assign add_74193 = array_index_74187[add_74181 > 32'h0000_0009 ? 4'h9 : add_74181[3:0]] + smul_74191;
  assign array_update_74195[0] = add_74181 == 32'h0000_0000 ? add_74193 : array_index_74187[0];
  assign array_update_74195[1] = add_74181 == 32'h0000_0001 ? add_74193 : array_index_74187[1];
  assign array_update_74195[2] = add_74181 == 32'h0000_0002 ? add_74193 : array_index_74187[2];
  assign array_update_74195[3] = add_74181 == 32'h0000_0003 ? add_74193 : array_index_74187[3];
  assign array_update_74195[4] = add_74181 == 32'h0000_0004 ? add_74193 : array_index_74187[4];
  assign array_update_74195[5] = add_74181 == 32'h0000_0005 ? add_74193 : array_index_74187[5];
  assign array_update_74195[6] = add_74181 == 32'h0000_0006 ? add_74193 : array_index_74187[6];
  assign array_update_74195[7] = add_74181 == 32'h0000_0007 ? add_74193 : array_index_74187[7];
  assign array_update_74195[8] = add_74181 == 32'h0000_0008 ? add_74193 : array_index_74187[8];
  assign array_update_74195[9] = add_74181 == 32'h0000_0009 ? add_74193 : array_index_74187[9];
  assign add_74196 = literal_74183 + 32'h0000_0001;
  assign array_update_74197[0] = add_73368 == 32'h0000_0000 ? array_update_74195 : array_update_74184[0];
  assign array_update_74197[1] = add_73368 == 32'h0000_0001 ? array_update_74195 : array_update_74184[1];
  assign array_update_74197[2] = add_73368 == 32'h0000_0002 ? array_update_74195 : array_update_74184[2];
  assign array_update_74197[3] = add_73368 == 32'h0000_0003 ? array_update_74195 : array_update_74184[3];
  assign array_update_74197[4] = add_73368 == 32'h0000_0004 ? array_update_74195 : array_update_74184[4];
  assign array_update_74197[5] = add_73368 == 32'h0000_0005 ? array_update_74195 : array_update_74184[5];
  assign array_update_74197[6] = add_73368 == 32'h0000_0006 ? array_update_74195 : array_update_74184[6];
  assign array_update_74197[7] = add_73368 == 32'h0000_0007 ? array_update_74195 : array_update_74184[7];
  assign array_update_74197[8] = add_73368 == 32'h0000_0008 ? array_update_74195 : array_update_74184[8];
  assign array_update_74197[9] = add_73368 == 32'h0000_0009 ? array_update_74195 : array_update_74184[9];
  assign array_index_74199 = array_update_72021[add_74196 > 32'h0000_0009 ? 4'h9 : add_74196[3:0]];
  assign array_index_74200 = array_update_74197[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_74204 = smul32b_32b_x_32b(array_index_73375[add_74196 > 32'h0000_0009 ? 4'h9 : add_74196[3:0]], array_index_74199[add_74181 > 32'h0000_0009 ? 4'h9 : add_74181[3:0]]);
  assign add_74206 = array_index_74200[add_74181 > 32'h0000_0009 ? 4'h9 : add_74181[3:0]] + smul_74204;
  assign array_update_74208[0] = add_74181 == 32'h0000_0000 ? add_74206 : array_index_74200[0];
  assign array_update_74208[1] = add_74181 == 32'h0000_0001 ? add_74206 : array_index_74200[1];
  assign array_update_74208[2] = add_74181 == 32'h0000_0002 ? add_74206 : array_index_74200[2];
  assign array_update_74208[3] = add_74181 == 32'h0000_0003 ? add_74206 : array_index_74200[3];
  assign array_update_74208[4] = add_74181 == 32'h0000_0004 ? add_74206 : array_index_74200[4];
  assign array_update_74208[5] = add_74181 == 32'h0000_0005 ? add_74206 : array_index_74200[5];
  assign array_update_74208[6] = add_74181 == 32'h0000_0006 ? add_74206 : array_index_74200[6];
  assign array_update_74208[7] = add_74181 == 32'h0000_0007 ? add_74206 : array_index_74200[7];
  assign array_update_74208[8] = add_74181 == 32'h0000_0008 ? add_74206 : array_index_74200[8];
  assign array_update_74208[9] = add_74181 == 32'h0000_0009 ? add_74206 : array_index_74200[9];
  assign add_74209 = add_74196 + 32'h0000_0001;
  assign array_update_74210[0] = add_73368 == 32'h0000_0000 ? array_update_74208 : array_update_74197[0];
  assign array_update_74210[1] = add_73368 == 32'h0000_0001 ? array_update_74208 : array_update_74197[1];
  assign array_update_74210[2] = add_73368 == 32'h0000_0002 ? array_update_74208 : array_update_74197[2];
  assign array_update_74210[3] = add_73368 == 32'h0000_0003 ? array_update_74208 : array_update_74197[3];
  assign array_update_74210[4] = add_73368 == 32'h0000_0004 ? array_update_74208 : array_update_74197[4];
  assign array_update_74210[5] = add_73368 == 32'h0000_0005 ? array_update_74208 : array_update_74197[5];
  assign array_update_74210[6] = add_73368 == 32'h0000_0006 ? array_update_74208 : array_update_74197[6];
  assign array_update_74210[7] = add_73368 == 32'h0000_0007 ? array_update_74208 : array_update_74197[7];
  assign array_update_74210[8] = add_73368 == 32'h0000_0008 ? array_update_74208 : array_update_74197[8];
  assign array_update_74210[9] = add_73368 == 32'h0000_0009 ? array_update_74208 : array_update_74197[9];
  assign array_index_74212 = array_update_72021[add_74209 > 32'h0000_0009 ? 4'h9 : add_74209[3:0]];
  assign array_index_74213 = array_update_74210[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_74217 = smul32b_32b_x_32b(array_index_73375[add_74209 > 32'h0000_0009 ? 4'h9 : add_74209[3:0]], array_index_74212[add_74181 > 32'h0000_0009 ? 4'h9 : add_74181[3:0]]);
  assign add_74219 = array_index_74213[add_74181 > 32'h0000_0009 ? 4'h9 : add_74181[3:0]] + smul_74217;
  assign array_update_74221[0] = add_74181 == 32'h0000_0000 ? add_74219 : array_index_74213[0];
  assign array_update_74221[1] = add_74181 == 32'h0000_0001 ? add_74219 : array_index_74213[1];
  assign array_update_74221[2] = add_74181 == 32'h0000_0002 ? add_74219 : array_index_74213[2];
  assign array_update_74221[3] = add_74181 == 32'h0000_0003 ? add_74219 : array_index_74213[3];
  assign array_update_74221[4] = add_74181 == 32'h0000_0004 ? add_74219 : array_index_74213[4];
  assign array_update_74221[5] = add_74181 == 32'h0000_0005 ? add_74219 : array_index_74213[5];
  assign array_update_74221[6] = add_74181 == 32'h0000_0006 ? add_74219 : array_index_74213[6];
  assign array_update_74221[7] = add_74181 == 32'h0000_0007 ? add_74219 : array_index_74213[7];
  assign array_update_74221[8] = add_74181 == 32'h0000_0008 ? add_74219 : array_index_74213[8];
  assign array_update_74221[9] = add_74181 == 32'h0000_0009 ? add_74219 : array_index_74213[9];
  assign add_74222 = add_74209 + 32'h0000_0001;
  assign array_update_74223[0] = add_73368 == 32'h0000_0000 ? array_update_74221 : array_update_74210[0];
  assign array_update_74223[1] = add_73368 == 32'h0000_0001 ? array_update_74221 : array_update_74210[1];
  assign array_update_74223[2] = add_73368 == 32'h0000_0002 ? array_update_74221 : array_update_74210[2];
  assign array_update_74223[3] = add_73368 == 32'h0000_0003 ? array_update_74221 : array_update_74210[3];
  assign array_update_74223[4] = add_73368 == 32'h0000_0004 ? array_update_74221 : array_update_74210[4];
  assign array_update_74223[5] = add_73368 == 32'h0000_0005 ? array_update_74221 : array_update_74210[5];
  assign array_update_74223[6] = add_73368 == 32'h0000_0006 ? array_update_74221 : array_update_74210[6];
  assign array_update_74223[7] = add_73368 == 32'h0000_0007 ? array_update_74221 : array_update_74210[7];
  assign array_update_74223[8] = add_73368 == 32'h0000_0008 ? array_update_74221 : array_update_74210[8];
  assign array_update_74223[9] = add_73368 == 32'h0000_0009 ? array_update_74221 : array_update_74210[9];
  assign array_index_74225 = array_update_72021[add_74222 > 32'h0000_0009 ? 4'h9 : add_74222[3:0]];
  assign array_index_74226 = array_update_74223[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_74230 = smul32b_32b_x_32b(array_index_73375[add_74222 > 32'h0000_0009 ? 4'h9 : add_74222[3:0]], array_index_74225[add_74181 > 32'h0000_0009 ? 4'h9 : add_74181[3:0]]);
  assign add_74232 = array_index_74226[add_74181 > 32'h0000_0009 ? 4'h9 : add_74181[3:0]] + smul_74230;
  assign array_update_74234[0] = add_74181 == 32'h0000_0000 ? add_74232 : array_index_74226[0];
  assign array_update_74234[1] = add_74181 == 32'h0000_0001 ? add_74232 : array_index_74226[1];
  assign array_update_74234[2] = add_74181 == 32'h0000_0002 ? add_74232 : array_index_74226[2];
  assign array_update_74234[3] = add_74181 == 32'h0000_0003 ? add_74232 : array_index_74226[3];
  assign array_update_74234[4] = add_74181 == 32'h0000_0004 ? add_74232 : array_index_74226[4];
  assign array_update_74234[5] = add_74181 == 32'h0000_0005 ? add_74232 : array_index_74226[5];
  assign array_update_74234[6] = add_74181 == 32'h0000_0006 ? add_74232 : array_index_74226[6];
  assign array_update_74234[7] = add_74181 == 32'h0000_0007 ? add_74232 : array_index_74226[7];
  assign array_update_74234[8] = add_74181 == 32'h0000_0008 ? add_74232 : array_index_74226[8];
  assign array_update_74234[9] = add_74181 == 32'h0000_0009 ? add_74232 : array_index_74226[9];
  assign add_74235 = add_74222 + 32'h0000_0001;
  assign array_update_74236[0] = add_73368 == 32'h0000_0000 ? array_update_74234 : array_update_74223[0];
  assign array_update_74236[1] = add_73368 == 32'h0000_0001 ? array_update_74234 : array_update_74223[1];
  assign array_update_74236[2] = add_73368 == 32'h0000_0002 ? array_update_74234 : array_update_74223[2];
  assign array_update_74236[3] = add_73368 == 32'h0000_0003 ? array_update_74234 : array_update_74223[3];
  assign array_update_74236[4] = add_73368 == 32'h0000_0004 ? array_update_74234 : array_update_74223[4];
  assign array_update_74236[5] = add_73368 == 32'h0000_0005 ? array_update_74234 : array_update_74223[5];
  assign array_update_74236[6] = add_73368 == 32'h0000_0006 ? array_update_74234 : array_update_74223[6];
  assign array_update_74236[7] = add_73368 == 32'h0000_0007 ? array_update_74234 : array_update_74223[7];
  assign array_update_74236[8] = add_73368 == 32'h0000_0008 ? array_update_74234 : array_update_74223[8];
  assign array_update_74236[9] = add_73368 == 32'h0000_0009 ? array_update_74234 : array_update_74223[9];
  assign array_index_74238 = array_update_72021[add_74235 > 32'h0000_0009 ? 4'h9 : add_74235[3:0]];
  assign array_index_74239 = array_update_74236[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_74243 = smul32b_32b_x_32b(array_index_73375[add_74235 > 32'h0000_0009 ? 4'h9 : add_74235[3:0]], array_index_74238[add_74181 > 32'h0000_0009 ? 4'h9 : add_74181[3:0]]);
  assign add_74245 = array_index_74239[add_74181 > 32'h0000_0009 ? 4'h9 : add_74181[3:0]] + smul_74243;
  assign array_update_74247[0] = add_74181 == 32'h0000_0000 ? add_74245 : array_index_74239[0];
  assign array_update_74247[1] = add_74181 == 32'h0000_0001 ? add_74245 : array_index_74239[1];
  assign array_update_74247[2] = add_74181 == 32'h0000_0002 ? add_74245 : array_index_74239[2];
  assign array_update_74247[3] = add_74181 == 32'h0000_0003 ? add_74245 : array_index_74239[3];
  assign array_update_74247[4] = add_74181 == 32'h0000_0004 ? add_74245 : array_index_74239[4];
  assign array_update_74247[5] = add_74181 == 32'h0000_0005 ? add_74245 : array_index_74239[5];
  assign array_update_74247[6] = add_74181 == 32'h0000_0006 ? add_74245 : array_index_74239[6];
  assign array_update_74247[7] = add_74181 == 32'h0000_0007 ? add_74245 : array_index_74239[7];
  assign array_update_74247[8] = add_74181 == 32'h0000_0008 ? add_74245 : array_index_74239[8];
  assign array_update_74247[9] = add_74181 == 32'h0000_0009 ? add_74245 : array_index_74239[9];
  assign add_74248 = add_74235 + 32'h0000_0001;
  assign array_update_74249[0] = add_73368 == 32'h0000_0000 ? array_update_74247 : array_update_74236[0];
  assign array_update_74249[1] = add_73368 == 32'h0000_0001 ? array_update_74247 : array_update_74236[1];
  assign array_update_74249[2] = add_73368 == 32'h0000_0002 ? array_update_74247 : array_update_74236[2];
  assign array_update_74249[3] = add_73368 == 32'h0000_0003 ? array_update_74247 : array_update_74236[3];
  assign array_update_74249[4] = add_73368 == 32'h0000_0004 ? array_update_74247 : array_update_74236[4];
  assign array_update_74249[5] = add_73368 == 32'h0000_0005 ? array_update_74247 : array_update_74236[5];
  assign array_update_74249[6] = add_73368 == 32'h0000_0006 ? array_update_74247 : array_update_74236[6];
  assign array_update_74249[7] = add_73368 == 32'h0000_0007 ? array_update_74247 : array_update_74236[7];
  assign array_update_74249[8] = add_73368 == 32'h0000_0008 ? array_update_74247 : array_update_74236[8];
  assign array_update_74249[9] = add_73368 == 32'h0000_0009 ? array_update_74247 : array_update_74236[9];
  assign array_index_74251 = array_update_72021[add_74248 > 32'h0000_0009 ? 4'h9 : add_74248[3:0]];
  assign array_index_74252 = array_update_74249[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_74256 = smul32b_32b_x_32b(array_index_73375[add_74248 > 32'h0000_0009 ? 4'h9 : add_74248[3:0]], array_index_74251[add_74181 > 32'h0000_0009 ? 4'h9 : add_74181[3:0]]);
  assign add_74258 = array_index_74252[add_74181 > 32'h0000_0009 ? 4'h9 : add_74181[3:0]] + smul_74256;
  assign array_update_74260[0] = add_74181 == 32'h0000_0000 ? add_74258 : array_index_74252[0];
  assign array_update_74260[1] = add_74181 == 32'h0000_0001 ? add_74258 : array_index_74252[1];
  assign array_update_74260[2] = add_74181 == 32'h0000_0002 ? add_74258 : array_index_74252[2];
  assign array_update_74260[3] = add_74181 == 32'h0000_0003 ? add_74258 : array_index_74252[3];
  assign array_update_74260[4] = add_74181 == 32'h0000_0004 ? add_74258 : array_index_74252[4];
  assign array_update_74260[5] = add_74181 == 32'h0000_0005 ? add_74258 : array_index_74252[5];
  assign array_update_74260[6] = add_74181 == 32'h0000_0006 ? add_74258 : array_index_74252[6];
  assign array_update_74260[7] = add_74181 == 32'h0000_0007 ? add_74258 : array_index_74252[7];
  assign array_update_74260[8] = add_74181 == 32'h0000_0008 ? add_74258 : array_index_74252[8];
  assign array_update_74260[9] = add_74181 == 32'h0000_0009 ? add_74258 : array_index_74252[9];
  assign add_74261 = add_74248 + 32'h0000_0001;
  assign array_update_74262[0] = add_73368 == 32'h0000_0000 ? array_update_74260 : array_update_74249[0];
  assign array_update_74262[1] = add_73368 == 32'h0000_0001 ? array_update_74260 : array_update_74249[1];
  assign array_update_74262[2] = add_73368 == 32'h0000_0002 ? array_update_74260 : array_update_74249[2];
  assign array_update_74262[3] = add_73368 == 32'h0000_0003 ? array_update_74260 : array_update_74249[3];
  assign array_update_74262[4] = add_73368 == 32'h0000_0004 ? array_update_74260 : array_update_74249[4];
  assign array_update_74262[5] = add_73368 == 32'h0000_0005 ? array_update_74260 : array_update_74249[5];
  assign array_update_74262[6] = add_73368 == 32'h0000_0006 ? array_update_74260 : array_update_74249[6];
  assign array_update_74262[7] = add_73368 == 32'h0000_0007 ? array_update_74260 : array_update_74249[7];
  assign array_update_74262[8] = add_73368 == 32'h0000_0008 ? array_update_74260 : array_update_74249[8];
  assign array_update_74262[9] = add_73368 == 32'h0000_0009 ? array_update_74260 : array_update_74249[9];
  assign array_index_74264 = array_update_72021[add_74261 > 32'h0000_0009 ? 4'h9 : add_74261[3:0]];
  assign array_index_74265 = array_update_74262[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_74269 = smul32b_32b_x_32b(array_index_73375[add_74261 > 32'h0000_0009 ? 4'h9 : add_74261[3:0]], array_index_74264[add_74181 > 32'h0000_0009 ? 4'h9 : add_74181[3:0]]);
  assign add_74271 = array_index_74265[add_74181 > 32'h0000_0009 ? 4'h9 : add_74181[3:0]] + smul_74269;
  assign array_update_74273[0] = add_74181 == 32'h0000_0000 ? add_74271 : array_index_74265[0];
  assign array_update_74273[1] = add_74181 == 32'h0000_0001 ? add_74271 : array_index_74265[1];
  assign array_update_74273[2] = add_74181 == 32'h0000_0002 ? add_74271 : array_index_74265[2];
  assign array_update_74273[3] = add_74181 == 32'h0000_0003 ? add_74271 : array_index_74265[3];
  assign array_update_74273[4] = add_74181 == 32'h0000_0004 ? add_74271 : array_index_74265[4];
  assign array_update_74273[5] = add_74181 == 32'h0000_0005 ? add_74271 : array_index_74265[5];
  assign array_update_74273[6] = add_74181 == 32'h0000_0006 ? add_74271 : array_index_74265[6];
  assign array_update_74273[7] = add_74181 == 32'h0000_0007 ? add_74271 : array_index_74265[7];
  assign array_update_74273[8] = add_74181 == 32'h0000_0008 ? add_74271 : array_index_74265[8];
  assign array_update_74273[9] = add_74181 == 32'h0000_0009 ? add_74271 : array_index_74265[9];
  assign add_74274 = add_74261 + 32'h0000_0001;
  assign array_update_74275[0] = add_73368 == 32'h0000_0000 ? array_update_74273 : array_update_74262[0];
  assign array_update_74275[1] = add_73368 == 32'h0000_0001 ? array_update_74273 : array_update_74262[1];
  assign array_update_74275[2] = add_73368 == 32'h0000_0002 ? array_update_74273 : array_update_74262[2];
  assign array_update_74275[3] = add_73368 == 32'h0000_0003 ? array_update_74273 : array_update_74262[3];
  assign array_update_74275[4] = add_73368 == 32'h0000_0004 ? array_update_74273 : array_update_74262[4];
  assign array_update_74275[5] = add_73368 == 32'h0000_0005 ? array_update_74273 : array_update_74262[5];
  assign array_update_74275[6] = add_73368 == 32'h0000_0006 ? array_update_74273 : array_update_74262[6];
  assign array_update_74275[7] = add_73368 == 32'h0000_0007 ? array_update_74273 : array_update_74262[7];
  assign array_update_74275[8] = add_73368 == 32'h0000_0008 ? array_update_74273 : array_update_74262[8];
  assign array_update_74275[9] = add_73368 == 32'h0000_0009 ? array_update_74273 : array_update_74262[9];
  assign array_index_74277 = array_update_72021[add_74274 > 32'h0000_0009 ? 4'h9 : add_74274[3:0]];
  assign array_index_74278 = array_update_74275[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_74282 = smul32b_32b_x_32b(array_index_73375[add_74274 > 32'h0000_0009 ? 4'h9 : add_74274[3:0]], array_index_74277[add_74181 > 32'h0000_0009 ? 4'h9 : add_74181[3:0]]);
  assign add_74284 = array_index_74278[add_74181 > 32'h0000_0009 ? 4'h9 : add_74181[3:0]] + smul_74282;
  assign array_update_74286[0] = add_74181 == 32'h0000_0000 ? add_74284 : array_index_74278[0];
  assign array_update_74286[1] = add_74181 == 32'h0000_0001 ? add_74284 : array_index_74278[1];
  assign array_update_74286[2] = add_74181 == 32'h0000_0002 ? add_74284 : array_index_74278[2];
  assign array_update_74286[3] = add_74181 == 32'h0000_0003 ? add_74284 : array_index_74278[3];
  assign array_update_74286[4] = add_74181 == 32'h0000_0004 ? add_74284 : array_index_74278[4];
  assign array_update_74286[5] = add_74181 == 32'h0000_0005 ? add_74284 : array_index_74278[5];
  assign array_update_74286[6] = add_74181 == 32'h0000_0006 ? add_74284 : array_index_74278[6];
  assign array_update_74286[7] = add_74181 == 32'h0000_0007 ? add_74284 : array_index_74278[7];
  assign array_update_74286[8] = add_74181 == 32'h0000_0008 ? add_74284 : array_index_74278[8];
  assign array_update_74286[9] = add_74181 == 32'h0000_0009 ? add_74284 : array_index_74278[9];
  assign add_74287 = add_74274 + 32'h0000_0001;
  assign array_update_74288[0] = add_73368 == 32'h0000_0000 ? array_update_74286 : array_update_74275[0];
  assign array_update_74288[1] = add_73368 == 32'h0000_0001 ? array_update_74286 : array_update_74275[1];
  assign array_update_74288[2] = add_73368 == 32'h0000_0002 ? array_update_74286 : array_update_74275[2];
  assign array_update_74288[3] = add_73368 == 32'h0000_0003 ? array_update_74286 : array_update_74275[3];
  assign array_update_74288[4] = add_73368 == 32'h0000_0004 ? array_update_74286 : array_update_74275[4];
  assign array_update_74288[5] = add_73368 == 32'h0000_0005 ? array_update_74286 : array_update_74275[5];
  assign array_update_74288[6] = add_73368 == 32'h0000_0006 ? array_update_74286 : array_update_74275[6];
  assign array_update_74288[7] = add_73368 == 32'h0000_0007 ? array_update_74286 : array_update_74275[7];
  assign array_update_74288[8] = add_73368 == 32'h0000_0008 ? array_update_74286 : array_update_74275[8];
  assign array_update_74288[9] = add_73368 == 32'h0000_0009 ? array_update_74286 : array_update_74275[9];
  assign array_index_74290 = array_update_72021[add_74287 > 32'h0000_0009 ? 4'h9 : add_74287[3:0]];
  assign array_index_74291 = array_update_74288[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_74295 = smul32b_32b_x_32b(array_index_73375[add_74287 > 32'h0000_0009 ? 4'h9 : add_74287[3:0]], array_index_74290[add_74181 > 32'h0000_0009 ? 4'h9 : add_74181[3:0]]);
  assign add_74297 = array_index_74291[add_74181 > 32'h0000_0009 ? 4'h9 : add_74181[3:0]] + smul_74295;
  assign array_update_74299[0] = add_74181 == 32'h0000_0000 ? add_74297 : array_index_74291[0];
  assign array_update_74299[1] = add_74181 == 32'h0000_0001 ? add_74297 : array_index_74291[1];
  assign array_update_74299[2] = add_74181 == 32'h0000_0002 ? add_74297 : array_index_74291[2];
  assign array_update_74299[3] = add_74181 == 32'h0000_0003 ? add_74297 : array_index_74291[3];
  assign array_update_74299[4] = add_74181 == 32'h0000_0004 ? add_74297 : array_index_74291[4];
  assign array_update_74299[5] = add_74181 == 32'h0000_0005 ? add_74297 : array_index_74291[5];
  assign array_update_74299[6] = add_74181 == 32'h0000_0006 ? add_74297 : array_index_74291[6];
  assign array_update_74299[7] = add_74181 == 32'h0000_0007 ? add_74297 : array_index_74291[7];
  assign array_update_74299[8] = add_74181 == 32'h0000_0008 ? add_74297 : array_index_74291[8];
  assign array_update_74299[9] = add_74181 == 32'h0000_0009 ? add_74297 : array_index_74291[9];
  assign add_74300 = add_74287 + 32'h0000_0001;
  assign array_update_74301[0] = add_73368 == 32'h0000_0000 ? array_update_74299 : array_update_74288[0];
  assign array_update_74301[1] = add_73368 == 32'h0000_0001 ? array_update_74299 : array_update_74288[1];
  assign array_update_74301[2] = add_73368 == 32'h0000_0002 ? array_update_74299 : array_update_74288[2];
  assign array_update_74301[3] = add_73368 == 32'h0000_0003 ? array_update_74299 : array_update_74288[3];
  assign array_update_74301[4] = add_73368 == 32'h0000_0004 ? array_update_74299 : array_update_74288[4];
  assign array_update_74301[5] = add_73368 == 32'h0000_0005 ? array_update_74299 : array_update_74288[5];
  assign array_update_74301[6] = add_73368 == 32'h0000_0006 ? array_update_74299 : array_update_74288[6];
  assign array_update_74301[7] = add_73368 == 32'h0000_0007 ? array_update_74299 : array_update_74288[7];
  assign array_update_74301[8] = add_73368 == 32'h0000_0008 ? array_update_74299 : array_update_74288[8];
  assign array_update_74301[9] = add_73368 == 32'h0000_0009 ? array_update_74299 : array_update_74288[9];
  assign array_index_74303 = array_update_72021[add_74300 > 32'h0000_0009 ? 4'h9 : add_74300[3:0]];
  assign array_index_74304 = array_update_74301[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_74308 = smul32b_32b_x_32b(array_index_73375[add_74300 > 32'h0000_0009 ? 4'h9 : add_74300[3:0]], array_index_74303[add_74181 > 32'h0000_0009 ? 4'h9 : add_74181[3:0]]);
  assign add_74310 = array_index_74304[add_74181 > 32'h0000_0009 ? 4'h9 : add_74181[3:0]] + smul_74308;
  assign array_update_74311[0] = add_74181 == 32'h0000_0000 ? add_74310 : array_index_74304[0];
  assign array_update_74311[1] = add_74181 == 32'h0000_0001 ? add_74310 : array_index_74304[1];
  assign array_update_74311[2] = add_74181 == 32'h0000_0002 ? add_74310 : array_index_74304[2];
  assign array_update_74311[3] = add_74181 == 32'h0000_0003 ? add_74310 : array_index_74304[3];
  assign array_update_74311[4] = add_74181 == 32'h0000_0004 ? add_74310 : array_index_74304[4];
  assign array_update_74311[5] = add_74181 == 32'h0000_0005 ? add_74310 : array_index_74304[5];
  assign array_update_74311[6] = add_74181 == 32'h0000_0006 ? add_74310 : array_index_74304[6];
  assign array_update_74311[7] = add_74181 == 32'h0000_0007 ? add_74310 : array_index_74304[7];
  assign array_update_74311[8] = add_74181 == 32'h0000_0008 ? add_74310 : array_index_74304[8];
  assign array_update_74311[9] = add_74181 == 32'h0000_0009 ? add_74310 : array_index_74304[9];
  assign array_update_74312[0] = add_73368 == 32'h0000_0000 ? array_update_74311 : array_update_74301[0];
  assign array_update_74312[1] = add_73368 == 32'h0000_0001 ? array_update_74311 : array_update_74301[1];
  assign array_update_74312[2] = add_73368 == 32'h0000_0002 ? array_update_74311 : array_update_74301[2];
  assign array_update_74312[3] = add_73368 == 32'h0000_0003 ? array_update_74311 : array_update_74301[3];
  assign array_update_74312[4] = add_73368 == 32'h0000_0004 ? array_update_74311 : array_update_74301[4];
  assign array_update_74312[5] = add_73368 == 32'h0000_0005 ? array_update_74311 : array_update_74301[5];
  assign array_update_74312[6] = add_73368 == 32'h0000_0006 ? array_update_74311 : array_update_74301[6];
  assign array_update_74312[7] = add_73368 == 32'h0000_0007 ? array_update_74311 : array_update_74301[7];
  assign array_update_74312[8] = add_73368 == 32'h0000_0008 ? array_update_74311 : array_update_74301[8];
  assign array_update_74312[9] = add_73368 == 32'h0000_0009 ? array_update_74311 : array_update_74301[9];
  assign array_index_74314 = array_update_74312[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign add_74316 = add_74181 + 32'h0000_0001;
  assign array_update_74317[0] = add_74316 == 32'h0000_0000 ? 32'h0000_0000 : array_index_74314[0];
  assign array_update_74317[1] = add_74316 == 32'h0000_0001 ? 32'h0000_0000 : array_index_74314[1];
  assign array_update_74317[2] = add_74316 == 32'h0000_0002 ? 32'h0000_0000 : array_index_74314[2];
  assign array_update_74317[3] = add_74316 == 32'h0000_0003 ? 32'h0000_0000 : array_index_74314[3];
  assign array_update_74317[4] = add_74316 == 32'h0000_0004 ? 32'h0000_0000 : array_index_74314[4];
  assign array_update_74317[5] = add_74316 == 32'h0000_0005 ? 32'h0000_0000 : array_index_74314[5];
  assign array_update_74317[6] = add_74316 == 32'h0000_0006 ? 32'h0000_0000 : array_index_74314[6];
  assign array_update_74317[7] = add_74316 == 32'h0000_0007 ? 32'h0000_0000 : array_index_74314[7];
  assign array_update_74317[8] = add_74316 == 32'h0000_0008 ? 32'h0000_0000 : array_index_74314[8];
  assign array_update_74317[9] = add_74316 == 32'h0000_0009 ? 32'h0000_0000 : array_index_74314[9];
  assign literal_74318 = 32'h0000_0000;
  assign array_update_74319[0] = add_73368 == 32'h0000_0000 ? array_update_74317 : array_update_74312[0];
  assign array_update_74319[1] = add_73368 == 32'h0000_0001 ? array_update_74317 : array_update_74312[1];
  assign array_update_74319[2] = add_73368 == 32'h0000_0002 ? array_update_74317 : array_update_74312[2];
  assign array_update_74319[3] = add_73368 == 32'h0000_0003 ? array_update_74317 : array_update_74312[3];
  assign array_update_74319[4] = add_73368 == 32'h0000_0004 ? array_update_74317 : array_update_74312[4];
  assign array_update_74319[5] = add_73368 == 32'h0000_0005 ? array_update_74317 : array_update_74312[5];
  assign array_update_74319[6] = add_73368 == 32'h0000_0006 ? array_update_74317 : array_update_74312[6];
  assign array_update_74319[7] = add_73368 == 32'h0000_0007 ? array_update_74317 : array_update_74312[7];
  assign array_update_74319[8] = add_73368 == 32'h0000_0008 ? array_update_74317 : array_update_74312[8];
  assign array_update_74319[9] = add_73368 == 32'h0000_0009 ? array_update_74317 : array_update_74312[9];
  assign array_index_74321 = array_update_72021[literal_74318 > 32'h0000_0009 ? 4'h9 : literal_74318[3:0]];
  assign array_index_74322 = array_update_74319[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_74326 = smul32b_32b_x_32b(array_index_73375[literal_74318 > 32'h0000_0009 ? 4'h9 : literal_74318[3:0]], array_index_74321[add_74316 > 32'h0000_0009 ? 4'h9 : add_74316[3:0]]);
  assign add_74328 = array_index_74322[add_74316 > 32'h0000_0009 ? 4'h9 : add_74316[3:0]] + smul_74326;
  assign array_update_74330[0] = add_74316 == 32'h0000_0000 ? add_74328 : array_index_74322[0];
  assign array_update_74330[1] = add_74316 == 32'h0000_0001 ? add_74328 : array_index_74322[1];
  assign array_update_74330[2] = add_74316 == 32'h0000_0002 ? add_74328 : array_index_74322[2];
  assign array_update_74330[3] = add_74316 == 32'h0000_0003 ? add_74328 : array_index_74322[3];
  assign array_update_74330[4] = add_74316 == 32'h0000_0004 ? add_74328 : array_index_74322[4];
  assign array_update_74330[5] = add_74316 == 32'h0000_0005 ? add_74328 : array_index_74322[5];
  assign array_update_74330[6] = add_74316 == 32'h0000_0006 ? add_74328 : array_index_74322[6];
  assign array_update_74330[7] = add_74316 == 32'h0000_0007 ? add_74328 : array_index_74322[7];
  assign array_update_74330[8] = add_74316 == 32'h0000_0008 ? add_74328 : array_index_74322[8];
  assign array_update_74330[9] = add_74316 == 32'h0000_0009 ? add_74328 : array_index_74322[9];
  assign add_74331 = literal_74318 + 32'h0000_0001;
  assign array_update_74332[0] = add_73368 == 32'h0000_0000 ? array_update_74330 : array_update_74319[0];
  assign array_update_74332[1] = add_73368 == 32'h0000_0001 ? array_update_74330 : array_update_74319[1];
  assign array_update_74332[2] = add_73368 == 32'h0000_0002 ? array_update_74330 : array_update_74319[2];
  assign array_update_74332[3] = add_73368 == 32'h0000_0003 ? array_update_74330 : array_update_74319[3];
  assign array_update_74332[4] = add_73368 == 32'h0000_0004 ? array_update_74330 : array_update_74319[4];
  assign array_update_74332[5] = add_73368 == 32'h0000_0005 ? array_update_74330 : array_update_74319[5];
  assign array_update_74332[6] = add_73368 == 32'h0000_0006 ? array_update_74330 : array_update_74319[6];
  assign array_update_74332[7] = add_73368 == 32'h0000_0007 ? array_update_74330 : array_update_74319[7];
  assign array_update_74332[8] = add_73368 == 32'h0000_0008 ? array_update_74330 : array_update_74319[8];
  assign array_update_74332[9] = add_73368 == 32'h0000_0009 ? array_update_74330 : array_update_74319[9];
  assign array_index_74334 = array_update_72021[add_74331 > 32'h0000_0009 ? 4'h9 : add_74331[3:0]];
  assign array_index_74335 = array_update_74332[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_74339 = smul32b_32b_x_32b(array_index_73375[add_74331 > 32'h0000_0009 ? 4'h9 : add_74331[3:0]], array_index_74334[add_74316 > 32'h0000_0009 ? 4'h9 : add_74316[3:0]]);
  assign add_74341 = array_index_74335[add_74316 > 32'h0000_0009 ? 4'h9 : add_74316[3:0]] + smul_74339;
  assign array_update_74343[0] = add_74316 == 32'h0000_0000 ? add_74341 : array_index_74335[0];
  assign array_update_74343[1] = add_74316 == 32'h0000_0001 ? add_74341 : array_index_74335[1];
  assign array_update_74343[2] = add_74316 == 32'h0000_0002 ? add_74341 : array_index_74335[2];
  assign array_update_74343[3] = add_74316 == 32'h0000_0003 ? add_74341 : array_index_74335[3];
  assign array_update_74343[4] = add_74316 == 32'h0000_0004 ? add_74341 : array_index_74335[4];
  assign array_update_74343[5] = add_74316 == 32'h0000_0005 ? add_74341 : array_index_74335[5];
  assign array_update_74343[6] = add_74316 == 32'h0000_0006 ? add_74341 : array_index_74335[6];
  assign array_update_74343[7] = add_74316 == 32'h0000_0007 ? add_74341 : array_index_74335[7];
  assign array_update_74343[8] = add_74316 == 32'h0000_0008 ? add_74341 : array_index_74335[8];
  assign array_update_74343[9] = add_74316 == 32'h0000_0009 ? add_74341 : array_index_74335[9];
  assign add_74344 = add_74331 + 32'h0000_0001;
  assign array_update_74345[0] = add_73368 == 32'h0000_0000 ? array_update_74343 : array_update_74332[0];
  assign array_update_74345[1] = add_73368 == 32'h0000_0001 ? array_update_74343 : array_update_74332[1];
  assign array_update_74345[2] = add_73368 == 32'h0000_0002 ? array_update_74343 : array_update_74332[2];
  assign array_update_74345[3] = add_73368 == 32'h0000_0003 ? array_update_74343 : array_update_74332[3];
  assign array_update_74345[4] = add_73368 == 32'h0000_0004 ? array_update_74343 : array_update_74332[4];
  assign array_update_74345[5] = add_73368 == 32'h0000_0005 ? array_update_74343 : array_update_74332[5];
  assign array_update_74345[6] = add_73368 == 32'h0000_0006 ? array_update_74343 : array_update_74332[6];
  assign array_update_74345[7] = add_73368 == 32'h0000_0007 ? array_update_74343 : array_update_74332[7];
  assign array_update_74345[8] = add_73368 == 32'h0000_0008 ? array_update_74343 : array_update_74332[8];
  assign array_update_74345[9] = add_73368 == 32'h0000_0009 ? array_update_74343 : array_update_74332[9];
  assign array_index_74347 = array_update_72021[add_74344 > 32'h0000_0009 ? 4'h9 : add_74344[3:0]];
  assign array_index_74348 = array_update_74345[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_74352 = smul32b_32b_x_32b(array_index_73375[add_74344 > 32'h0000_0009 ? 4'h9 : add_74344[3:0]], array_index_74347[add_74316 > 32'h0000_0009 ? 4'h9 : add_74316[3:0]]);
  assign add_74354 = array_index_74348[add_74316 > 32'h0000_0009 ? 4'h9 : add_74316[3:0]] + smul_74352;
  assign array_update_74356[0] = add_74316 == 32'h0000_0000 ? add_74354 : array_index_74348[0];
  assign array_update_74356[1] = add_74316 == 32'h0000_0001 ? add_74354 : array_index_74348[1];
  assign array_update_74356[2] = add_74316 == 32'h0000_0002 ? add_74354 : array_index_74348[2];
  assign array_update_74356[3] = add_74316 == 32'h0000_0003 ? add_74354 : array_index_74348[3];
  assign array_update_74356[4] = add_74316 == 32'h0000_0004 ? add_74354 : array_index_74348[4];
  assign array_update_74356[5] = add_74316 == 32'h0000_0005 ? add_74354 : array_index_74348[5];
  assign array_update_74356[6] = add_74316 == 32'h0000_0006 ? add_74354 : array_index_74348[6];
  assign array_update_74356[7] = add_74316 == 32'h0000_0007 ? add_74354 : array_index_74348[7];
  assign array_update_74356[8] = add_74316 == 32'h0000_0008 ? add_74354 : array_index_74348[8];
  assign array_update_74356[9] = add_74316 == 32'h0000_0009 ? add_74354 : array_index_74348[9];
  assign add_74357 = add_74344 + 32'h0000_0001;
  assign array_update_74358[0] = add_73368 == 32'h0000_0000 ? array_update_74356 : array_update_74345[0];
  assign array_update_74358[1] = add_73368 == 32'h0000_0001 ? array_update_74356 : array_update_74345[1];
  assign array_update_74358[2] = add_73368 == 32'h0000_0002 ? array_update_74356 : array_update_74345[2];
  assign array_update_74358[3] = add_73368 == 32'h0000_0003 ? array_update_74356 : array_update_74345[3];
  assign array_update_74358[4] = add_73368 == 32'h0000_0004 ? array_update_74356 : array_update_74345[4];
  assign array_update_74358[5] = add_73368 == 32'h0000_0005 ? array_update_74356 : array_update_74345[5];
  assign array_update_74358[6] = add_73368 == 32'h0000_0006 ? array_update_74356 : array_update_74345[6];
  assign array_update_74358[7] = add_73368 == 32'h0000_0007 ? array_update_74356 : array_update_74345[7];
  assign array_update_74358[8] = add_73368 == 32'h0000_0008 ? array_update_74356 : array_update_74345[8];
  assign array_update_74358[9] = add_73368 == 32'h0000_0009 ? array_update_74356 : array_update_74345[9];
  assign array_index_74360 = array_update_72021[add_74357 > 32'h0000_0009 ? 4'h9 : add_74357[3:0]];
  assign array_index_74361 = array_update_74358[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_74365 = smul32b_32b_x_32b(array_index_73375[add_74357 > 32'h0000_0009 ? 4'h9 : add_74357[3:0]], array_index_74360[add_74316 > 32'h0000_0009 ? 4'h9 : add_74316[3:0]]);
  assign add_74367 = array_index_74361[add_74316 > 32'h0000_0009 ? 4'h9 : add_74316[3:0]] + smul_74365;
  assign array_update_74369[0] = add_74316 == 32'h0000_0000 ? add_74367 : array_index_74361[0];
  assign array_update_74369[1] = add_74316 == 32'h0000_0001 ? add_74367 : array_index_74361[1];
  assign array_update_74369[2] = add_74316 == 32'h0000_0002 ? add_74367 : array_index_74361[2];
  assign array_update_74369[3] = add_74316 == 32'h0000_0003 ? add_74367 : array_index_74361[3];
  assign array_update_74369[4] = add_74316 == 32'h0000_0004 ? add_74367 : array_index_74361[4];
  assign array_update_74369[5] = add_74316 == 32'h0000_0005 ? add_74367 : array_index_74361[5];
  assign array_update_74369[6] = add_74316 == 32'h0000_0006 ? add_74367 : array_index_74361[6];
  assign array_update_74369[7] = add_74316 == 32'h0000_0007 ? add_74367 : array_index_74361[7];
  assign array_update_74369[8] = add_74316 == 32'h0000_0008 ? add_74367 : array_index_74361[8];
  assign array_update_74369[9] = add_74316 == 32'h0000_0009 ? add_74367 : array_index_74361[9];
  assign add_74370 = add_74357 + 32'h0000_0001;
  assign array_update_74371[0] = add_73368 == 32'h0000_0000 ? array_update_74369 : array_update_74358[0];
  assign array_update_74371[1] = add_73368 == 32'h0000_0001 ? array_update_74369 : array_update_74358[1];
  assign array_update_74371[2] = add_73368 == 32'h0000_0002 ? array_update_74369 : array_update_74358[2];
  assign array_update_74371[3] = add_73368 == 32'h0000_0003 ? array_update_74369 : array_update_74358[3];
  assign array_update_74371[4] = add_73368 == 32'h0000_0004 ? array_update_74369 : array_update_74358[4];
  assign array_update_74371[5] = add_73368 == 32'h0000_0005 ? array_update_74369 : array_update_74358[5];
  assign array_update_74371[6] = add_73368 == 32'h0000_0006 ? array_update_74369 : array_update_74358[6];
  assign array_update_74371[7] = add_73368 == 32'h0000_0007 ? array_update_74369 : array_update_74358[7];
  assign array_update_74371[8] = add_73368 == 32'h0000_0008 ? array_update_74369 : array_update_74358[8];
  assign array_update_74371[9] = add_73368 == 32'h0000_0009 ? array_update_74369 : array_update_74358[9];
  assign array_index_74373 = array_update_72021[add_74370 > 32'h0000_0009 ? 4'h9 : add_74370[3:0]];
  assign array_index_74374 = array_update_74371[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_74378 = smul32b_32b_x_32b(array_index_73375[add_74370 > 32'h0000_0009 ? 4'h9 : add_74370[3:0]], array_index_74373[add_74316 > 32'h0000_0009 ? 4'h9 : add_74316[3:0]]);
  assign add_74380 = array_index_74374[add_74316 > 32'h0000_0009 ? 4'h9 : add_74316[3:0]] + smul_74378;
  assign array_update_74382[0] = add_74316 == 32'h0000_0000 ? add_74380 : array_index_74374[0];
  assign array_update_74382[1] = add_74316 == 32'h0000_0001 ? add_74380 : array_index_74374[1];
  assign array_update_74382[2] = add_74316 == 32'h0000_0002 ? add_74380 : array_index_74374[2];
  assign array_update_74382[3] = add_74316 == 32'h0000_0003 ? add_74380 : array_index_74374[3];
  assign array_update_74382[4] = add_74316 == 32'h0000_0004 ? add_74380 : array_index_74374[4];
  assign array_update_74382[5] = add_74316 == 32'h0000_0005 ? add_74380 : array_index_74374[5];
  assign array_update_74382[6] = add_74316 == 32'h0000_0006 ? add_74380 : array_index_74374[6];
  assign array_update_74382[7] = add_74316 == 32'h0000_0007 ? add_74380 : array_index_74374[7];
  assign array_update_74382[8] = add_74316 == 32'h0000_0008 ? add_74380 : array_index_74374[8];
  assign array_update_74382[9] = add_74316 == 32'h0000_0009 ? add_74380 : array_index_74374[9];
  assign add_74383 = add_74370 + 32'h0000_0001;
  assign array_update_74384[0] = add_73368 == 32'h0000_0000 ? array_update_74382 : array_update_74371[0];
  assign array_update_74384[1] = add_73368 == 32'h0000_0001 ? array_update_74382 : array_update_74371[1];
  assign array_update_74384[2] = add_73368 == 32'h0000_0002 ? array_update_74382 : array_update_74371[2];
  assign array_update_74384[3] = add_73368 == 32'h0000_0003 ? array_update_74382 : array_update_74371[3];
  assign array_update_74384[4] = add_73368 == 32'h0000_0004 ? array_update_74382 : array_update_74371[4];
  assign array_update_74384[5] = add_73368 == 32'h0000_0005 ? array_update_74382 : array_update_74371[5];
  assign array_update_74384[6] = add_73368 == 32'h0000_0006 ? array_update_74382 : array_update_74371[6];
  assign array_update_74384[7] = add_73368 == 32'h0000_0007 ? array_update_74382 : array_update_74371[7];
  assign array_update_74384[8] = add_73368 == 32'h0000_0008 ? array_update_74382 : array_update_74371[8];
  assign array_update_74384[9] = add_73368 == 32'h0000_0009 ? array_update_74382 : array_update_74371[9];
  assign array_index_74386 = array_update_72021[add_74383 > 32'h0000_0009 ? 4'h9 : add_74383[3:0]];
  assign array_index_74387 = array_update_74384[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_74391 = smul32b_32b_x_32b(array_index_73375[add_74383 > 32'h0000_0009 ? 4'h9 : add_74383[3:0]], array_index_74386[add_74316 > 32'h0000_0009 ? 4'h9 : add_74316[3:0]]);
  assign add_74393 = array_index_74387[add_74316 > 32'h0000_0009 ? 4'h9 : add_74316[3:0]] + smul_74391;
  assign array_update_74395[0] = add_74316 == 32'h0000_0000 ? add_74393 : array_index_74387[0];
  assign array_update_74395[1] = add_74316 == 32'h0000_0001 ? add_74393 : array_index_74387[1];
  assign array_update_74395[2] = add_74316 == 32'h0000_0002 ? add_74393 : array_index_74387[2];
  assign array_update_74395[3] = add_74316 == 32'h0000_0003 ? add_74393 : array_index_74387[3];
  assign array_update_74395[4] = add_74316 == 32'h0000_0004 ? add_74393 : array_index_74387[4];
  assign array_update_74395[5] = add_74316 == 32'h0000_0005 ? add_74393 : array_index_74387[5];
  assign array_update_74395[6] = add_74316 == 32'h0000_0006 ? add_74393 : array_index_74387[6];
  assign array_update_74395[7] = add_74316 == 32'h0000_0007 ? add_74393 : array_index_74387[7];
  assign array_update_74395[8] = add_74316 == 32'h0000_0008 ? add_74393 : array_index_74387[8];
  assign array_update_74395[9] = add_74316 == 32'h0000_0009 ? add_74393 : array_index_74387[9];
  assign add_74396 = add_74383 + 32'h0000_0001;
  assign array_update_74397[0] = add_73368 == 32'h0000_0000 ? array_update_74395 : array_update_74384[0];
  assign array_update_74397[1] = add_73368 == 32'h0000_0001 ? array_update_74395 : array_update_74384[1];
  assign array_update_74397[2] = add_73368 == 32'h0000_0002 ? array_update_74395 : array_update_74384[2];
  assign array_update_74397[3] = add_73368 == 32'h0000_0003 ? array_update_74395 : array_update_74384[3];
  assign array_update_74397[4] = add_73368 == 32'h0000_0004 ? array_update_74395 : array_update_74384[4];
  assign array_update_74397[5] = add_73368 == 32'h0000_0005 ? array_update_74395 : array_update_74384[5];
  assign array_update_74397[6] = add_73368 == 32'h0000_0006 ? array_update_74395 : array_update_74384[6];
  assign array_update_74397[7] = add_73368 == 32'h0000_0007 ? array_update_74395 : array_update_74384[7];
  assign array_update_74397[8] = add_73368 == 32'h0000_0008 ? array_update_74395 : array_update_74384[8];
  assign array_update_74397[9] = add_73368 == 32'h0000_0009 ? array_update_74395 : array_update_74384[9];
  assign array_index_74399 = array_update_72021[add_74396 > 32'h0000_0009 ? 4'h9 : add_74396[3:0]];
  assign array_index_74400 = array_update_74397[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_74404 = smul32b_32b_x_32b(array_index_73375[add_74396 > 32'h0000_0009 ? 4'h9 : add_74396[3:0]], array_index_74399[add_74316 > 32'h0000_0009 ? 4'h9 : add_74316[3:0]]);
  assign add_74406 = array_index_74400[add_74316 > 32'h0000_0009 ? 4'h9 : add_74316[3:0]] + smul_74404;
  assign array_update_74408[0] = add_74316 == 32'h0000_0000 ? add_74406 : array_index_74400[0];
  assign array_update_74408[1] = add_74316 == 32'h0000_0001 ? add_74406 : array_index_74400[1];
  assign array_update_74408[2] = add_74316 == 32'h0000_0002 ? add_74406 : array_index_74400[2];
  assign array_update_74408[3] = add_74316 == 32'h0000_0003 ? add_74406 : array_index_74400[3];
  assign array_update_74408[4] = add_74316 == 32'h0000_0004 ? add_74406 : array_index_74400[4];
  assign array_update_74408[5] = add_74316 == 32'h0000_0005 ? add_74406 : array_index_74400[5];
  assign array_update_74408[6] = add_74316 == 32'h0000_0006 ? add_74406 : array_index_74400[6];
  assign array_update_74408[7] = add_74316 == 32'h0000_0007 ? add_74406 : array_index_74400[7];
  assign array_update_74408[8] = add_74316 == 32'h0000_0008 ? add_74406 : array_index_74400[8];
  assign array_update_74408[9] = add_74316 == 32'h0000_0009 ? add_74406 : array_index_74400[9];
  assign add_74409 = add_74396 + 32'h0000_0001;
  assign array_update_74410[0] = add_73368 == 32'h0000_0000 ? array_update_74408 : array_update_74397[0];
  assign array_update_74410[1] = add_73368 == 32'h0000_0001 ? array_update_74408 : array_update_74397[1];
  assign array_update_74410[2] = add_73368 == 32'h0000_0002 ? array_update_74408 : array_update_74397[2];
  assign array_update_74410[3] = add_73368 == 32'h0000_0003 ? array_update_74408 : array_update_74397[3];
  assign array_update_74410[4] = add_73368 == 32'h0000_0004 ? array_update_74408 : array_update_74397[4];
  assign array_update_74410[5] = add_73368 == 32'h0000_0005 ? array_update_74408 : array_update_74397[5];
  assign array_update_74410[6] = add_73368 == 32'h0000_0006 ? array_update_74408 : array_update_74397[6];
  assign array_update_74410[7] = add_73368 == 32'h0000_0007 ? array_update_74408 : array_update_74397[7];
  assign array_update_74410[8] = add_73368 == 32'h0000_0008 ? array_update_74408 : array_update_74397[8];
  assign array_update_74410[9] = add_73368 == 32'h0000_0009 ? array_update_74408 : array_update_74397[9];
  assign array_index_74412 = array_update_72021[add_74409 > 32'h0000_0009 ? 4'h9 : add_74409[3:0]];
  assign array_index_74413 = array_update_74410[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_74417 = smul32b_32b_x_32b(array_index_73375[add_74409 > 32'h0000_0009 ? 4'h9 : add_74409[3:0]], array_index_74412[add_74316 > 32'h0000_0009 ? 4'h9 : add_74316[3:0]]);
  assign add_74419 = array_index_74413[add_74316 > 32'h0000_0009 ? 4'h9 : add_74316[3:0]] + smul_74417;
  assign array_update_74421[0] = add_74316 == 32'h0000_0000 ? add_74419 : array_index_74413[0];
  assign array_update_74421[1] = add_74316 == 32'h0000_0001 ? add_74419 : array_index_74413[1];
  assign array_update_74421[2] = add_74316 == 32'h0000_0002 ? add_74419 : array_index_74413[2];
  assign array_update_74421[3] = add_74316 == 32'h0000_0003 ? add_74419 : array_index_74413[3];
  assign array_update_74421[4] = add_74316 == 32'h0000_0004 ? add_74419 : array_index_74413[4];
  assign array_update_74421[5] = add_74316 == 32'h0000_0005 ? add_74419 : array_index_74413[5];
  assign array_update_74421[6] = add_74316 == 32'h0000_0006 ? add_74419 : array_index_74413[6];
  assign array_update_74421[7] = add_74316 == 32'h0000_0007 ? add_74419 : array_index_74413[7];
  assign array_update_74421[8] = add_74316 == 32'h0000_0008 ? add_74419 : array_index_74413[8];
  assign array_update_74421[9] = add_74316 == 32'h0000_0009 ? add_74419 : array_index_74413[9];
  assign add_74422 = add_74409 + 32'h0000_0001;
  assign array_update_74423[0] = add_73368 == 32'h0000_0000 ? array_update_74421 : array_update_74410[0];
  assign array_update_74423[1] = add_73368 == 32'h0000_0001 ? array_update_74421 : array_update_74410[1];
  assign array_update_74423[2] = add_73368 == 32'h0000_0002 ? array_update_74421 : array_update_74410[2];
  assign array_update_74423[3] = add_73368 == 32'h0000_0003 ? array_update_74421 : array_update_74410[3];
  assign array_update_74423[4] = add_73368 == 32'h0000_0004 ? array_update_74421 : array_update_74410[4];
  assign array_update_74423[5] = add_73368 == 32'h0000_0005 ? array_update_74421 : array_update_74410[5];
  assign array_update_74423[6] = add_73368 == 32'h0000_0006 ? array_update_74421 : array_update_74410[6];
  assign array_update_74423[7] = add_73368 == 32'h0000_0007 ? array_update_74421 : array_update_74410[7];
  assign array_update_74423[8] = add_73368 == 32'h0000_0008 ? array_update_74421 : array_update_74410[8];
  assign array_update_74423[9] = add_73368 == 32'h0000_0009 ? array_update_74421 : array_update_74410[9];
  assign array_index_74425 = array_update_72021[add_74422 > 32'h0000_0009 ? 4'h9 : add_74422[3:0]];
  assign array_index_74426 = array_update_74423[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_74430 = smul32b_32b_x_32b(array_index_73375[add_74422 > 32'h0000_0009 ? 4'h9 : add_74422[3:0]], array_index_74425[add_74316 > 32'h0000_0009 ? 4'h9 : add_74316[3:0]]);
  assign add_74432 = array_index_74426[add_74316 > 32'h0000_0009 ? 4'h9 : add_74316[3:0]] + smul_74430;
  assign array_update_74434[0] = add_74316 == 32'h0000_0000 ? add_74432 : array_index_74426[0];
  assign array_update_74434[1] = add_74316 == 32'h0000_0001 ? add_74432 : array_index_74426[1];
  assign array_update_74434[2] = add_74316 == 32'h0000_0002 ? add_74432 : array_index_74426[2];
  assign array_update_74434[3] = add_74316 == 32'h0000_0003 ? add_74432 : array_index_74426[3];
  assign array_update_74434[4] = add_74316 == 32'h0000_0004 ? add_74432 : array_index_74426[4];
  assign array_update_74434[5] = add_74316 == 32'h0000_0005 ? add_74432 : array_index_74426[5];
  assign array_update_74434[6] = add_74316 == 32'h0000_0006 ? add_74432 : array_index_74426[6];
  assign array_update_74434[7] = add_74316 == 32'h0000_0007 ? add_74432 : array_index_74426[7];
  assign array_update_74434[8] = add_74316 == 32'h0000_0008 ? add_74432 : array_index_74426[8];
  assign array_update_74434[9] = add_74316 == 32'h0000_0009 ? add_74432 : array_index_74426[9];
  assign add_74435 = add_74422 + 32'h0000_0001;
  assign array_update_74436[0] = add_73368 == 32'h0000_0000 ? array_update_74434 : array_update_74423[0];
  assign array_update_74436[1] = add_73368 == 32'h0000_0001 ? array_update_74434 : array_update_74423[1];
  assign array_update_74436[2] = add_73368 == 32'h0000_0002 ? array_update_74434 : array_update_74423[2];
  assign array_update_74436[3] = add_73368 == 32'h0000_0003 ? array_update_74434 : array_update_74423[3];
  assign array_update_74436[4] = add_73368 == 32'h0000_0004 ? array_update_74434 : array_update_74423[4];
  assign array_update_74436[5] = add_73368 == 32'h0000_0005 ? array_update_74434 : array_update_74423[5];
  assign array_update_74436[6] = add_73368 == 32'h0000_0006 ? array_update_74434 : array_update_74423[6];
  assign array_update_74436[7] = add_73368 == 32'h0000_0007 ? array_update_74434 : array_update_74423[7];
  assign array_update_74436[8] = add_73368 == 32'h0000_0008 ? array_update_74434 : array_update_74423[8];
  assign array_update_74436[9] = add_73368 == 32'h0000_0009 ? array_update_74434 : array_update_74423[9];
  assign array_index_74438 = array_update_72021[add_74435 > 32'h0000_0009 ? 4'h9 : add_74435[3:0]];
  assign array_index_74439 = array_update_74436[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_74443 = smul32b_32b_x_32b(array_index_73375[add_74435 > 32'h0000_0009 ? 4'h9 : add_74435[3:0]], array_index_74438[add_74316 > 32'h0000_0009 ? 4'h9 : add_74316[3:0]]);
  assign add_74445 = array_index_74439[add_74316 > 32'h0000_0009 ? 4'h9 : add_74316[3:0]] + smul_74443;
  assign array_update_74446[0] = add_74316 == 32'h0000_0000 ? add_74445 : array_index_74439[0];
  assign array_update_74446[1] = add_74316 == 32'h0000_0001 ? add_74445 : array_index_74439[1];
  assign array_update_74446[2] = add_74316 == 32'h0000_0002 ? add_74445 : array_index_74439[2];
  assign array_update_74446[3] = add_74316 == 32'h0000_0003 ? add_74445 : array_index_74439[3];
  assign array_update_74446[4] = add_74316 == 32'h0000_0004 ? add_74445 : array_index_74439[4];
  assign array_update_74446[5] = add_74316 == 32'h0000_0005 ? add_74445 : array_index_74439[5];
  assign array_update_74446[6] = add_74316 == 32'h0000_0006 ? add_74445 : array_index_74439[6];
  assign array_update_74446[7] = add_74316 == 32'h0000_0007 ? add_74445 : array_index_74439[7];
  assign array_update_74446[8] = add_74316 == 32'h0000_0008 ? add_74445 : array_index_74439[8];
  assign array_update_74446[9] = add_74316 == 32'h0000_0009 ? add_74445 : array_index_74439[9];
  assign array_update_74447[0] = add_73368 == 32'h0000_0000 ? array_update_74446 : array_update_74436[0];
  assign array_update_74447[1] = add_73368 == 32'h0000_0001 ? array_update_74446 : array_update_74436[1];
  assign array_update_74447[2] = add_73368 == 32'h0000_0002 ? array_update_74446 : array_update_74436[2];
  assign array_update_74447[3] = add_73368 == 32'h0000_0003 ? array_update_74446 : array_update_74436[3];
  assign array_update_74447[4] = add_73368 == 32'h0000_0004 ? array_update_74446 : array_update_74436[4];
  assign array_update_74447[5] = add_73368 == 32'h0000_0005 ? array_update_74446 : array_update_74436[5];
  assign array_update_74447[6] = add_73368 == 32'h0000_0006 ? array_update_74446 : array_update_74436[6];
  assign array_update_74447[7] = add_73368 == 32'h0000_0007 ? array_update_74446 : array_update_74436[7];
  assign array_update_74447[8] = add_73368 == 32'h0000_0008 ? array_update_74446 : array_update_74436[8];
  assign array_update_74447[9] = add_73368 == 32'h0000_0009 ? array_update_74446 : array_update_74436[9];
  assign array_index_74449 = array_update_74447[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign add_74451 = add_74316 + 32'h0000_0001;
  assign array_update_74452[0] = add_74451 == 32'h0000_0000 ? 32'h0000_0000 : array_index_74449[0];
  assign array_update_74452[1] = add_74451 == 32'h0000_0001 ? 32'h0000_0000 : array_index_74449[1];
  assign array_update_74452[2] = add_74451 == 32'h0000_0002 ? 32'h0000_0000 : array_index_74449[2];
  assign array_update_74452[3] = add_74451 == 32'h0000_0003 ? 32'h0000_0000 : array_index_74449[3];
  assign array_update_74452[4] = add_74451 == 32'h0000_0004 ? 32'h0000_0000 : array_index_74449[4];
  assign array_update_74452[5] = add_74451 == 32'h0000_0005 ? 32'h0000_0000 : array_index_74449[5];
  assign array_update_74452[6] = add_74451 == 32'h0000_0006 ? 32'h0000_0000 : array_index_74449[6];
  assign array_update_74452[7] = add_74451 == 32'h0000_0007 ? 32'h0000_0000 : array_index_74449[7];
  assign array_update_74452[8] = add_74451 == 32'h0000_0008 ? 32'h0000_0000 : array_index_74449[8];
  assign array_update_74452[9] = add_74451 == 32'h0000_0009 ? 32'h0000_0000 : array_index_74449[9];
  assign literal_74453 = 32'h0000_0000;
  assign array_update_74454[0] = add_73368 == 32'h0000_0000 ? array_update_74452 : array_update_74447[0];
  assign array_update_74454[1] = add_73368 == 32'h0000_0001 ? array_update_74452 : array_update_74447[1];
  assign array_update_74454[2] = add_73368 == 32'h0000_0002 ? array_update_74452 : array_update_74447[2];
  assign array_update_74454[3] = add_73368 == 32'h0000_0003 ? array_update_74452 : array_update_74447[3];
  assign array_update_74454[4] = add_73368 == 32'h0000_0004 ? array_update_74452 : array_update_74447[4];
  assign array_update_74454[5] = add_73368 == 32'h0000_0005 ? array_update_74452 : array_update_74447[5];
  assign array_update_74454[6] = add_73368 == 32'h0000_0006 ? array_update_74452 : array_update_74447[6];
  assign array_update_74454[7] = add_73368 == 32'h0000_0007 ? array_update_74452 : array_update_74447[7];
  assign array_update_74454[8] = add_73368 == 32'h0000_0008 ? array_update_74452 : array_update_74447[8];
  assign array_update_74454[9] = add_73368 == 32'h0000_0009 ? array_update_74452 : array_update_74447[9];
  assign array_index_74456 = array_update_72021[literal_74453 > 32'h0000_0009 ? 4'h9 : literal_74453[3:0]];
  assign array_index_74457 = array_update_74454[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_74461 = smul32b_32b_x_32b(array_index_73375[literal_74453 > 32'h0000_0009 ? 4'h9 : literal_74453[3:0]], array_index_74456[add_74451 > 32'h0000_0009 ? 4'h9 : add_74451[3:0]]);
  assign add_74463 = array_index_74457[add_74451 > 32'h0000_0009 ? 4'h9 : add_74451[3:0]] + smul_74461;
  assign array_update_74465[0] = add_74451 == 32'h0000_0000 ? add_74463 : array_index_74457[0];
  assign array_update_74465[1] = add_74451 == 32'h0000_0001 ? add_74463 : array_index_74457[1];
  assign array_update_74465[2] = add_74451 == 32'h0000_0002 ? add_74463 : array_index_74457[2];
  assign array_update_74465[3] = add_74451 == 32'h0000_0003 ? add_74463 : array_index_74457[3];
  assign array_update_74465[4] = add_74451 == 32'h0000_0004 ? add_74463 : array_index_74457[4];
  assign array_update_74465[5] = add_74451 == 32'h0000_0005 ? add_74463 : array_index_74457[5];
  assign array_update_74465[6] = add_74451 == 32'h0000_0006 ? add_74463 : array_index_74457[6];
  assign array_update_74465[7] = add_74451 == 32'h0000_0007 ? add_74463 : array_index_74457[7];
  assign array_update_74465[8] = add_74451 == 32'h0000_0008 ? add_74463 : array_index_74457[8];
  assign array_update_74465[9] = add_74451 == 32'h0000_0009 ? add_74463 : array_index_74457[9];
  assign add_74466 = literal_74453 + 32'h0000_0001;
  assign array_update_74467[0] = add_73368 == 32'h0000_0000 ? array_update_74465 : array_update_74454[0];
  assign array_update_74467[1] = add_73368 == 32'h0000_0001 ? array_update_74465 : array_update_74454[1];
  assign array_update_74467[2] = add_73368 == 32'h0000_0002 ? array_update_74465 : array_update_74454[2];
  assign array_update_74467[3] = add_73368 == 32'h0000_0003 ? array_update_74465 : array_update_74454[3];
  assign array_update_74467[4] = add_73368 == 32'h0000_0004 ? array_update_74465 : array_update_74454[4];
  assign array_update_74467[5] = add_73368 == 32'h0000_0005 ? array_update_74465 : array_update_74454[5];
  assign array_update_74467[6] = add_73368 == 32'h0000_0006 ? array_update_74465 : array_update_74454[6];
  assign array_update_74467[7] = add_73368 == 32'h0000_0007 ? array_update_74465 : array_update_74454[7];
  assign array_update_74467[8] = add_73368 == 32'h0000_0008 ? array_update_74465 : array_update_74454[8];
  assign array_update_74467[9] = add_73368 == 32'h0000_0009 ? array_update_74465 : array_update_74454[9];
  assign array_index_74469 = array_update_72021[add_74466 > 32'h0000_0009 ? 4'h9 : add_74466[3:0]];
  assign array_index_74470 = array_update_74467[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_74474 = smul32b_32b_x_32b(array_index_73375[add_74466 > 32'h0000_0009 ? 4'h9 : add_74466[3:0]], array_index_74469[add_74451 > 32'h0000_0009 ? 4'h9 : add_74451[3:0]]);
  assign add_74476 = array_index_74470[add_74451 > 32'h0000_0009 ? 4'h9 : add_74451[3:0]] + smul_74474;
  assign array_update_74478[0] = add_74451 == 32'h0000_0000 ? add_74476 : array_index_74470[0];
  assign array_update_74478[1] = add_74451 == 32'h0000_0001 ? add_74476 : array_index_74470[1];
  assign array_update_74478[2] = add_74451 == 32'h0000_0002 ? add_74476 : array_index_74470[2];
  assign array_update_74478[3] = add_74451 == 32'h0000_0003 ? add_74476 : array_index_74470[3];
  assign array_update_74478[4] = add_74451 == 32'h0000_0004 ? add_74476 : array_index_74470[4];
  assign array_update_74478[5] = add_74451 == 32'h0000_0005 ? add_74476 : array_index_74470[5];
  assign array_update_74478[6] = add_74451 == 32'h0000_0006 ? add_74476 : array_index_74470[6];
  assign array_update_74478[7] = add_74451 == 32'h0000_0007 ? add_74476 : array_index_74470[7];
  assign array_update_74478[8] = add_74451 == 32'h0000_0008 ? add_74476 : array_index_74470[8];
  assign array_update_74478[9] = add_74451 == 32'h0000_0009 ? add_74476 : array_index_74470[9];
  assign add_74479 = add_74466 + 32'h0000_0001;
  assign array_update_74480[0] = add_73368 == 32'h0000_0000 ? array_update_74478 : array_update_74467[0];
  assign array_update_74480[1] = add_73368 == 32'h0000_0001 ? array_update_74478 : array_update_74467[1];
  assign array_update_74480[2] = add_73368 == 32'h0000_0002 ? array_update_74478 : array_update_74467[2];
  assign array_update_74480[3] = add_73368 == 32'h0000_0003 ? array_update_74478 : array_update_74467[3];
  assign array_update_74480[4] = add_73368 == 32'h0000_0004 ? array_update_74478 : array_update_74467[4];
  assign array_update_74480[5] = add_73368 == 32'h0000_0005 ? array_update_74478 : array_update_74467[5];
  assign array_update_74480[6] = add_73368 == 32'h0000_0006 ? array_update_74478 : array_update_74467[6];
  assign array_update_74480[7] = add_73368 == 32'h0000_0007 ? array_update_74478 : array_update_74467[7];
  assign array_update_74480[8] = add_73368 == 32'h0000_0008 ? array_update_74478 : array_update_74467[8];
  assign array_update_74480[9] = add_73368 == 32'h0000_0009 ? array_update_74478 : array_update_74467[9];
  assign array_index_74482 = array_update_72021[add_74479 > 32'h0000_0009 ? 4'h9 : add_74479[3:0]];
  assign array_index_74483 = array_update_74480[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_74487 = smul32b_32b_x_32b(array_index_73375[add_74479 > 32'h0000_0009 ? 4'h9 : add_74479[3:0]], array_index_74482[add_74451 > 32'h0000_0009 ? 4'h9 : add_74451[3:0]]);
  assign add_74489 = array_index_74483[add_74451 > 32'h0000_0009 ? 4'h9 : add_74451[3:0]] + smul_74487;
  assign array_update_74491[0] = add_74451 == 32'h0000_0000 ? add_74489 : array_index_74483[0];
  assign array_update_74491[1] = add_74451 == 32'h0000_0001 ? add_74489 : array_index_74483[1];
  assign array_update_74491[2] = add_74451 == 32'h0000_0002 ? add_74489 : array_index_74483[2];
  assign array_update_74491[3] = add_74451 == 32'h0000_0003 ? add_74489 : array_index_74483[3];
  assign array_update_74491[4] = add_74451 == 32'h0000_0004 ? add_74489 : array_index_74483[4];
  assign array_update_74491[5] = add_74451 == 32'h0000_0005 ? add_74489 : array_index_74483[5];
  assign array_update_74491[6] = add_74451 == 32'h0000_0006 ? add_74489 : array_index_74483[6];
  assign array_update_74491[7] = add_74451 == 32'h0000_0007 ? add_74489 : array_index_74483[7];
  assign array_update_74491[8] = add_74451 == 32'h0000_0008 ? add_74489 : array_index_74483[8];
  assign array_update_74491[9] = add_74451 == 32'h0000_0009 ? add_74489 : array_index_74483[9];
  assign add_74492 = add_74479 + 32'h0000_0001;
  assign array_update_74493[0] = add_73368 == 32'h0000_0000 ? array_update_74491 : array_update_74480[0];
  assign array_update_74493[1] = add_73368 == 32'h0000_0001 ? array_update_74491 : array_update_74480[1];
  assign array_update_74493[2] = add_73368 == 32'h0000_0002 ? array_update_74491 : array_update_74480[2];
  assign array_update_74493[3] = add_73368 == 32'h0000_0003 ? array_update_74491 : array_update_74480[3];
  assign array_update_74493[4] = add_73368 == 32'h0000_0004 ? array_update_74491 : array_update_74480[4];
  assign array_update_74493[5] = add_73368 == 32'h0000_0005 ? array_update_74491 : array_update_74480[5];
  assign array_update_74493[6] = add_73368 == 32'h0000_0006 ? array_update_74491 : array_update_74480[6];
  assign array_update_74493[7] = add_73368 == 32'h0000_0007 ? array_update_74491 : array_update_74480[7];
  assign array_update_74493[8] = add_73368 == 32'h0000_0008 ? array_update_74491 : array_update_74480[8];
  assign array_update_74493[9] = add_73368 == 32'h0000_0009 ? array_update_74491 : array_update_74480[9];
  assign array_index_74495 = array_update_72021[add_74492 > 32'h0000_0009 ? 4'h9 : add_74492[3:0]];
  assign array_index_74496 = array_update_74493[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_74500 = smul32b_32b_x_32b(array_index_73375[add_74492 > 32'h0000_0009 ? 4'h9 : add_74492[3:0]], array_index_74495[add_74451 > 32'h0000_0009 ? 4'h9 : add_74451[3:0]]);
  assign add_74502 = array_index_74496[add_74451 > 32'h0000_0009 ? 4'h9 : add_74451[3:0]] + smul_74500;
  assign array_update_74504[0] = add_74451 == 32'h0000_0000 ? add_74502 : array_index_74496[0];
  assign array_update_74504[1] = add_74451 == 32'h0000_0001 ? add_74502 : array_index_74496[1];
  assign array_update_74504[2] = add_74451 == 32'h0000_0002 ? add_74502 : array_index_74496[2];
  assign array_update_74504[3] = add_74451 == 32'h0000_0003 ? add_74502 : array_index_74496[3];
  assign array_update_74504[4] = add_74451 == 32'h0000_0004 ? add_74502 : array_index_74496[4];
  assign array_update_74504[5] = add_74451 == 32'h0000_0005 ? add_74502 : array_index_74496[5];
  assign array_update_74504[6] = add_74451 == 32'h0000_0006 ? add_74502 : array_index_74496[6];
  assign array_update_74504[7] = add_74451 == 32'h0000_0007 ? add_74502 : array_index_74496[7];
  assign array_update_74504[8] = add_74451 == 32'h0000_0008 ? add_74502 : array_index_74496[8];
  assign array_update_74504[9] = add_74451 == 32'h0000_0009 ? add_74502 : array_index_74496[9];
  assign add_74505 = add_74492 + 32'h0000_0001;
  assign array_update_74506[0] = add_73368 == 32'h0000_0000 ? array_update_74504 : array_update_74493[0];
  assign array_update_74506[1] = add_73368 == 32'h0000_0001 ? array_update_74504 : array_update_74493[1];
  assign array_update_74506[2] = add_73368 == 32'h0000_0002 ? array_update_74504 : array_update_74493[2];
  assign array_update_74506[3] = add_73368 == 32'h0000_0003 ? array_update_74504 : array_update_74493[3];
  assign array_update_74506[4] = add_73368 == 32'h0000_0004 ? array_update_74504 : array_update_74493[4];
  assign array_update_74506[5] = add_73368 == 32'h0000_0005 ? array_update_74504 : array_update_74493[5];
  assign array_update_74506[6] = add_73368 == 32'h0000_0006 ? array_update_74504 : array_update_74493[6];
  assign array_update_74506[7] = add_73368 == 32'h0000_0007 ? array_update_74504 : array_update_74493[7];
  assign array_update_74506[8] = add_73368 == 32'h0000_0008 ? array_update_74504 : array_update_74493[8];
  assign array_update_74506[9] = add_73368 == 32'h0000_0009 ? array_update_74504 : array_update_74493[9];
  assign array_index_74508 = array_update_72021[add_74505 > 32'h0000_0009 ? 4'h9 : add_74505[3:0]];
  assign array_index_74509 = array_update_74506[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_74513 = smul32b_32b_x_32b(array_index_73375[add_74505 > 32'h0000_0009 ? 4'h9 : add_74505[3:0]], array_index_74508[add_74451 > 32'h0000_0009 ? 4'h9 : add_74451[3:0]]);
  assign add_74515 = array_index_74509[add_74451 > 32'h0000_0009 ? 4'h9 : add_74451[3:0]] + smul_74513;
  assign array_update_74517[0] = add_74451 == 32'h0000_0000 ? add_74515 : array_index_74509[0];
  assign array_update_74517[1] = add_74451 == 32'h0000_0001 ? add_74515 : array_index_74509[1];
  assign array_update_74517[2] = add_74451 == 32'h0000_0002 ? add_74515 : array_index_74509[2];
  assign array_update_74517[3] = add_74451 == 32'h0000_0003 ? add_74515 : array_index_74509[3];
  assign array_update_74517[4] = add_74451 == 32'h0000_0004 ? add_74515 : array_index_74509[4];
  assign array_update_74517[5] = add_74451 == 32'h0000_0005 ? add_74515 : array_index_74509[5];
  assign array_update_74517[6] = add_74451 == 32'h0000_0006 ? add_74515 : array_index_74509[6];
  assign array_update_74517[7] = add_74451 == 32'h0000_0007 ? add_74515 : array_index_74509[7];
  assign array_update_74517[8] = add_74451 == 32'h0000_0008 ? add_74515 : array_index_74509[8];
  assign array_update_74517[9] = add_74451 == 32'h0000_0009 ? add_74515 : array_index_74509[9];
  assign add_74518 = add_74505 + 32'h0000_0001;
  assign array_update_74519[0] = add_73368 == 32'h0000_0000 ? array_update_74517 : array_update_74506[0];
  assign array_update_74519[1] = add_73368 == 32'h0000_0001 ? array_update_74517 : array_update_74506[1];
  assign array_update_74519[2] = add_73368 == 32'h0000_0002 ? array_update_74517 : array_update_74506[2];
  assign array_update_74519[3] = add_73368 == 32'h0000_0003 ? array_update_74517 : array_update_74506[3];
  assign array_update_74519[4] = add_73368 == 32'h0000_0004 ? array_update_74517 : array_update_74506[4];
  assign array_update_74519[5] = add_73368 == 32'h0000_0005 ? array_update_74517 : array_update_74506[5];
  assign array_update_74519[6] = add_73368 == 32'h0000_0006 ? array_update_74517 : array_update_74506[6];
  assign array_update_74519[7] = add_73368 == 32'h0000_0007 ? array_update_74517 : array_update_74506[7];
  assign array_update_74519[8] = add_73368 == 32'h0000_0008 ? array_update_74517 : array_update_74506[8];
  assign array_update_74519[9] = add_73368 == 32'h0000_0009 ? array_update_74517 : array_update_74506[9];
  assign array_index_74521 = array_update_72021[add_74518 > 32'h0000_0009 ? 4'h9 : add_74518[3:0]];
  assign array_index_74522 = array_update_74519[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_74526 = smul32b_32b_x_32b(array_index_73375[add_74518 > 32'h0000_0009 ? 4'h9 : add_74518[3:0]], array_index_74521[add_74451 > 32'h0000_0009 ? 4'h9 : add_74451[3:0]]);
  assign add_74528 = array_index_74522[add_74451 > 32'h0000_0009 ? 4'h9 : add_74451[3:0]] + smul_74526;
  assign array_update_74530[0] = add_74451 == 32'h0000_0000 ? add_74528 : array_index_74522[0];
  assign array_update_74530[1] = add_74451 == 32'h0000_0001 ? add_74528 : array_index_74522[1];
  assign array_update_74530[2] = add_74451 == 32'h0000_0002 ? add_74528 : array_index_74522[2];
  assign array_update_74530[3] = add_74451 == 32'h0000_0003 ? add_74528 : array_index_74522[3];
  assign array_update_74530[4] = add_74451 == 32'h0000_0004 ? add_74528 : array_index_74522[4];
  assign array_update_74530[5] = add_74451 == 32'h0000_0005 ? add_74528 : array_index_74522[5];
  assign array_update_74530[6] = add_74451 == 32'h0000_0006 ? add_74528 : array_index_74522[6];
  assign array_update_74530[7] = add_74451 == 32'h0000_0007 ? add_74528 : array_index_74522[7];
  assign array_update_74530[8] = add_74451 == 32'h0000_0008 ? add_74528 : array_index_74522[8];
  assign array_update_74530[9] = add_74451 == 32'h0000_0009 ? add_74528 : array_index_74522[9];
  assign add_74531 = add_74518 + 32'h0000_0001;
  assign array_update_74532[0] = add_73368 == 32'h0000_0000 ? array_update_74530 : array_update_74519[0];
  assign array_update_74532[1] = add_73368 == 32'h0000_0001 ? array_update_74530 : array_update_74519[1];
  assign array_update_74532[2] = add_73368 == 32'h0000_0002 ? array_update_74530 : array_update_74519[2];
  assign array_update_74532[3] = add_73368 == 32'h0000_0003 ? array_update_74530 : array_update_74519[3];
  assign array_update_74532[4] = add_73368 == 32'h0000_0004 ? array_update_74530 : array_update_74519[4];
  assign array_update_74532[5] = add_73368 == 32'h0000_0005 ? array_update_74530 : array_update_74519[5];
  assign array_update_74532[6] = add_73368 == 32'h0000_0006 ? array_update_74530 : array_update_74519[6];
  assign array_update_74532[7] = add_73368 == 32'h0000_0007 ? array_update_74530 : array_update_74519[7];
  assign array_update_74532[8] = add_73368 == 32'h0000_0008 ? array_update_74530 : array_update_74519[8];
  assign array_update_74532[9] = add_73368 == 32'h0000_0009 ? array_update_74530 : array_update_74519[9];
  assign array_index_74534 = array_update_72021[add_74531 > 32'h0000_0009 ? 4'h9 : add_74531[3:0]];
  assign array_index_74535 = array_update_74532[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_74539 = smul32b_32b_x_32b(array_index_73375[add_74531 > 32'h0000_0009 ? 4'h9 : add_74531[3:0]], array_index_74534[add_74451 > 32'h0000_0009 ? 4'h9 : add_74451[3:0]]);
  assign add_74541 = array_index_74535[add_74451 > 32'h0000_0009 ? 4'h9 : add_74451[3:0]] + smul_74539;
  assign array_update_74543[0] = add_74451 == 32'h0000_0000 ? add_74541 : array_index_74535[0];
  assign array_update_74543[1] = add_74451 == 32'h0000_0001 ? add_74541 : array_index_74535[1];
  assign array_update_74543[2] = add_74451 == 32'h0000_0002 ? add_74541 : array_index_74535[2];
  assign array_update_74543[3] = add_74451 == 32'h0000_0003 ? add_74541 : array_index_74535[3];
  assign array_update_74543[4] = add_74451 == 32'h0000_0004 ? add_74541 : array_index_74535[4];
  assign array_update_74543[5] = add_74451 == 32'h0000_0005 ? add_74541 : array_index_74535[5];
  assign array_update_74543[6] = add_74451 == 32'h0000_0006 ? add_74541 : array_index_74535[6];
  assign array_update_74543[7] = add_74451 == 32'h0000_0007 ? add_74541 : array_index_74535[7];
  assign array_update_74543[8] = add_74451 == 32'h0000_0008 ? add_74541 : array_index_74535[8];
  assign array_update_74543[9] = add_74451 == 32'h0000_0009 ? add_74541 : array_index_74535[9];
  assign add_74544 = add_74531 + 32'h0000_0001;
  assign array_update_74545[0] = add_73368 == 32'h0000_0000 ? array_update_74543 : array_update_74532[0];
  assign array_update_74545[1] = add_73368 == 32'h0000_0001 ? array_update_74543 : array_update_74532[1];
  assign array_update_74545[2] = add_73368 == 32'h0000_0002 ? array_update_74543 : array_update_74532[2];
  assign array_update_74545[3] = add_73368 == 32'h0000_0003 ? array_update_74543 : array_update_74532[3];
  assign array_update_74545[4] = add_73368 == 32'h0000_0004 ? array_update_74543 : array_update_74532[4];
  assign array_update_74545[5] = add_73368 == 32'h0000_0005 ? array_update_74543 : array_update_74532[5];
  assign array_update_74545[6] = add_73368 == 32'h0000_0006 ? array_update_74543 : array_update_74532[6];
  assign array_update_74545[7] = add_73368 == 32'h0000_0007 ? array_update_74543 : array_update_74532[7];
  assign array_update_74545[8] = add_73368 == 32'h0000_0008 ? array_update_74543 : array_update_74532[8];
  assign array_update_74545[9] = add_73368 == 32'h0000_0009 ? array_update_74543 : array_update_74532[9];
  assign array_index_74547 = array_update_72021[add_74544 > 32'h0000_0009 ? 4'h9 : add_74544[3:0]];
  assign array_index_74548 = array_update_74545[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_74552 = smul32b_32b_x_32b(array_index_73375[add_74544 > 32'h0000_0009 ? 4'h9 : add_74544[3:0]], array_index_74547[add_74451 > 32'h0000_0009 ? 4'h9 : add_74451[3:0]]);
  assign add_74554 = array_index_74548[add_74451 > 32'h0000_0009 ? 4'h9 : add_74451[3:0]] + smul_74552;
  assign array_update_74556[0] = add_74451 == 32'h0000_0000 ? add_74554 : array_index_74548[0];
  assign array_update_74556[1] = add_74451 == 32'h0000_0001 ? add_74554 : array_index_74548[1];
  assign array_update_74556[2] = add_74451 == 32'h0000_0002 ? add_74554 : array_index_74548[2];
  assign array_update_74556[3] = add_74451 == 32'h0000_0003 ? add_74554 : array_index_74548[3];
  assign array_update_74556[4] = add_74451 == 32'h0000_0004 ? add_74554 : array_index_74548[4];
  assign array_update_74556[5] = add_74451 == 32'h0000_0005 ? add_74554 : array_index_74548[5];
  assign array_update_74556[6] = add_74451 == 32'h0000_0006 ? add_74554 : array_index_74548[6];
  assign array_update_74556[7] = add_74451 == 32'h0000_0007 ? add_74554 : array_index_74548[7];
  assign array_update_74556[8] = add_74451 == 32'h0000_0008 ? add_74554 : array_index_74548[8];
  assign array_update_74556[9] = add_74451 == 32'h0000_0009 ? add_74554 : array_index_74548[9];
  assign add_74557 = add_74544 + 32'h0000_0001;
  assign array_update_74558[0] = add_73368 == 32'h0000_0000 ? array_update_74556 : array_update_74545[0];
  assign array_update_74558[1] = add_73368 == 32'h0000_0001 ? array_update_74556 : array_update_74545[1];
  assign array_update_74558[2] = add_73368 == 32'h0000_0002 ? array_update_74556 : array_update_74545[2];
  assign array_update_74558[3] = add_73368 == 32'h0000_0003 ? array_update_74556 : array_update_74545[3];
  assign array_update_74558[4] = add_73368 == 32'h0000_0004 ? array_update_74556 : array_update_74545[4];
  assign array_update_74558[5] = add_73368 == 32'h0000_0005 ? array_update_74556 : array_update_74545[5];
  assign array_update_74558[6] = add_73368 == 32'h0000_0006 ? array_update_74556 : array_update_74545[6];
  assign array_update_74558[7] = add_73368 == 32'h0000_0007 ? array_update_74556 : array_update_74545[7];
  assign array_update_74558[8] = add_73368 == 32'h0000_0008 ? array_update_74556 : array_update_74545[8];
  assign array_update_74558[9] = add_73368 == 32'h0000_0009 ? array_update_74556 : array_update_74545[9];
  assign array_index_74560 = array_update_72021[add_74557 > 32'h0000_0009 ? 4'h9 : add_74557[3:0]];
  assign array_index_74561 = array_update_74558[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_74565 = smul32b_32b_x_32b(array_index_73375[add_74557 > 32'h0000_0009 ? 4'h9 : add_74557[3:0]], array_index_74560[add_74451 > 32'h0000_0009 ? 4'h9 : add_74451[3:0]]);
  assign add_74567 = array_index_74561[add_74451 > 32'h0000_0009 ? 4'h9 : add_74451[3:0]] + smul_74565;
  assign array_update_74569[0] = add_74451 == 32'h0000_0000 ? add_74567 : array_index_74561[0];
  assign array_update_74569[1] = add_74451 == 32'h0000_0001 ? add_74567 : array_index_74561[1];
  assign array_update_74569[2] = add_74451 == 32'h0000_0002 ? add_74567 : array_index_74561[2];
  assign array_update_74569[3] = add_74451 == 32'h0000_0003 ? add_74567 : array_index_74561[3];
  assign array_update_74569[4] = add_74451 == 32'h0000_0004 ? add_74567 : array_index_74561[4];
  assign array_update_74569[5] = add_74451 == 32'h0000_0005 ? add_74567 : array_index_74561[5];
  assign array_update_74569[6] = add_74451 == 32'h0000_0006 ? add_74567 : array_index_74561[6];
  assign array_update_74569[7] = add_74451 == 32'h0000_0007 ? add_74567 : array_index_74561[7];
  assign array_update_74569[8] = add_74451 == 32'h0000_0008 ? add_74567 : array_index_74561[8];
  assign array_update_74569[9] = add_74451 == 32'h0000_0009 ? add_74567 : array_index_74561[9];
  assign add_74570 = add_74557 + 32'h0000_0001;
  assign array_update_74571[0] = add_73368 == 32'h0000_0000 ? array_update_74569 : array_update_74558[0];
  assign array_update_74571[1] = add_73368 == 32'h0000_0001 ? array_update_74569 : array_update_74558[1];
  assign array_update_74571[2] = add_73368 == 32'h0000_0002 ? array_update_74569 : array_update_74558[2];
  assign array_update_74571[3] = add_73368 == 32'h0000_0003 ? array_update_74569 : array_update_74558[3];
  assign array_update_74571[4] = add_73368 == 32'h0000_0004 ? array_update_74569 : array_update_74558[4];
  assign array_update_74571[5] = add_73368 == 32'h0000_0005 ? array_update_74569 : array_update_74558[5];
  assign array_update_74571[6] = add_73368 == 32'h0000_0006 ? array_update_74569 : array_update_74558[6];
  assign array_update_74571[7] = add_73368 == 32'h0000_0007 ? array_update_74569 : array_update_74558[7];
  assign array_update_74571[8] = add_73368 == 32'h0000_0008 ? array_update_74569 : array_update_74558[8];
  assign array_update_74571[9] = add_73368 == 32'h0000_0009 ? array_update_74569 : array_update_74558[9];
  assign array_index_74573 = array_update_72021[add_74570 > 32'h0000_0009 ? 4'h9 : add_74570[3:0]];
  assign array_index_74574 = array_update_74571[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_74578 = smul32b_32b_x_32b(array_index_73375[add_74570 > 32'h0000_0009 ? 4'h9 : add_74570[3:0]], array_index_74573[add_74451 > 32'h0000_0009 ? 4'h9 : add_74451[3:0]]);
  assign add_74580 = array_index_74574[add_74451 > 32'h0000_0009 ? 4'h9 : add_74451[3:0]] + smul_74578;
  assign array_update_74581[0] = add_74451 == 32'h0000_0000 ? add_74580 : array_index_74574[0];
  assign array_update_74581[1] = add_74451 == 32'h0000_0001 ? add_74580 : array_index_74574[1];
  assign array_update_74581[2] = add_74451 == 32'h0000_0002 ? add_74580 : array_index_74574[2];
  assign array_update_74581[3] = add_74451 == 32'h0000_0003 ? add_74580 : array_index_74574[3];
  assign array_update_74581[4] = add_74451 == 32'h0000_0004 ? add_74580 : array_index_74574[4];
  assign array_update_74581[5] = add_74451 == 32'h0000_0005 ? add_74580 : array_index_74574[5];
  assign array_update_74581[6] = add_74451 == 32'h0000_0006 ? add_74580 : array_index_74574[6];
  assign array_update_74581[7] = add_74451 == 32'h0000_0007 ? add_74580 : array_index_74574[7];
  assign array_update_74581[8] = add_74451 == 32'h0000_0008 ? add_74580 : array_index_74574[8];
  assign array_update_74581[9] = add_74451 == 32'h0000_0009 ? add_74580 : array_index_74574[9];
  assign array_update_74582[0] = add_73368 == 32'h0000_0000 ? array_update_74581 : array_update_74571[0];
  assign array_update_74582[1] = add_73368 == 32'h0000_0001 ? array_update_74581 : array_update_74571[1];
  assign array_update_74582[2] = add_73368 == 32'h0000_0002 ? array_update_74581 : array_update_74571[2];
  assign array_update_74582[3] = add_73368 == 32'h0000_0003 ? array_update_74581 : array_update_74571[3];
  assign array_update_74582[4] = add_73368 == 32'h0000_0004 ? array_update_74581 : array_update_74571[4];
  assign array_update_74582[5] = add_73368 == 32'h0000_0005 ? array_update_74581 : array_update_74571[5];
  assign array_update_74582[6] = add_73368 == 32'h0000_0006 ? array_update_74581 : array_update_74571[6];
  assign array_update_74582[7] = add_73368 == 32'h0000_0007 ? array_update_74581 : array_update_74571[7];
  assign array_update_74582[8] = add_73368 == 32'h0000_0008 ? array_update_74581 : array_update_74571[8];
  assign array_update_74582[9] = add_73368 == 32'h0000_0009 ? array_update_74581 : array_update_74571[9];
  assign array_index_74584 = array_update_74582[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign add_74586 = add_74451 + 32'h0000_0001;
  assign array_update_74587[0] = add_74586 == 32'h0000_0000 ? 32'h0000_0000 : array_index_74584[0];
  assign array_update_74587[1] = add_74586 == 32'h0000_0001 ? 32'h0000_0000 : array_index_74584[1];
  assign array_update_74587[2] = add_74586 == 32'h0000_0002 ? 32'h0000_0000 : array_index_74584[2];
  assign array_update_74587[3] = add_74586 == 32'h0000_0003 ? 32'h0000_0000 : array_index_74584[3];
  assign array_update_74587[4] = add_74586 == 32'h0000_0004 ? 32'h0000_0000 : array_index_74584[4];
  assign array_update_74587[5] = add_74586 == 32'h0000_0005 ? 32'h0000_0000 : array_index_74584[5];
  assign array_update_74587[6] = add_74586 == 32'h0000_0006 ? 32'h0000_0000 : array_index_74584[6];
  assign array_update_74587[7] = add_74586 == 32'h0000_0007 ? 32'h0000_0000 : array_index_74584[7];
  assign array_update_74587[8] = add_74586 == 32'h0000_0008 ? 32'h0000_0000 : array_index_74584[8];
  assign array_update_74587[9] = add_74586 == 32'h0000_0009 ? 32'h0000_0000 : array_index_74584[9];
  assign literal_74588 = 32'h0000_0000;
  assign array_update_74589[0] = add_73368 == 32'h0000_0000 ? array_update_74587 : array_update_74582[0];
  assign array_update_74589[1] = add_73368 == 32'h0000_0001 ? array_update_74587 : array_update_74582[1];
  assign array_update_74589[2] = add_73368 == 32'h0000_0002 ? array_update_74587 : array_update_74582[2];
  assign array_update_74589[3] = add_73368 == 32'h0000_0003 ? array_update_74587 : array_update_74582[3];
  assign array_update_74589[4] = add_73368 == 32'h0000_0004 ? array_update_74587 : array_update_74582[4];
  assign array_update_74589[5] = add_73368 == 32'h0000_0005 ? array_update_74587 : array_update_74582[5];
  assign array_update_74589[6] = add_73368 == 32'h0000_0006 ? array_update_74587 : array_update_74582[6];
  assign array_update_74589[7] = add_73368 == 32'h0000_0007 ? array_update_74587 : array_update_74582[7];
  assign array_update_74589[8] = add_73368 == 32'h0000_0008 ? array_update_74587 : array_update_74582[8];
  assign array_update_74589[9] = add_73368 == 32'h0000_0009 ? array_update_74587 : array_update_74582[9];
  assign array_index_74591 = array_update_72021[literal_74588 > 32'h0000_0009 ? 4'h9 : literal_74588[3:0]];
  assign array_index_74592 = array_update_74589[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_74596 = smul32b_32b_x_32b(array_index_73375[literal_74588 > 32'h0000_0009 ? 4'h9 : literal_74588[3:0]], array_index_74591[add_74586 > 32'h0000_0009 ? 4'h9 : add_74586[3:0]]);
  assign add_74598 = array_index_74592[add_74586 > 32'h0000_0009 ? 4'h9 : add_74586[3:0]] + smul_74596;
  assign array_update_74600[0] = add_74586 == 32'h0000_0000 ? add_74598 : array_index_74592[0];
  assign array_update_74600[1] = add_74586 == 32'h0000_0001 ? add_74598 : array_index_74592[1];
  assign array_update_74600[2] = add_74586 == 32'h0000_0002 ? add_74598 : array_index_74592[2];
  assign array_update_74600[3] = add_74586 == 32'h0000_0003 ? add_74598 : array_index_74592[3];
  assign array_update_74600[4] = add_74586 == 32'h0000_0004 ? add_74598 : array_index_74592[4];
  assign array_update_74600[5] = add_74586 == 32'h0000_0005 ? add_74598 : array_index_74592[5];
  assign array_update_74600[6] = add_74586 == 32'h0000_0006 ? add_74598 : array_index_74592[6];
  assign array_update_74600[7] = add_74586 == 32'h0000_0007 ? add_74598 : array_index_74592[7];
  assign array_update_74600[8] = add_74586 == 32'h0000_0008 ? add_74598 : array_index_74592[8];
  assign array_update_74600[9] = add_74586 == 32'h0000_0009 ? add_74598 : array_index_74592[9];
  assign add_74601 = literal_74588 + 32'h0000_0001;
  assign array_update_74602[0] = add_73368 == 32'h0000_0000 ? array_update_74600 : array_update_74589[0];
  assign array_update_74602[1] = add_73368 == 32'h0000_0001 ? array_update_74600 : array_update_74589[1];
  assign array_update_74602[2] = add_73368 == 32'h0000_0002 ? array_update_74600 : array_update_74589[2];
  assign array_update_74602[3] = add_73368 == 32'h0000_0003 ? array_update_74600 : array_update_74589[3];
  assign array_update_74602[4] = add_73368 == 32'h0000_0004 ? array_update_74600 : array_update_74589[4];
  assign array_update_74602[5] = add_73368 == 32'h0000_0005 ? array_update_74600 : array_update_74589[5];
  assign array_update_74602[6] = add_73368 == 32'h0000_0006 ? array_update_74600 : array_update_74589[6];
  assign array_update_74602[7] = add_73368 == 32'h0000_0007 ? array_update_74600 : array_update_74589[7];
  assign array_update_74602[8] = add_73368 == 32'h0000_0008 ? array_update_74600 : array_update_74589[8];
  assign array_update_74602[9] = add_73368 == 32'h0000_0009 ? array_update_74600 : array_update_74589[9];
  assign array_index_74604 = array_update_72021[add_74601 > 32'h0000_0009 ? 4'h9 : add_74601[3:0]];
  assign array_index_74605 = array_update_74602[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_74609 = smul32b_32b_x_32b(array_index_73375[add_74601 > 32'h0000_0009 ? 4'h9 : add_74601[3:0]], array_index_74604[add_74586 > 32'h0000_0009 ? 4'h9 : add_74586[3:0]]);
  assign add_74611 = array_index_74605[add_74586 > 32'h0000_0009 ? 4'h9 : add_74586[3:0]] + smul_74609;
  assign array_update_74613[0] = add_74586 == 32'h0000_0000 ? add_74611 : array_index_74605[0];
  assign array_update_74613[1] = add_74586 == 32'h0000_0001 ? add_74611 : array_index_74605[1];
  assign array_update_74613[2] = add_74586 == 32'h0000_0002 ? add_74611 : array_index_74605[2];
  assign array_update_74613[3] = add_74586 == 32'h0000_0003 ? add_74611 : array_index_74605[3];
  assign array_update_74613[4] = add_74586 == 32'h0000_0004 ? add_74611 : array_index_74605[4];
  assign array_update_74613[5] = add_74586 == 32'h0000_0005 ? add_74611 : array_index_74605[5];
  assign array_update_74613[6] = add_74586 == 32'h0000_0006 ? add_74611 : array_index_74605[6];
  assign array_update_74613[7] = add_74586 == 32'h0000_0007 ? add_74611 : array_index_74605[7];
  assign array_update_74613[8] = add_74586 == 32'h0000_0008 ? add_74611 : array_index_74605[8];
  assign array_update_74613[9] = add_74586 == 32'h0000_0009 ? add_74611 : array_index_74605[9];
  assign add_74614 = add_74601 + 32'h0000_0001;
  assign array_update_74615[0] = add_73368 == 32'h0000_0000 ? array_update_74613 : array_update_74602[0];
  assign array_update_74615[1] = add_73368 == 32'h0000_0001 ? array_update_74613 : array_update_74602[1];
  assign array_update_74615[2] = add_73368 == 32'h0000_0002 ? array_update_74613 : array_update_74602[2];
  assign array_update_74615[3] = add_73368 == 32'h0000_0003 ? array_update_74613 : array_update_74602[3];
  assign array_update_74615[4] = add_73368 == 32'h0000_0004 ? array_update_74613 : array_update_74602[4];
  assign array_update_74615[5] = add_73368 == 32'h0000_0005 ? array_update_74613 : array_update_74602[5];
  assign array_update_74615[6] = add_73368 == 32'h0000_0006 ? array_update_74613 : array_update_74602[6];
  assign array_update_74615[7] = add_73368 == 32'h0000_0007 ? array_update_74613 : array_update_74602[7];
  assign array_update_74615[8] = add_73368 == 32'h0000_0008 ? array_update_74613 : array_update_74602[8];
  assign array_update_74615[9] = add_73368 == 32'h0000_0009 ? array_update_74613 : array_update_74602[9];
  assign array_index_74617 = array_update_72021[add_74614 > 32'h0000_0009 ? 4'h9 : add_74614[3:0]];
  assign array_index_74618 = array_update_74615[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_74622 = smul32b_32b_x_32b(array_index_73375[add_74614 > 32'h0000_0009 ? 4'h9 : add_74614[3:0]], array_index_74617[add_74586 > 32'h0000_0009 ? 4'h9 : add_74586[3:0]]);
  assign add_74624 = array_index_74618[add_74586 > 32'h0000_0009 ? 4'h9 : add_74586[3:0]] + smul_74622;
  assign array_update_74626[0] = add_74586 == 32'h0000_0000 ? add_74624 : array_index_74618[0];
  assign array_update_74626[1] = add_74586 == 32'h0000_0001 ? add_74624 : array_index_74618[1];
  assign array_update_74626[2] = add_74586 == 32'h0000_0002 ? add_74624 : array_index_74618[2];
  assign array_update_74626[3] = add_74586 == 32'h0000_0003 ? add_74624 : array_index_74618[3];
  assign array_update_74626[4] = add_74586 == 32'h0000_0004 ? add_74624 : array_index_74618[4];
  assign array_update_74626[5] = add_74586 == 32'h0000_0005 ? add_74624 : array_index_74618[5];
  assign array_update_74626[6] = add_74586 == 32'h0000_0006 ? add_74624 : array_index_74618[6];
  assign array_update_74626[7] = add_74586 == 32'h0000_0007 ? add_74624 : array_index_74618[7];
  assign array_update_74626[8] = add_74586 == 32'h0000_0008 ? add_74624 : array_index_74618[8];
  assign array_update_74626[9] = add_74586 == 32'h0000_0009 ? add_74624 : array_index_74618[9];
  assign add_74627 = add_74614 + 32'h0000_0001;
  assign array_update_74628[0] = add_73368 == 32'h0000_0000 ? array_update_74626 : array_update_74615[0];
  assign array_update_74628[1] = add_73368 == 32'h0000_0001 ? array_update_74626 : array_update_74615[1];
  assign array_update_74628[2] = add_73368 == 32'h0000_0002 ? array_update_74626 : array_update_74615[2];
  assign array_update_74628[3] = add_73368 == 32'h0000_0003 ? array_update_74626 : array_update_74615[3];
  assign array_update_74628[4] = add_73368 == 32'h0000_0004 ? array_update_74626 : array_update_74615[4];
  assign array_update_74628[5] = add_73368 == 32'h0000_0005 ? array_update_74626 : array_update_74615[5];
  assign array_update_74628[6] = add_73368 == 32'h0000_0006 ? array_update_74626 : array_update_74615[6];
  assign array_update_74628[7] = add_73368 == 32'h0000_0007 ? array_update_74626 : array_update_74615[7];
  assign array_update_74628[8] = add_73368 == 32'h0000_0008 ? array_update_74626 : array_update_74615[8];
  assign array_update_74628[9] = add_73368 == 32'h0000_0009 ? array_update_74626 : array_update_74615[9];
  assign array_index_74630 = array_update_72021[add_74627 > 32'h0000_0009 ? 4'h9 : add_74627[3:0]];
  assign array_index_74631 = array_update_74628[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_74635 = smul32b_32b_x_32b(array_index_73375[add_74627 > 32'h0000_0009 ? 4'h9 : add_74627[3:0]], array_index_74630[add_74586 > 32'h0000_0009 ? 4'h9 : add_74586[3:0]]);
  assign add_74637 = array_index_74631[add_74586 > 32'h0000_0009 ? 4'h9 : add_74586[3:0]] + smul_74635;
  assign array_update_74639[0] = add_74586 == 32'h0000_0000 ? add_74637 : array_index_74631[0];
  assign array_update_74639[1] = add_74586 == 32'h0000_0001 ? add_74637 : array_index_74631[1];
  assign array_update_74639[2] = add_74586 == 32'h0000_0002 ? add_74637 : array_index_74631[2];
  assign array_update_74639[3] = add_74586 == 32'h0000_0003 ? add_74637 : array_index_74631[3];
  assign array_update_74639[4] = add_74586 == 32'h0000_0004 ? add_74637 : array_index_74631[4];
  assign array_update_74639[5] = add_74586 == 32'h0000_0005 ? add_74637 : array_index_74631[5];
  assign array_update_74639[6] = add_74586 == 32'h0000_0006 ? add_74637 : array_index_74631[6];
  assign array_update_74639[7] = add_74586 == 32'h0000_0007 ? add_74637 : array_index_74631[7];
  assign array_update_74639[8] = add_74586 == 32'h0000_0008 ? add_74637 : array_index_74631[8];
  assign array_update_74639[9] = add_74586 == 32'h0000_0009 ? add_74637 : array_index_74631[9];
  assign add_74640 = add_74627 + 32'h0000_0001;
  assign array_update_74641[0] = add_73368 == 32'h0000_0000 ? array_update_74639 : array_update_74628[0];
  assign array_update_74641[1] = add_73368 == 32'h0000_0001 ? array_update_74639 : array_update_74628[1];
  assign array_update_74641[2] = add_73368 == 32'h0000_0002 ? array_update_74639 : array_update_74628[2];
  assign array_update_74641[3] = add_73368 == 32'h0000_0003 ? array_update_74639 : array_update_74628[3];
  assign array_update_74641[4] = add_73368 == 32'h0000_0004 ? array_update_74639 : array_update_74628[4];
  assign array_update_74641[5] = add_73368 == 32'h0000_0005 ? array_update_74639 : array_update_74628[5];
  assign array_update_74641[6] = add_73368 == 32'h0000_0006 ? array_update_74639 : array_update_74628[6];
  assign array_update_74641[7] = add_73368 == 32'h0000_0007 ? array_update_74639 : array_update_74628[7];
  assign array_update_74641[8] = add_73368 == 32'h0000_0008 ? array_update_74639 : array_update_74628[8];
  assign array_update_74641[9] = add_73368 == 32'h0000_0009 ? array_update_74639 : array_update_74628[9];
  assign array_index_74643 = array_update_72021[add_74640 > 32'h0000_0009 ? 4'h9 : add_74640[3:0]];
  assign array_index_74644 = array_update_74641[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_74648 = smul32b_32b_x_32b(array_index_73375[add_74640 > 32'h0000_0009 ? 4'h9 : add_74640[3:0]], array_index_74643[add_74586 > 32'h0000_0009 ? 4'h9 : add_74586[3:0]]);
  assign add_74650 = array_index_74644[add_74586 > 32'h0000_0009 ? 4'h9 : add_74586[3:0]] + smul_74648;
  assign array_update_74652[0] = add_74586 == 32'h0000_0000 ? add_74650 : array_index_74644[0];
  assign array_update_74652[1] = add_74586 == 32'h0000_0001 ? add_74650 : array_index_74644[1];
  assign array_update_74652[2] = add_74586 == 32'h0000_0002 ? add_74650 : array_index_74644[2];
  assign array_update_74652[3] = add_74586 == 32'h0000_0003 ? add_74650 : array_index_74644[3];
  assign array_update_74652[4] = add_74586 == 32'h0000_0004 ? add_74650 : array_index_74644[4];
  assign array_update_74652[5] = add_74586 == 32'h0000_0005 ? add_74650 : array_index_74644[5];
  assign array_update_74652[6] = add_74586 == 32'h0000_0006 ? add_74650 : array_index_74644[6];
  assign array_update_74652[7] = add_74586 == 32'h0000_0007 ? add_74650 : array_index_74644[7];
  assign array_update_74652[8] = add_74586 == 32'h0000_0008 ? add_74650 : array_index_74644[8];
  assign array_update_74652[9] = add_74586 == 32'h0000_0009 ? add_74650 : array_index_74644[9];
  assign add_74653 = add_74640 + 32'h0000_0001;
  assign array_update_74654[0] = add_73368 == 32'h0000_0000 ? array_update_74652 : array_update_74641[0];
  assign array_update_74654[1] = add_73368 == 32'h0000_0001 ? array_update_74652 : array_update_74641[1];
  assign array_update_74654[2] = add_73368 == 32'h0000_0002 ? array_update_74652 : array_update_74641[2];
  assign array_update_74654[3] = add_73368 == 32'h0000_0003 ? array_update_74652 : array_update_74641[3];
  assign array_update_74654[4] = add_73368 == 32'h0000_0004 ? array_update_74652 : array_update_74641[4];
  assign array_update_74654[5] = add_73368 == 32'h0000_0005 ? array_update_74652 : array_update_74641[5];
  assign array_update_74654[6] = add_73368 == 32'h0000_0006 ? array_update_74652 : array_update_74641[6];
  assign array_update_74654[7] = add_73368 == 32'h0000_0007 ? array_update_74652 : array_update_74641[7];
  assign array_update_74654[8] = add_73368 == 32'h0000_0008 ? array_update_74652 : array_update_74641[8];
  assign array_update_74654[9] = add_73368 == 32'h0000_0009 ? array_update_74652 : array_update_74641[9];
  assign array_index_74656 = array_update_72021[add_74653 > 32'h0000_0009 ? 4'h9 : add_74653[3:0]];
  assign array_index_74657 = array_update_74654[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_74661 = smul32b_32b_x_32b(array_index_73375[add_74653 > 32'h0000_0009 ? 4'h9 : add_74653[3:0]], array_index_74656[add_74586 > 32'h0000_0009 ? 4'h9 : add_74586[3:0]]);
  assign add_74663 = array_index_74657[add_74586 > 32'h0000_0009 ? 4'h9 : add_74586[3:0]] + smul_74661;
  assign array_update_74665[0] = add_74586 == 32'h0000_0000 ? add_74663 : array_index_74657[0];
  assign array_update_74665[1] = add_74586 == 32'h0000_0001 ? add_74663 : array_index_74657[1];
  assign array_update_74665[2] = add_74586 == 32'h0000_0002 ? add_74663 : array_index_74657[2];
  assign array_update_74665[3] = add_74586 == 32'h0000_0003 ? add_74663 : array_index_74657[3];
  assign array_update_74665[4] = add_74586 == 32'h0000_0004 ? add_74663 : array_index_74657[4];
  assign array_update_74665[5] = add_74586 == 32'h0000_0005 ? add_74663 : array_index_74657[5];
  assign array_update_74665[6] = add_74586 == 32'h0000_0006 ? add_74663 : array_index_74657[6];
  assign array_update_74665[7] = add_74586 == 32'h0000_0007 ? add_74663 : array_index_74657[7];
  assign array_update_74665[8] = add_74586 == 32'h0000_0008 ? add_74663 : array_index_74657[8];
  assign array_update_74665[9] = add_74586 == 32'h0000_0009 ? add_74663 : array_index_74657[9];
  assign add_74666 = add_74653 + 32'h0000_0001;
  assign array_update_74667[0] = add_73368 == 32'h0000_0000 ? array_update_74665 : array_update_74654[0];
  assign array_update_74667[1] = add_73368 == 32'h0000_0001 ? array_update_74665 : array_update_74654[1];
  assign array_update_74667[2] = add_73368 == 32'h0000_0002 ? array_update_74665 : array_update_74654[2];
  assign array_update_74667[3] = add_73368 == 32'h0000_0003 ? array_update_74665 : array_update_74654[3];
  assign array_update_74667[4] = add_73368 == 32'h0000_0004 ? array_update_74665 : array_update_74654[4];
  assign array_update_74667[5] = add_73368 == 32'h0000_0005 ? array_update_74665 : array_update_74654[5];
  assign array_update_74667[6] = add_73368 == 32'h0000_0006 ? array_update_74665 : array_update_74654[6];
  assign array_update_74667[7] = add_73368 == 32'h0000_0007 ? array_update_74665 : array_update_74654[7];
  assign array_update_74667[8] = add_73368 == 32'h0000_0008 ? array_update_74665 : array_update_74654[8];
  assign array_update_74667[9] = add_73368 == 32'h0000_0009 ? array_update_74665 : array_update_74654[9];
  assign array_index_74669 = array_update_72021[add_74666 > 32'h0000_0009 ? 4'h9 : add_74666[3:0]];
  assign array_index_74670 = array_update_74667[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_74674 = smul32b_32b_x_32b(array_index_73375[add_74666 > 32'h0000_0009 ? 4'h9 : add_74666[3:0]], array_index_74669[add_74586 > 32'h0000_0009 ? 4'h9 : add_74586[3:0]]);
  assign add_74676 = array_index_74670[add_74586 > 32'h0000_0009 ? 4'h9 : add_74586[3:0]] + smul_74674;
  assign array_update_74678[0] = add_74586 == 32'h0000_0000 ? add_74676 : array_index_74670[0];
  assign array_update_74678[1] = add_74586 == 32'h0000_0001 ? add_74676 : array_index_74670[1];
  assign array_update_74678[2] = add_74586 == 32'h0000_0002 ? add_74676 : array_index_74670[2];
  assign array_update_74678[3] = add_74586 == 32'h0000_0003 ? add_74676 : array_index_74670[3];
  assign array_update_74678[4] = add_74586 == 32'h0000_0004 ? add_74676 : array_index_74670[4];
  assign array_update_74678[5] = add_74586 == 32'h0000_0005 ? add_74676 : array_index_74670[5];
  assign array_update_74678[6] = add_74586 == 32'h0000_0006 ? add_74676 : array_index_74670[6];
  assign array_update_74678[7] = add_74586 == 32'h0000_0007 ? add_74676 : array_index_74670[7];
  assign array_update_74678[8] = add_74586 == 32'h0000_0008 ? add_74676 : array_index_74670[8];
  assign array_update_74678[9] = add_74586 == 32'h0000_0009 ? add_74676 : array_index_74670[9];
  assign add_74679 = add_74666 + 32'h0000_0001;
  assign array_update_74680[0] = add_73368 == 32'h0000_0000 ? array_update_74678 : array_update_74667[0];
  assign array_update_74680[1] = add_73368 == 32'h0000_0001 ? array_update_74678 : array_update_74667[1];
  assign array_update_74680[2] = add_73368 == 32'h0000_0002 ? array_update_74678 : array_update_74667[2];
  assign array_update_74680[3] = add_73368 == 32'h0000_0003 ? array_update_74678 : array_update_74667[3];
  assign array_update_74680[4] = add_73368 == 32'h0000_0004 ? array_update_74678 : array_update_74667[4];
  assign array_update_74680[5] = add_73368 == 32'h0000_0005 ? array_update_74678 : array_update_74667[5];
  assign array_update_74680[6] = add_73368 == 32'h0000_0006 ? array_update_74678 : array_update_74667[6];
  assign array_update_74680[7] = add_73368 == 32'h0000_0007 ? array_update_74678 : array_update_74667[7];
  assign array_update_74680[8] = add_73368 == 32'h0000_0008 ? array_update_74678 : array_update_74667[8];
  assign array_update_74680[9] = add_73368 == 32'h0000_0009 ? array_update_74678 : array_update_74667[9];
  assign array_index_74682 = array_update_72021[add_74679 > 32'h0000_0009 ? 4'h9 : add_74679[3:0]];
  assign array_index_74683 = array_update_74680[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_74687 = smul32b_32b_x_32b(array_index_73375[add_74679 > 32'h0000_0009 ? 4'h9 : add_74679[3:0]], array_index_74682[add_74586 > 32'h0000_0009 ? 4'h9 : add_74586[3:0]]);
  assign add_74689 = array_index_74683[add_74586 > 32'h0000_0009 ? 4'h9 : add_74586[3:0]] + smul_74687;
  assign array_update_74691[0] = add_74586 == 32'h0000_0000 ? add_74689 : array_index_74683[0];
  assign array_update_74691[1] = add_74586 == 32'h0000_0001 ? add_74689 : array_index_74683[1];
  assign array_update_74691[2] = add_74586 == 32'h0000_0002 ? add_74689 : array_index_74683[2];
  assign array_update_74691[3] = add_74586 == 32'h0000_0003 ? add_74689 : array_index_74683[3];
  assign array_update_74691[4] = add_74586 == 32'h0000_0004 ? add_74689 : array_index_74683[4];
  assign array_update_74691[5] = add_74586 == 32'h0000_0005 ? add_74689 : array_index_74683[5];
  assign array_update_74691[6] = add_74586 == 32'h0000_0006 ? add_74689 : array_index_74683[6];
  assign array_update_74691[7] = add_74586 == 32'h0000_0007 ? add_74689 : array_index_74683[7];
  assign array_update_74691[8] = add_74586 == 32'h0000_0008 ? add_74689 : array_index_74683[8];
  assign array_update_74691[9] = add_74586 == 32'h0000_0009 ? add_74689 : array_index_74683[9];
  assign add_74692 = add_74679 + 32'h0000_0001;
  assign array_update_74693[0] = add_73368 == 32'h0000_0000 ? array_update_74691 : array_update_74680[0];
  assign array_update_74693[1] = add_73368 == 32'h0000_0001 ? array_update_74691 : array_update_74680[1];
  assign array_update_74693[2] = add_73368 == 32'h0000_0002 ? array_update_74691 : array_update_74680[2];
  assign array_update_74693[3] = add_73368 == 32'h0000_0003 ? array_update_74691 : array_update_74680[3];
  assign array_update_74693[4] = add_73368 == 32'h0000_0004 ? array_update_74691 : array_update_74680[4];
  assign array_update_74693[5] = add_73368 == 32'h0000_0005 ? array_update_74691 : array_update_74680[5];
  assign array_update_74693[6] = add_73368 == 32'h0000_0006 ? array_update_74691 : array_update_74680[6];
  assign array_update_74693[7] = add_73368 == 32'h0000_0007 ? array_update_74691 : array_update_74680[7];
  assign array_update_74693[8] = add_73368 == 32'h0000_0008 ? array_update_74691 : array_update_74680[8];
  assign array_update_74693[9] = add_73368 == 32'h0000_0009 ? array_update_74691 : array_update_74680[9];
  assign array_index_74695 = array_update_72021[add_74692 > 32'h0000_0009 ? 4'h9 : add_74692[3:0]];
  assign array_index_74696 = array_update_74693[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_74700 = smul32b_32b_x_32b(array_index_73375[add_74692 > 32'h0000_0009 ? 4'h9 : add_74692[3:0]], array_index_74695[add_74586 > 32'h0000_0009 ? 4'h9 : add_74586[3:0]]);
  assign add_74702 = array_index_74696[add_74586 > 32'h0000_0009 ? 4'h9 : add_74586[3:0]] + smul_74700;
  assign array_update_74704[0] = add_74586 == 32'h0000_0000 ? add_74702 : array_index_74696[0];
  assign array_update_74704[1] = add_74586 == 32'h0000_0001 ? add_74702 : array_index_74696[1];
  assign array_update_74704[2] = add_74586 == 32'h0000_0002 ? add_74702 : array_index_74696[2];
  assign array_update_74704[3] = add_74586 == 32'h0000_0003 ? add_74702 : array_index_74696[3];
  assign array_update_74704[4] = add_74586 == 32'h0000_0004 ? add_74702 : array_index_74696[4];
  assign array_update_74704[5] = add_74586 == 32'h0000_0005 ? add_74702 : array_index_74696[5];
  assign array_update_74704[6] = add_74586 == 32'h0000_0006 ? add_74702 : array_index_74696[6];
  assign array_update_74704[7] = add_74586 == 32'h0000_0007 ? add_74702 : array_index_74696[7];
  assign array_update_74704[8] = add_74586 == 32'h0000_0008 ? add_74702 : array_index_74696[8];
  assign array_update_74704[9] = add_74586 == 32'h0000_0009 ? add_74702 : array_index_74696[9];
  assign add_74705 = add_74692 + 32'h0000_0001;
  assign array_update_74706[0] = add_73368 == 32'h0000_0000 ? array_update_74704 : array_update_74693[0];
  assign array_update_74706[1] = add_73368 == 32'h0000_0001 ? array_update_74704 : array_update_74693[1];
  assign array_update_74706[2] = add_73368 == 32'h0000_0002 ? array_update_74704 : array_update_74693[2];
  assign array_update_74706[3] = add_73368 == 32'h0000_0003 ? array_update_74704 : array_update_74693[3];
  assign array_update_74706[4] = add_73368 == 32'h0000_0004 ? array_update_74704 : array_update_74693[4];
  assign array_update_74706[5] = add_73368 == 32'h0000_0005 ? array_update_74704 : array_update_74693[5];
  assign array_update_74706[6] = add_73368 == 32'h0000_0006 ? array_update_74704 : array_update_74693[6];
  assign array_update_74706[7] = add_73368 == 32'h0000_0007 ? array_update_74704 : array_update_74693[7];
  assign array_update_74706[8] = add_73368 == 32'h0000_0008 ? array_update_74704 : array_update_74693[8];
  assign array_update_74706[9] = add_73368 == 32'h0000_0009 ? array_update_74704 : array_update_74693[9];
  assign array_index_74708 = array_update_72021[add_74705 > 32'h0000_0009 ? 4'h9 : add_74705[3:0]];
  assign array_index_74709 = array_update_74706[add_73368 > 32'h0000_0009 ? 4'h9 : add_73368[3:0]];
  assign smul_74713 = smul32b_32b_x_32b(array_index_73375[add_74705 > 32'h0000_0009 ? 4'h9 : add_74705[3:0]], array_index_74708[add_74586 > 32'h0000_0009 ? 4'h9 : add_74586[3:0]]);
  assign add_74715 = array_index_74709[add_74586 > 32'h0000_0009 ? 4'h9 : add_74586[3:0]] + smul_74713;
  assign array_update_74716[0] = add_74586 == 32'h0000_0000 ? add_74715 : array_index_74709[0];
  assign array_update_74716[1] = add_74586 == 32'h0000_0001 ? add_74715 : array_index_74709[1];
  assign array_update_74716[2] = add_74586 == 32'h0000_0002 ? add_74715 : array_index_74709[2];
  assign array_update_74716[3] = add_74586 == 32'h0000_0003 ? add_74715 : array_index_74709[3];
  assign array_update_74716[4] = add_74586 == 32'h0000_0004 ? add_74715 : array_index_74709[4];
  assign array_update_74716[5] = add_74586 == 32'h0000_0005 ? add_74715 : array_index_74709[5];
  assign array_update_74716[6] = add_74586 == 32'h0000_0006 ? add_74715 : array_index_74709[6];
  assign array_update_74716[7] = add_74586 == 32'h0000_0007 ? add_74715 : array_index_74709[7];
  assign array_update_74716[8] = add_74586 == 32'h0000_0008 ? add_74715 : array_index_74709[8];
  assign array_update_74716[9] = add_74586 == 32'h0000_0009 ? add_74715 : array_index_74709[9];
  assign array_update_74718[0] = add_73368 == 32'h0000_0000 ? array_update_74716 : array_update_74706[0];
  assign array_update_74718[1] = add_73368 == 32'h0000_0001 ? array_update_74716 : array_update_74706[1];
  assign array_update_74718[2] = add_73368 == 32'h0000_0002 ? array_update_74716 : array_update_74706[2];
  assign array_update_74718[3] = add_73368 == 32'h0000_0003 ? array_update_74716 : array_update_74706[3];
  assign array_update_74718[4] = add_73368 == 32'h0000_0004 ? array_update_74716 : array_update_74706[4];
  assign array_update_74718[5] = add_73368 == 32'h0000_0005 ? array_update_74716 : array_update_74706[5];
  assign array_update_74718[6] = add_73368 == 32'h0000_0006 ? array_update_74716 : array_update_74706[6];
  assign array_update_74718[7] = add_73368 == 32'h0000_0007 ? array_update_74716 : array_update_74706[7];
  assign array_update_74718[8] = add_73368 == 32'h0000_0008 ? array_update_74716 : array_update_74706[8];
  assign array_update_74718[9] = add_73368 == 32'h0000_0009 ? array_update_74716 : array_update_74706[9];
  assign add_74719 = add_73368 + 32'h0000_0001;
  assign array_index_74720 = array_update_74718[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign literal_74722 = 32'h0000_0000;
  assign array_update_74723[0] = literal_74722 == 32'h0000_0000 ? 32'h0000_0000 : array_index_74720[0];
  assign array_update_74723[1] = literal_74722 == 32'h0000_0001 ? 32'h0000_0000 : array_index_74720[1];
  assign array_update_74723[2] = literal_74722 == 32'h0000_0002 ? 32'h0000_0000 : array_index_74720[2];
  assign array_update_74723[3] = literal_74722 == 32'h0000_0003 ? 32'h0000_0000 : array_index_74720[3];
  assign array_update_74723[4] = literal_74722 == 32'h0000_0004 ? 32'h0000_0000 : array_index_74720[4];
  assign array_update_74723[5] = literal_74722 == 32'h0000_0005 ? 32'h0000_0000 : array_index_74720[5];
  assign array_update_74723[6] = literal_74722 == 32'h0000_0006 ? 32'h0000_0000 : array_index_74720[6];
  assign array_update_74723[7] = literal_74722 == 32'h0000_0007 ? 32'h0000_0000 : array_index_74720[7];
  assign array_update_74723[8] = literal_74722 == 32'h0000_0008 ? 32'h0000_0000 : array_index_74720[8];
  assign array_update_74723[9] = literal_74722 == 32'h0000_0009 ? 32'h0000_0000 : array_index_74720[9];
  assign literal_74724 = 32'h0000_0000;
  assign array_update_74725[0] = add_74719 == 32'h0000_0000 ? array_update_74723 : array_update_74718[0];
  assign array_update_74725[1] = add_74719 == 32'h0000_0001 ? array_update_74723 : array_update_74718[1];
  assign array_update_74725[2] = add_74719 == 32'h0000_0002 ? array_update_74723 : array_update_74718[2];
  assign array_update_74725[3] = add_74719 == 32'h0000_0003 ? array_update_74723 : array_update_74718[3];
  assign array_update_74725[4] = add_74719 == 32'h0000_0004 ? array_update_74723 : array_update_74718[4];
  assign array_update_74725[5] = add_74719 == 32'h0000_0005 ? array_update_74723 : array_update_74718[5];
  assign array_update_74725[6] = add_74719 == 32'h0000_0006 ? array_update_74723 : array_update_74718[6];
  assign array_update_74725[7] = add_74719 == 32'h0000_0007 ? array_update_74723 : array_update_74718[7];
  assign array_update_74725[8] = add_74719 == 32'h0000_0008 ? array_update_74723 : array_update_74718[8];
  assign array_update_74725[9] = add_74719 == 32'h0000_0009 ? array_update_74723 : array_update_74718[9];
  assign array_index_74726 = array_update_72020[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign array_index_74727 = array_update_72021[literal_74724 > 32'h0000_0009 ? 4'h9 : literal_74724[3:0]];
  assign array_index_74728 = array_update_74725[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_74732 = smul32b_32b_x_32b(array_index_74726[literal_74724 > 32'h0000_0009 ? 4'h9 : literal_74724[3:0]], array_index_74727[literal_74722 > 32'h0000_0009 ? 4'h9 : literal_74722[3:0]]);
  assign add_74734 = array_index_74728[literal_74722 > 32'h0000_0009 ? 4'h9 : literal_74722[3:0]] + smul_74732;
  assign array_update_74736[0] = literal_74722 == 32'h0000_0000 ? add_74734 : array_index_74728[0];
  assign array_update_74736[1] = literal_74722 == 32'h0000_0001 ? add_74734 : array_index_74728[1];
  assign array_update_74736[2] = literal_74722 == 32'h0000_0002 ? add_74734 : array_index_74728[2];
  assign array_update_74736[3] = literal_74722 == 32'h0000_0003 ? add_74734 : array_index_74728[3];
  assign array_update_74736[4] = literal_74722 == 32'h0000_0004 ? add_74734 : array_index_74728[4];
  assign array_update_74736[5] = literal_74722 == 32'h0000_0005 ? add_74734 : array_index_74728[5];
  assign array_update_74736[6] = literal_74722 == 32'h0000_0006 ? add_74734 : array_index_74728[6];
  assign array_update_74736[7] = literal_74722 == 32'h0000_0007 ? add_74734 : array_index_74728[7];
  assign array_update_74736[8] = literal_74722 == 32'h0000_0008 ? add_74734 : array_index_74728[8];
  assign array_update_74736[9] = literal_74722 == 32'h0000_0009 ? add_74734 : array_index_74728[9];
  assign add_74737 = literal_74724 + 32'h0000_0001;
  assign array_update_74738[0] = add_74719 == 32'h0000_0000 ? array_update_74736 : array_update_74725[0];
  assign array_update_74738[1] = add_74719 == 32'h0000_0001 ? array_update_74736 : array_update_74725[1];
  assign array_update_74738[2] = add_74719 == 32'h0000_0002 ? array_update_74736 : array_update_74725[2];
  assign array_update_74738[3] = add_74719 == 32'h0000_0003 ? array_update_74736 : array_update_74725[3];
  assign array_update_74738[4] = add_74719 == 32'h0000_0004 ? array_update_74736 : array_update_74725[4];
  assign array_update_74738[5] = add_74719 == 32'h0000_0005 ? array_update_74736 : array_update_74725[5];
  assign array_update_74738[6] = add_74719 == 32'h0000_0006 ? array_update_74736 : array_update_74725[6];
  assign array_update_74738[7] = add_74719 == 32'h0000_0007 ? array_update_74736 : array_update_74725[7];
  assign array_update_74738[8] = add_74719 == 32'h0000_0008 ? array_update_74736 : array_update_74725[8];
  assign array_update_74738[9] = add_74719 == 32'h0000_0009 ? array_update_74736 : array_update_74725[9];
  assign array_index_74740 = array_update_72021[add_74737 > 32'h0000_0009 ? 4'h9 : add_74737[3:0]];
  assign array_index_74741 = array_update_74738[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_74745 = smul32b_32b_x_32b(array_index_74726[add_74737 > 32'h0000_0009 ? 4'h9 : add_74737[3:0]], array_index_74740[literal_74722 > 32'h0000_0009 ? 4'h9 : literal_74722[3:0]]);
  assign add_74747 = array_index_74741[literal_74722 > 32'h0000_0009 ? 4'h9 : literal_74722[3:0]] + smul_74745;
  assign array_update_74749[0] = literal_74722 == 32'h0000_0000 ? add_74747 : array_index_74741[0];
  assign array_update_74749[1] = literal_74722 == 32'h0000_0001 ? add_74747 : array_index_74741[1];
  assign array_update_74749[2] = literal_74722 == 32'h0000_0002 ? add_74747 : array_index_74741[2];
  assign array_update_74749[3] = literal_74722 == 32'h0000_0003 ? add_74747 : array_index_74741[3];
  assign array_update_74749[4] = literal_74722 == 32'h0000_0004 ? add_74747 : array_index_74741[4];
  assign array_update_74749[5] = literal_74722 == 32'h0000_0005 ? add_74747 : array_index_74741[5];
  assign array_update_74749[6] = literal_74722 == 32'h0000_0006 ? add_74747 : array_index_74741[6];
  assign array_update_74749[7] = literal_74722 == 32'h0000_0007 ? add_74747 : array_index_74741[7];
  assign array_update_74749[8] = literal_74722 == 32'h0000_0008 ? add_74747 : array_index_74741[8];
  assign array_update_74749[9] = literal_74722 == 32'h0000_0009 ? add_74747 : array_index_74741[9];
  assign add_74750 = add_74737 + 32'h0000_0001;
  assign array_update_74751[0] = add_74719 == 32'h0000_0000 ? array_update_74749 : array_update_74738[0];
  assign array_update_74751[1] = add_74719 == 32'h0000_0001 ? array_update_74749 : array_update_74738[1];
  assign array_update_74751[2] = add_74719 == 32'h0000_0002 ? array_update_74749 : array_update_74738[2];
  assign array_update_74751[3] = add_74719 == 32'h0000_0003 ? array_update_74749 : array_update_74738[3];
  assign array_update_74751[4] = add_74719 == 32'h0000_0004 ? array_update_74749 : array_update_74738[4];
  assign array_update_74751[5] = add_74719 == 32'h0000_0005 ? array_update_74749 : array_update_74738[5];
  assign array_update_74751[6] = add_74719 == 32'h0000_0006 ? array_update_74749 : array_update_74738[6];
  assign array_update_74751[7] = add_74719 == 32'h0000_0007 ? array_update_74749 : array_update_74738[7];
  assign array_update_74751[8] = add_74719 == 32'h0000_0008 ? array_update_74749 : array_update_74738[8];
  assign array_update_74751[9] = add_74719 == 32'h0000_0009 ? array_update_74749 : array_update_74738[9];
  assign array_index_74753 = array_update_72021[add_74750 > 32'h0000_0009 ? 4'h9 : add_74750[3:0]];
  assign array_index_74754 = array_update_74751[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_74758 = smul32b_32b_x_32b(array_index_74726[add_74750 > 32'h0000_0009 ? 4'h9 : add_74750[3:0]], array_index_74753[literal_74722 > 32'h0000_0009 ? 4'h9 : literal_74722[3:0]]);
  assign add_74760 = array_index_74754[literal_74722 > 32'h0000_0009 ? 4'h9 : literal_74722[3:0]] + smul_74758;
  assign array_update_74762[0] = literal_74722 == 32'h0000_0000 ? add_74760 : array_index_74754[0];
  assign array_update_74762[1] = literal_74722 == 32'h0000_0001 ? add_74760 : array_index_74754[1];
  assign array_update_74762[2] = literal_74722 == 32'h0000_0002 ? add_74760 : array_index_74754[2];
  assign array_update_74762[3] = literal_74722 == 32'h0000_0003 ? add_74760 : array_index_74754[3];
  assign array_update_74762[4] = literal_74722 == 32'h0000_0004 ? add_74760 : array_index_74754[4];
  assign array_update_74762[5] = literal_74722 == 32'h0000_0005 ? add_74760 : array_index_74754[5];
  assign array_update_74762[6] = literal_74722 == 32'h0000_0006 ? add_74760 : array_index_74754[6];
  assign array_update_74762[7] = literal_74722 == 32'h0000_0007 ? add_74760 : array_index_74754[7];
  assign array_update_74762[8] = literal_74722 == 32'h0000_0008 ? add_74760 : array_index_74754[8];
  assign array_update_74762[9] = literal_74722 == 32'h0000_0009 ? add_74760 : array_index_74754[9];
  assign add_74763 = add_74750 + 32'h0000_0001;
  assign array_update_74764[0] = add_74719 == 32'h0000_0000 ? array_update_74762 : array_update_74751[0];
  assign array_update_74764[1] = add_74719 == 32'h0000_0001 ? array_update_74762 : array_update_74751[1];
  assign array_update_74764[2] = add_74719 == 32'h0000_0002 ? array_update_74762 : array_update_74751[2];
  assign array_update_74764[3] = add_74719 == 32'h0000_0003 ? array_update_74762 : array_update_74751[3];
  assign array_update_74764[4] = add_74719 == 32'h0000_0004 ? array_update_74762 : array_update_74751[4];
  assign array_update_74764[5] = add_74719 == 32'h0000_0005 ? array_update_74762 : array_update_74751[5];
  assign array_update_74764[6] = add_74719 == 32'h0000_0006 ? array_update_74762 : array_update_74751[6];
  assign array_update_74764[7] = add_74719 == 32'h0000_0007 ? array_update_74762 : array_update_74751[7];
  assign array_update_74764[8] = add_74719 == 32'h0000_0008 ? array_update_74762 : array_update_74751[8];
  assign array_update_74764[9] = add_74719 == 32'h0000_0009 ? array_update_74762 : array_update_74751[9];
  assign array_index_74766 = array_update_72021[add_74763 > 32'h0000_0009 ? 4'h9 : add_74763[3:0]];
  assign array_index_74767 = array_update_74764[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_74771 = smul32b_32b_x_32b(array_index_74726[add_74763 > 32'h0000_0009 ? 4'h9 : add_74763[3:0]], array_index_74766[literal_74722 > 32'h0000_0009 ? 4'h9 : literal_74722[3:0]]);
  assign add_74773 = array_index_74767[literal_74722 > 32'h0000_0009 ? 4'h9 : literal_74722[3:0]] + smul_74771;
  assign array_update_74775[0] = literal_74722 == 32'h0000_0000 ? add_74773 : array_index_74767[0];
  assign array_update_74775[1] = literal_74722 == 32'h0000_0001 ? add_74773 : array_index_74767[1];
  assign array_update_74775[2] = literal_74722 == 32'h0000_0002 ? add_74773 : array_index_74767[2];
  assign array_update_74775[3] = literal_74722 == 32'h0000_0003 ? add_74773 : array_index_74767[3];
  assign array_update_74775[4] = literal_74722 == 32'h0000_0004 ? add_74773 : array_index_74767[4];
  assign array_update_74775[5] = literal_74722 == 32'h0000_0005 ? add_74773 : array_index_74767[5];
  assign array_update_74775[6] = literal_74722 == 32'h0000_0006 ? add_74773 : array_index_74767[6];
  assign array_update_74775[7] = literal_74722 == 32'h0000_0007 ? add_74773 : array_index_74767[7];
  assign array_update_74775[8] = literal_74722 == 32'h0000_0008 ? add_74773 : array_index_74767[8];
  assign array_update_74775[9] = literal_74722 == 32'h0000_0009 ? add_74773 : array_index_74767[9];
  assign add_74776 = add_74763 + 32'h0000_0001;
  assign array_update_74777[0] = add_74719 == 32'h0000_0000 ? array_update_74775 : array_update_74764[0];
  assign array_update_74777[1] = add_74719 == 32'h0000_0001 ? array_update_74775 : array_update_74764[1];
  assign array_update_74777[2] = add_74719 == 32'h0000_0002 ? array_update_74775 : array_update_74764[2];
  assign array_update_74777[3] = add_74719 == 32'h0000_0003 ? array_update_74775 : array_update_74764[3];
  assign array_update_74777[4] = add_74719 == 32'h0000_0004 ? array_update_74775 : array_update_74764[4];
  assign array_update_74777[5] = add_74719 == 32'h0000_0005 ? array_update_74775 : array_update_74764[5];
  assign array_update_74777[6] = add_74719 == 32'h0000_0006 ? array_update_74775 : array_update_74764[6];
  assign array_update_74777[7] = add_74719 == 32'h0000_0007 ? array_update_74775 : array_update_74764[7];
  assign array_update_74777[8] = add_74719 == 32'h0000_0008 ? array_update_74775 : array_update_74764[8];
  assign array_update_74777[9] = add_74719 == 32'h0000_0009 ? array_update_74775 : array_update_74764[9];
  assign array_index_74779 = array_update_72021[add_74776 > 32'h0000_0009 ? 4'h9 : add_74776[3:0]];
  assign array_index_74780 = array_update_74777[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_74784 = smul32b_32b_x_32b(array_index_74726[add_74776 > 32'h0000_0009 ? 4'h9 : add_74776[3:0]], array_index_74779[literal_74722 > 32'h0000_0009 ? 4'h9 : literal_74722[3:0]]);
  assign add_74786 = array_index_74780[literal_74722 > 32'h0000_0009 ? 4'h9 : literal_74722[3:0]] + smul_74784;
  assign array_update_74788[0] = literal_74722 == 32'h0000_0000 ? add_74786 : array_index_74780[0];
  assign array_update_74788[1] = literal_74722 == 32'h0000_0001 ? add_74786 : array_index_74780[1];
  assign array_update_74788[2] = literal_74722 == 32'h0000_0002 ? add_74786 : array_index_74780[2];
  assign array_update_74788[3] = literal_74722 == 32'h0000_0003 ? add_74786 : array_index_74780[3];
  assign array_update_74788[4] = literal_74722 == 32'h0000_0004 ? add_74786 : array_index_74780[4];
  assign array_update_74788[5] = literal_74722 == 32'h0000_0005 ? add_74786 : array_index_74780[5];
  assign array_update_74788[6] = literal_74722 == 32'h0000_0006 ? add_74786 : array_index_74780[6];
  assign array_update_74788[7] = literal_74722 == 32'h0000_0007 ? add_74786 : array_index_74780[7];
  assign array_update_74788[8] = literal_74722 == 32'h0000_0008 ? add_74786 : array_index_74780[8];
  assign array_update_74788[9] = literal_74722 == 32'h0000_0009 ? add_74786 : array_index_74780[9];
  assign add_74789 = add_74776 + 32'h0000_0001;
  assign array_update_74790[0] = add_74719 == 32'h0000_0000 ? array_update_74788 : array_update_74777[0];
  assign array_update_74790[1] = add_74719 == 32'h0000_0001 ? array_update_74788 : array_update_74777[1];
  assign array_update_74790[2] = add_74719 == 32'h0000_0002 ? array_update_74788 : array_update_74777[2];
  assign array_update_74790[3] = add_74719 == 32'h0000_0003 ? array_update_74788 : array_update_74777[3];
  assign array_update_74790[4] = add_74719 == 32'h0000_0004 ? array_update_74788 : array_update_74777[4];
  assign array_update_74790[5] = add_74719 == 32'h0000_0005 ? array_update_74788 : array_update_74777[5];
  assign array_update_74790[6] = add_74719 == 32'h0000_0006 ? array_update_74788 : array_update_74777[6];
  assign array_update_74790[7] = add_74719 == 32'h0000_0007 ? array_update_74788 : array_update_74777[7];
  assign array_update_74790[8] = add_74719 == 32'h0000_0008 ? array_update_74788 : array_update_74777[8];
  assign array_update_74790[9] = add_74719 == 32'h0000_0009 ? array_update_74788 : array_update_74777[9];
  assign array_index_74792 = array_update_72021[add_74789 > 32'h0000_0009 ? 4'h9 : add_74789[3:0]];
  assign array_index_74793 = array_update_74790[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_74797 = smul32b_32b_x_32b(array_index_74726[add_74789 > 32'h0000_0009 ? 4'h9 : add_74789[3:0]], array_index_74792[literal_74722 > 32'h0000_0009 ? 4'h9 : literal_74722[3:0]]);
  assign add_74799 = array_index_74793[literal_74722 > 32'h0000_0009 ? 4'h9 : literal_74722[3:0]] + smul_74797;
  assign array_update_74801[0] = literal_74722 == 32'h0000_0000 ? add_74799 : array_index_74793[0];
  assign array_update_74801[1] = literal_74722 == 32'h0000_0001 ? add_74799 : array_index_74793[1];
  assign array_update_74801[2] = literal_74722 == 32'h0000_0002 ? add_74799 : array_index_74793[2];
  assign array_update_74801[3] = literal_74722 == 32'h0000_0003 ? add_74799 : array_index_74793[3];
  assign array_update_74801[4] = literal_74722 == 32'h0000_0004 ? add_74799 : array_index_74793[4];
  assign array_update_74801[5] = literal_74722 == 32'h0000_0005 ? add_74799 : array_index_74793[5];
  assign array_update_74801[6] = literal_74722 == 32'h0000_0006 ? add_74799 : array_index_74793[6];
  assign array_update_74801[7] = literal_74722 == 32'h0000_0007 ? add_74799 : array_index_74793[7];
  assign array_update_74801[8] = literal_74722 == 32'h0000_0008 ? add_74799 : array_index_74793[8];
  assign array_update_74801[9] = literal_74722 == 32'h0000_0009 ? add_74799 : array_index_74793[9];
  assign add_74802 = add_74789 + 32'h0000_0001;
  assign array_update_74803[0] = add_74719 == 32'h0000_0000 ? array_update_74801 : array_update_74790[0];
  assign array_update_74803[1] = add_74719 == 32'h0000_0001 ? array_update_74801 : array_update_74790[1];
  assign array_update_74803[2] = add_74719 == 32'h0000_0002 ? array_update_74801 : array_update_74790[2];
  assign array_update_74803[3] = add_74719 == 32'h0000_0003 ? array_update_74801 : array_update_74790[3];
  assign array_update_74803[4] = add_74719 == 32'h0000_0004 ? array_update_74801 : array_update_74790[4];
  assign array_update_74803[5] = add_74719 == 32'h0000_0005 ? array_update_74801 : array_update_74790[5];
  assign array_update_74803[6] = add_74719 == 32'h0000_0006 ? array_update_74801 : array_update_74790[6];
  assign array_update_74803[7] = add_74719 == 32'h0000_0007 ? array_update_74801 : array_update_74790[7];
  assign array_update_74803[8] = add_74719 == 32'h0000_0008 ? array_update_74801 : array_update_74790[8];
  assign array_update_74803[9] = add_74719 == 32'h0000_0009 ? array_update_74801 : array_update_74790[9];
  assign array_index_74805 = array_update_72021[add_74802 > 32'h0000_0009 ? 4'h9 : add_74802[3:0]];
  assign array_index_74806 = array_update_74803[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_74810 = smul32b_32b_x_32b(array_index_74726[add_74802 > 32'h0000_0009 ? 4'h9 : add_74802[3:0]], array_index_74805[literal_74722 > 32'h0000_0009 ? 4'h9 : literal_74722[3:0]]);
  assign add_74812 = array_index_74806[literal_74722 > 32'h0000_0009 ? 4'h9 : literal_74722[3:0]] + smul_74810;
  assign array_update_74814[0] = literal_74722 == 32'h0000_0000 ? add_74812 : array_index_74806[0];
  assign array_update_74814[1] = literal_74722 == 32'h0000_0001 ? add_74812 : array_index_74806[1];
  assign array_update_74814[2] = literal_74722 == 32'h0000_0002 ? add_74812 : array_index_74806[2];
  assign array_update_74814[3] = literal_74722 == 32'h0000_0003 ? add_74812 : array_index_74806[3];
  assign array_update_74814[4] = literal_74722 == 32'h0000_0004 ? add_74812 : array_index_74806[4];
  assign array_update_74814[5] = literal_74722 == 32'h0000_0005 ? add_74812 : array_index_74806[5];
  assign array_update_74814[6] = literal_74722 == 32'h0000_0006 ? add_74812 : array_index_74806[6];
  assign array_update_74814[7] = literal_74722 == 32'h0000_0007 ? add_74812 : array_index_74806[7];
  assign array_update_74814[8] = literal_74722 == 32'h0000_0008 ? add_74812 : array_index_74806[8];
  assign array_update_74814[9] = literal_74722 == 32'h0000_0009 ? add_74812 : array_index_74806[9];
  assign add_74815 = add_74802 + 32'h0000_0001;
  assign array_update_74816[0] = add_74719 == 32'h0000_0000 ? array_update_74814 : array_update_74803[0];
  assign array_update_74816[1] = add_74719 == 32'h0000_0001 ? array_update_74814 : array_update_74803[1];
  assign array_update_74816[2] = add_74719 == 32'h0000_0002 ? array_update_74814 : array_update_74803[2];
  assign array_update_74816[3] = add_74719 == 32'h0000_0003 ? array_update_74814 : array_update_74803[3];
  assign array_update_74816[4] = add_74719 == 32'h0000_0004 ? array_update_74814 : array_update_74803[4];
  assign array_update_74816[5] = add_74719 == 32'h0000_0005 ? array_update_74814 : array_update_74803[5];
  assign array_update_74816[6] = add_74719 == 32'h0000_0006 ? array_update_74814 : array_update_74803[6];
  assign array_update_74816[7] = add_74719 == 32'h0000_0007 ? array_update_74814 : array_update_74803[7];
  assign array_update_74816[8] = add_74719 == 32'h0000_0008 ? array_update_74814 : array_update_74803[8];
  assign array_update_74816[9] = add_74719 == 32'h0000_0009 ? array_update_74814 : array_update_74803[9];
  assign array_index_74818 = array_update_72021[add_74815 > 32'h0000_0009 ? 4'h9 : add_74815[3:0]];
  assign array_index_74819 = array_update_74816[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_74823 = smul32b_32b_x_32b(array_index_74726[add_74815 > 32'h0000_0009 ? 4'h9 : add_74815[3:0]], array_index_74818[literal_74722 > 32'h0000_0009 ? 4'h9 : literal_74722[3:0]]);
  assign add_74825 = array_index_74819[literal_74722 > 32'h0000_0009 ? 4'h9 : literal_74722[3:0]] + smul_74823;
  assign array_update_74827[0] = literal_74722 == 32'h0000_0000 ? add_74825 : array_index_74819[0];
  assign array_update_74827[1] = literal_74722 == 32'h0000_0001 ? add_74825 : array_index_74819[1];
  assign array_update_74827[2] = literal_74722 == 32'h0000_0002 ? add_74825 : array_index_74819[2];
  assign array_update_74827[3] = literal_74722 == 32'h0000_0003 ? add_74825 : array_index_74819[3];
  assign array_update_74827[4] = literal_74722 == 32'h0000_0004 ? add_74825 : array_index_74819[4];
  assign array_update_74827[5] = literal_74722 == 32'h0000_0005 ? add_74825 : array_index_74819[5];
  assign array_update_74827[6] = literal_74722 == 32'h0000_0006 ? add_74825 : array_index_74819[6];
  assign array_update_74827[7] = literal_74722 == 32'h0000_0007 ? add_74825 : array_index_74819[7];
  assign array_update_74827[8] = literal_74722 == 32'h0000_0008 ? add_74825 : array_index_74819[8];
  assign array_update_74827[9] = literal_74722 == 32'h0000_0009 ? add_74825 : array_index_74819[9];
  assign add_74828 = add_74815 + 32'h0000_0001;
  assign array_update_74829[0] = add_74719 == 32'h0000_0000 ? array_update_74827 : array_update_74816[0];
  assign array_update_74829[1] = add_74719 == 32'h0000_0001 ? array_update_74827 : array_update_74816[1];
  assign array_update_74829[2] = add_74719 == 32'h0000_0002 ? array_update_74827 : array_update_74816[2];
  assign array_update_74829[3] = add_74719 == 32'h0000_0003 ? array_update_74827 : array_update_74816[3];
  assign array_update_74829[4] = add_74719 == 32'h0000_0004 ? array_update_74827 : array_update_74816[4];
  assign array_update_74829[5] = add_74719 == 32'h0000_0005 ? array_update_74827 : array_update_74816[5];
  assign array_update_74829[6] = add_74719 == 32'h0000_0006 ? array_update_74827 : array_update_74816[6];
  assign array_update_74829[7] = add_74719 == 32'h0000_0007 ? array_update_74827 : array_update_74816[7];
  assign array_update_74829[8] = add_74719 == 32'h0000_0008 ? array_update_74827 : array_update_74816[8];
  assign array_update_74829[9] = add_74719 == 32'h0000_0009 ? array_update_74827 : array_update_74816[9];
  assign array_index_74831 = array_update_72021[add_74828 > 32'h0000_0009 ? 4'h9 : add_74828[3:0]];
  assign array_index_74832 = array_update_74829[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_74836 = smul32b_32b_x_32b(array_index_74726[add_74828 > 32'h0000_0009 ? 4'h9 : add_74828[3:0]], array_index_74831[literal_74722 > 32'h0000_0009 ? 4'h9 : literal_74722[3:0]]);
  assign add_74838 = array_index_74832[literal_74722 > 32'h0000_0009 ? 4'h9 : literal_74722[3:0]] + smul_74836;
  assign array_update_74840[0] = literal_74722 == 32'h0000_0000 ? add_74838 : array_index_74832[0];
  assign array_update_74840[1] = literal_74722 == 32'h0000_0001 ? add_74838 : array_index_74832[1];
  assign array_update_74840[2] = literal_74722 == 32'h0000_0002 ? add_74838 : array_index_74832[2];
  assign array_update_74840[3] = literal_74722 == 32'h0000_0003 ? add_74838 : array_index_74832[3];
  assign array_update_74840[4] = literal_74722 == 32'h0000_0004 ? add_74838 : array_index_74832[4];
  assign array_update_74840[5] = literal_74722 == 32'h0000_0005 ? add_74838 : array_index_74832[5];
  assign array_update_74840[6] = literal_74722 == 32'h0000_0006 ? add_74838 : array_index_74832[6];
  assign array_update_74840[7] = literal_74722 == 32'h0000_0007 ? add_74838 : array_index_74832[7];
  assign array_update_74840[8] = literal_74722 == 32'h0000_0008 ? add_74838 : array_index_74832[8];
  assign array_update_74840[9] = literal_74722 == 32'h0000_0009 ? add_74838 : array_index_74832[9];
  assign add_74841 = add_74828 + 32'h0000_0001;
  assign array_update_74842[0] = add_74719 == 32'h0000_0000 ? array_update_74840 : array_update_74829[0];
  assign array_update_74842[1] = add_74719 == 32'h0000_0001 ? array_update_74840 : array_update_74829[1];
  assign array_update_74842[2] = add_74719 == 32'h0000_0002 ? array_update_74840 : array_update_74829[2];
  assign array_update_74842[3] = add_74719 == 32'h0000_0003 ? array_update_74840 : array_update_74829[3];
  assign array_update_74842[4] = add_74719 == 32'h0000_0004 ? array_update_74840 : array_update_74829[4];
  assign array_update_74842[5] = add_74719 == 32'h0000_0005 ? array_update_74840 : array_update_74829[5];
  assign array_update_74842[6] = add_74719 == 32'h0000_0006 ? array_update_74840 : array_update_74829[6];
  assign array_update_74842[7] = add_74719 == 32'h0000_0007 ? array_update_74840 : array_update_74829[7];
  assign array_update_74842[8] = add_74719 == 32'h0000_0008 ? array_update_74840 : array_update_74829[8];
  assign array_update_74842[9] = add_74719 == 32'h0000_0009 ? array_update_74840 : array_update_74829[9];
  assign array_index_74844 = array_update_72021[add_74841 > 32'h0000_0009 ? 4'h9 : add_74841[3:0]];
  assign array_index_74845 = array_update_74842[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_74849 = smul32b_32b_x_32b(array_index_74726[add_74841 > 32'h0000_0009 ? 4'h9 : add_74841[3:0]], array_index_74844[literal_74722 > 32'h0000_0009 ? 4'h9 : literal_74722[3:0]]);
  assign add_74851 = array_index_74845[literal_74722 > 32'h0000_0009 ? 4'h9 : literal_74722[3:0]] + smul_74849;
  assign array_update_74852[0] = literal_74722 == 32'h0000_0000 ? add_74851 : array_index_74845[0];
  assign array_update_74852[1] = literal_74722 == 32'h0000_0001 ? add_74851 : array_index_74845[1];
  assign array_update_74852[2] = literal_74722 == 32'h0000_0002 ? add_74851 : array_index_74845[2];
  assign array_update_74852[3] = literal_74722 == 32'h0000_0003 ? add_74851 : array_index_74845[3];
  assign array_update_74852[4] = literal_74722 == 32'h0000_0004 ? add_74851 : array_index_74845[4];
  assign array_update_74852[5] = literal_74722 == 32'h0000_0005 ? add_74851 : array_index_74845[5];
  assign array_update_74852[6] = literal_74722 == 32'h0000_0006 ? add_74851 : array_index_74845[6];
  assign array_update_74852[7] = literal_74722 == 32'h0000_0007 ? add_74851 : array_index_74845[7];
  assign array_update_74852[8] = literal_74722 == 32'h0000_0008 ? add_74851 : array_index_74845[8];
  assign array_update_74852[9] = literal_74722 == 32'h0000_0009 ? add_74851 : array_index_74845[9];
  assign array_update_74853[0] = add_74719 == 32'h0000_0000 ? array_update_74852 : array_update_74842[0];
  assign array_update_74853[1] = add_74719 == 32'h0000_0001 ? array_update_74852 : array_update_74842[1];
  assign array_update_74853[2] = add_74719 == 32'h0000_0002 ? array_update_74852 : array_update_74842[2];
  assign array_update_74853[3] = add_74719 == 32'h0000_0003 ? array_update_74852 : array_update_74842[3];
  assign array_update_74853[4] = add_74719 == 32'h0000_0004 ? array_update_74852 : array_update_74842[4];
  assign array_update_74853[5] = add_74719 == 32'h0000_0005 ? array_update_74852 : array_update_74842[5];
  assign array_update_74853[6] = add_74719 == 32'h0000_0006 ? array_update_74852 : array_update_74842[6];
  assign array_update_74853[7] = add_74719 == 32'h0000_0007 ? array_update_74852 : array_update_74842[7];
  assign array_update_74853[8] = add_74719 == 32'h0000_0008 ? array_update_74852 : array_update_74842[8];
  assign array_update_74853[9] = add_74719 == 32'h0000_0009 ? array_update_74852 : array_update_74842[9];
  assign array_index_74855 = array_update_74853[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign add_74857 = literal_74722 + 32'h0000_0001;
  assign array_update_74858[0] = add_74857 == 32'h0000_0000 ? 32'h0000_0000 : array_index_74855[0];
  assign array_update_74858[1] = add_74857 == 32'h0000_0001 ? 32'h0000_0000 : array_index_74855[1];
  assign array_update_74858[2] = add_74857 == 32'h0000_0002 ? 32'h0000_0000 : array_index_74855[2];
  assign array_update_74858[3] = add_74857 == 32'h0000_0003 ? 32'h0000_0000 : array_index_74855[3];
  assign array_update_74858[4] = add_74857 == 32'h0000_0004 ? 32'h0000_0000 : array_index_74855[4];
  assign array_update_74858[5] = add_74857 == 32'h0000_0005 ? 32'h0000_0000 : array_index_74855[5];
  assign array_update_74858[6] = add_74857 == 32'h0000_0006 ? 32'h0000_0000 : array_index_74855[6];
  assign array_update_74858[7] = add_74857 == 32'h0000_0007 ? 32'h0000_0000 : array_index_74855[7];
  assign array_update_74858[8] = add_74857 == 32'h0000_0008 ? 32'h0000_0000 : array_index_74855[8];
  assign array_update_74858[9] = add_74857 == 32'h0000_0009 ? 32'h0000_0000 : array_index_74855[9];
  assign literal_74859 = 32'h0000_0000;
  assign array_update_74860[0] = add_74719 == 32'h0000_0000 ? array_update_74858 : array_update_74853[0];
  assign array_update_74860[1] = add_74719 == 32'h0000_0001 ? array_update_74858 : array_update_74853[1];
  assign array_update_74860[2] = add_74719 == 32'h0000_0002 ? array_update_74858 : array_update_74853[2];
  assign array_update_74860[3] = add_74719 == 32'h0000_0003 ? array_update_74858 : array_update_74853[3];
  assign array_update_74860[4] = add_74719 == 32'h0000_0004 ? array_update_74858 : array_update_74853[4];
  assign array_update_74860[5] = add_74719 == 32'h0000_0005 ? array_update_74858 : array_update_74853[5];
  assign array_update_74860[6] = add_74719 == 32'h0000_0006 ? array_update_74858 : array_update_74853[6];
  assign array_update_74860[7] = add_74719 == 32'h0000_0007 ? array_update_74858 : array_update_74853[7];
  assign array_update_74860[8] = add_74719 == 32'h0000_0008 ? array_update_74858 : array_update_74853[8];
  assign array_update_74860[9] = add_74719 == 32'h0000_0009 ? array_update_74858 : array_update_74853[9];
  assign array_index_74862 = array_update_72021[literal_74859 > 32'h0000_0009 ? 4'h9 : literal_74859[3:0]];
  assign array_index_74863 = array_update_74860[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_74867 = smul32b_32b_x_32b(array_index_74726[literal_74859 > 32'h0000_0009 ? 4'h9 : literal_74859[3:0]], array_index_74862[add_74857 > 32'h0000_0009 ? 4'h9 : add_74857[3:0]]);
  assign add_74869 = array_index_74863[add_74857 > 32'h0000_0009 ? 4'h9 : add_74857[3:0]] + smul_74867;
  assign array_update_74871[0] = add_74857 == 32'h0000_0000 ? add_74869 : array_index_74863[0];
  assign array_update_74871[1] = add_74857 == 32'h0000_0001 ? add_74869 : array_index_74863[1];
  assign array_update_74871[2] = add_74857 == 32'h0000_0002 ? add_74869 : array_index_74863[2];
  assign array_update_74871[3] = add_74857 == 32'h0000_0003 ? add_74869 : array_index_74863[3];
  assign array_update_74871[4] = add_74857 == 32'h0000_0004 ? add_74869 : array_index_74863[4];
  assign array_update_74871[5] = add_74857 == 32'h0000_0005 ? add_74869 : array_index_74863[5];
  assign array_update_74871[6] = add_74857 == 32'h0000_0006 ? add_74869 : array_index_74863[6];
  assign array_update_74871[7] = add_74857 == 32'h0000_0007 ? add_74869 : array_index_74863[7];
  assign array_update_74871[8] = add_74857 == 32'h0000_0008 ? add_74869 : array_index_74863[8];
  assign array_update_74871[9] = add_74857 == 32'h0000_0009 ? add_74869 : array_index_74863[9];
  assign add_74872 = literal_74859 + 32'h0000_0001;
  assign array_update_74873[0] = add_74719 == 32'h0000_0000 ? array_update_74871 : array_update_74860[0];
  assign array_update_74873[1] = add_74719 == 32'h0000_0001 ? array_update_74871 : array_update_74860[1];
  assign array_update_74873[2] = add_74719 == 32'h0000_0002 ? array_update_74871 : array_update_74860[2];
  assign array_update_74873[3] = add_74719 == 32'h0000_0003 ? array_update_74871 : array_update_74860[3];
  assign array_update_74873[4] = add_74719 == 32'h0000_0004 ? array_update_74871 : array_update_74860[4];
  assign array_update_74873[5] = add_74719 == 32'h0000_0005 ? array_update_74871 : array_update_74860[5];
  assign array_update_74873[6] = add_74719 == 32'h0000_0006 ? array_update_74871 : array_update_74860[6];
  assign array_update_74873[7] = add_74719 == 32'h0000_0007 ? array_update_74871 : array_update_74860[7];
  assign array_update_74873[8] = add_74719 == 32'h0000_0008 ? array_update_74871 : array_update_74860[8];
  assign array_update_74873[9] = add_74719 == 32'h0000_0009 ? array_update_74871 : array_update_74860[9];
  assign array_index_74875 = array_update_72021[add_74872 > 32'h0000_0009 ? 4'h9 : add_74872[3:0]];
  assign array_index_74876 = array_update_74873[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_74880 = smul32b_32b_x_32b(array_index_74726[add_74872 > 32'h0000_0009 ? 4'h9 : add_74872[3:0]], array_index_74875[add_74857 > 32'h0000_0009 ? 4'h9 : add_74857[3:0]]);
  assign add_74882 = array_index_74876[add_74857 > 32'h0000_0009 ? 4'h9 : add_74857[3:0]] + smul_74880;
  assign array_update_74884[0] = add_74857 == 32'h0000_0000 ? add_74882 : array_index_74876[0];
  assign array_update_74884[1] = add_74857 == 32'h0000_0001 ? add_74882 : array_index_74876[1];
  assign array_update_74884[2] = add_74857 == 32'h0000_0002 ? add_74882 : array_index_74876[2];
  assign array_update_74884[3] = add_74857 == 32'h0000_0003 ? add_74882 : array_index_74876[3];
  assign array_update_74884[4] = add_74857 == 32'h0000_0004 ? add_74882 : array_index_74876[4];
  assign array_update_74884[5] = add_74857 == 32'h0000_0005 ? add_74882 : array_index_74876[5];
  assign array_update_74884[6] = add_74857 == 32'h0000_0006 ? add_74882 : array_index_74876[6];
  assign array_update_74884[7] = add_74857 == 32'h0000_0007 ? add_74882 : array_index_74876[7];
  assign array_update_74884[8] = add_74857 == 32'h0000_0008 ? add_74882 : array_index_74876[8];
  assign array_update_74884[9] = add_74857 == 32'h0000_0009 ? add_74882 : array_index_74876[9];
  assign add_74885 = add_74872 + 32'h0000_0001;
  assign array_update_74886[0] = add_74719 == 32'h0000_0000 ? array_update_74884 : array_update_74873[0];
  assign array_update_74886[1] = add_74719 == 32'h0000_0001 ? array_update_74884 : array_update_74873[1];
  assign array_update_74886[2] = add_74719 == 32'h0000_0002 ? array_update_74884 : array_update_74873[2];
  assign array_update_74886[3] = add_74719 == 32'h0000_0003 ? array_update_74884 : array_update_74873[3];
  assign array_update_74886[4] = add_74719 == 32'h0000_0004 ? array_update_74884 : array_update_74873[4];
  assign array_update_74886[5] = add_74719 == 32'h0000_0005 ? array_update_74884 : array_update_74873[5];
  assign array_update_74886[6] = add_74719 == 32'h0000_0006 ? array_update_74884 : array_update_74873[6];
  assign array_update_74886[7] = add_74719 == 32'h0000_0007 ? array_update_74884 : array_update_74873[7];
  assign array_update_74886[8] = add_74719 == 32'h0000_0008 ? array_update_74884 : array_update_74873[8];
  assign array_update_74886[9] = add_74719 == 32'h0000_0009 ? array_update_74884 : array_update_74873[9];
  assign array_index_74888 = array_update_72021[add_74885 > 32'h0000_0009 ? 4'h9 : add_74885[3:0]];
  assign array_index_74889 = array_update_74886[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_74893 = smul32b_32b_x_32b(array_index_74726[add_74885 > 32'h0000_0009 ? 4'h9 : add_74885[3:0]], array_index_74888[add_74857 > 32'h0000_0009 ? 4'h9 : add_74857[3:0]]);
  assign add_74895 = array_index_74889[add_74857 > 32'h0000_0009 ? 4'h9 : add_74857[3:0]] + smul_74893;
  assign array_update_74897[0] = add_74857 == 32'h0000_0000 ? add_74895 : array_index_74889[0];
  assign array_update_74897[1] = add_74857 == 32'h0000_0001 ? add_74895 : array_index_74889[1];
  assign array_update_74897[2] = add_74857 == 32'h0000_0002 ? add_74895 : array_index_74889[2];
  assign array_update_74897[3] = add_74857 == 32'h0000_0003 ? add_74895 : array_index_74889[3];
  assign array_update_74897[4] = add_74857 == 32'h0000_0004 ? add_74895 : array_index_74889[4];
  assign array_update_74897[5] = add_74857 == 32'h0000_0005 ? add_74895 : array_index_74889[5];
  assign array_update_74897[6] = add_74857 == 32'h0000_0006 ? add_74895 : array_index_74889[6];
  assign array_update_74897[7] = add_74857 == 32'h0000_0007 ? add_74895 : array_index_74889[7];
  assign array_update_74897[8] = add_74857 == 32'h0000_0008 ? add_74895 : array_index_74889[8];
  assign array_update_74897[9] = add_74857 == 32'h0000_0009 ? add_74895 : array_index_74889[9];
  assign add_74898 = add_74885 + 32'h0000_0001;
  assign array_update_74899[0] = add_74719 == 32'h0000_0000 ? array_update_74897 : array_update_74886[0];
  assign array_update_74899[1] = add_74719 == 32'h0000_0001 ? array_update_74897 : array_update_74886[1];
  assign array_update_74899[2] = add_74719 == 32'h0000_0002 ? array_update_74897 : array_update_74886[2];
  assign array_update_74899[3] = add_74719 == 32'h0000_0003 ? array_update_74897 : array_update_74886[3];
  assign array_update_74899[4] = add_74719 == 32'h0000_0004 ? array_update_74897 : array_update_74886[4];
  assign array_update_74899[5] = add_74719 == 32'h0000_0005 ? array_update_74897 : array_update_74886[5];
  assign array_update_74899[6] = add_74719 == 32'h0000_0006 ? array_update_74897 : array_update_74886[6];
  assign array_update_74899[7] = add_74719 == 32'h0000_0007 ? array_update_74897 : array_update_74886[7];
  assign array_update_74899[8] = add_74719 == 32'h0000_0008 ? array_update_74897 : array_update_74886[8];
  assign array_update_74899[9] = add_74719 == 32'h0000_0009 ? array_update_74897 : array_update_74886[9];
  assign array_index_74901 = array_update_72021[add_74898 > 32'h0000_0009 ? 4'h9 : add_74898[3:0]];
  assign array_index_74902 = array_update_74899[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_74906 = smul32b_32b_x_32b(array_index_74726[add_74898 > 32'h0000_0009 ? 4'h9 : add_74898[3:0]], array_index_74901[add_74857 > 32'h0000_0009 ? 4'h9 : add_74857[3:0]]);
  assign add_74908 = array_index_74902[add_74857 > 32'h0000_0009 ? 4'h9 : add_74857[3:0]] + smul_74906;
  assign array_update_74910[0] = add_74857 == 32'h0000_0000 ? add_74908 : array_index_74902[0];
  assign array_update_74910[1] = add_74857 == 32'h0000_0001 ? add_74908 : array_index_74902[1];
  assign array_update_74910[2] = add_74857 == 32'h0000_0002 ? add_74908 : array_index_74902[2];
  assign array_update_74910[3] = add_74857 == 32'h0000_0003 ? add_74908 : array_index_74902[3];
  assign array_update_74910[4] = add_74857 == 32'h0000_0004 ? add_74908 : array_index_74902[4];
  assign array_update_74910[5] = add_74857 == 32'h0000_0005 ? add_74908 : array_index_74902[5];
  assign array_update_74910[6] = add_74857 == 32'h0000_0006 ? add_74908 : array_index_74902[6];
  assign array_update_74910[7] = add_74857 == 32'h0000_0007 ? add_74908 : array_index_74902[7];
  assign array_update_74910[8] = add_74857 == 32'h0000_0008 ? add_74908 : array_index_74902[8];
  assign array_update_74910[9] = add_74857 == 32'h0000_0009 ? add_74908 : array_index_74902[9];
  assign add_74911 = add_74898 + 32'h0000_0001;
  assign array_update_74912[0] = add_74719 == 32'h0000_0000 ? array_update_74910 : array_update_74899[0];
  assign array_update_74912[1] = add_74719 == 32'h0000_0001 ? array_update_74910 : array_update_74899[1];
  assign array_update_74912[2] = add_74719 == 32'h0000_0002 ? array_update_74910 : array_update_74899[2];
  assign array_update_74912[3] = add_74719 == 32'h0000_0003 ? array_update_74910 : array_update_74899[3];
  assign array_update_74912[4] = add_74719 == 32'h0000_0004 ? array_update_74910 : array_update_74899[4];
  assign array_update_74912[5] = add_74719 == 32'h0000_0005 ? array_update_74910 : array_update_74899[5];
  assign array_update_74912[6] = add_74719 == 32'h0000_0006 ? array_update_74910 : array_update_74899[6];
  assign array_update_74912[7] = add_74719 == 32'h0000_0007 ? array_update_74910 : array_update_74899[7];
  assign array_update_74912[8] = add_74719 == 32'h0000_0008 ? array_update_74910 : array_update_74899[8];
  assign array_update_74912[9] = add_74719 == 32'h0000_0009 ? array_update_74910 : array_update_74899[9];
  assign array_index_74914 = array_update_72021[add_74911 > 32'h0000_0009 ? 4'h9 : add_74911[3:0]];
  assign array_index_74915 = array_update_74912[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_74919 = smul32b_32b_x_32b(array_index_74726[add_74911 > 32'h0000_0009 ? 4'h9 : add_74911[3:0]], array_index_74914[add_74857 > 32'h0000_0009 ? 4'h9 : add_74857[3:0]]);
  assign add_74921 = array_index_74915[add_74857 > 32'h0000_0009 ? 4'h9 : add_74857[3:0]] + smul_74919;
  assign array_update_74923[0] = add_74857 == 32'h0000_0000 ? add_74921 : array_index_74915[0];
  assign array_update_74923[1] = add_74857 == 32'h0000_0001 ? add_74921 : array_index_74915[1];
  assign array_update_74923[2] = add_74857 == 32'h0000_0002 ? add_74921 : array_index_74915[2];
  assign array_update_74923[3] = add_74857 == 32'h0000_0003 ? add_74921 : array_index_74915[3];
  assign array_update_74923[4] = add_74857 == 32'h0000_0004 ? add_74921 : array_index_74915[4];
  assign array_update_74923[5] = add_74857 == 32'h0000_0005 ? add_74921 : array_index_74915[5];
  assign array_update_74923[6] = add_74857 == 32'h0000_0006 ? add_74921 : array_index_74915[6];
  assign array_update_74923[7] = add_74857 == 32'h0000_0007 ? add_74921 : array_index_74915[7];
  assign array_update_74923[8] = add_74857 == 32'h0000_0008 ? add_74921 : array_index_74915[8];
  assign array_update_74923[9] = add_74857 == 32'h0000_0009 ? add_74921 : array_index_74915[9];
  assign add_74924 = add_74911 + 32'h0000_0001;
  assign array_update_74925[0] = add_74719 == 32'h0000_0000 ? array_update_74923 : array_update_74912[0];
  assign array_update_74925[1] = add_74719 == 32'h0000_0001 ? array_update_74923 : array_update_74912[1];
  assign array_update_74925[2] = add_74719 == 32'h0000_0002 ? array_update_74923 : array_update_74912[2];
  assign array_update_74925[3] = add_74719 == 32'h0000_0003 ? array_update_74923 : array_update_74912[3];
  assign array_update_74925[4] = add_74719 == 32'h0000_0004 ? array_update_74923 : array_update_74912[4];
  assign array_update_74925[5] = add_74719 == 32'h0000_0005 ? array_update_74923 : array_update_74912[5];
  assign array_update_74925[6] = add_74719 == 32'h0000_0006 ? array_update_74923 : array_update_74912[6];
  assign array_update_74925[7] = add_74719 == 32'h0000_0007 ? array_update_74923 : array_update_74912[7];
  assign array_update_74925[8] = add_74719 == 32'h0000_0008 ? array_update_74923 : array_update_74912[8];
  assign array_update_74925[9] = add_74719 == 32'h0000_0009 ? array_update_74923 : array_update_74912[9];
  assign array_index_74927 = array_update_72021[add_74924 > 32'h0000_0009 ? 4'h9 : add_74924[3:0]];
  assign array_index_74928 = array_update_74925[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_74932 = smul32b_32b_x_32b(array_index_74726[add_74924 > 32'h0000_0009 ? 4'h9 : add_74924[3:0]], array_index_74927[add_74857 > 32'h0000_0009 ? 4'h9 : add_74857[3:0]]);
  assign add_74934 = array_index_74928[add_74857 > 32'h0000_0009 ? 4'h9 : add_74857[3:0]] + smul_74932;
  assign array_update_74936[0] = add_74857 == 32'h0000_0000 ? add_74934 : array_index_74928[0];
  assign array_update_74936[1] = add_74857 == 32'h0000_0001 ? add_74934 : array_index_74928[1];
  assign array_update_74936[2] = add_74857 == 32'h0000_0002 ? add_74934 : array_index_74928[2];
  assign array_update_74936[3] = add_74857 == 32'h0000_0003 ? add_74934 : array_index_74928[3];
  assign array_update_74936[4] = add_74857 == 32'h0000_0004 ? add_74934 : array_index_74928[4];
  assign array_update_74936[5] = add_74857 == 32'h0000_0005 ? add_74934 : array_index_74928[5];
  assign array_update_74936[6] = add_74857 == 32'h0000_0006 ? add_74934 : array_index_74928[6];
  assign array_update_74936[7] = add_74857 == 32'h0000_0007 ? add_74934 : array_index_74928[7];
  assign array_update_74936[8] = add_74857 == 32'h0000_0008 ? add_74934 : array_index_74928[8];
  assign array_update_74936[9] = add_74857 == 32'h0000_0009 ? add_74934 : array_index_74928[9];
  assign add_74937 = add_74924 + 32'h0000_0001;
  assign array_update_74938[0] = add_74719 == 32'h0000_0000 ? array_update_74936 : array_update_74925[0];
  assign array_update_74938[1] = add_74719 == 32'h0000_0001 ? array_update_74936 : array_update_74925[1];
  assign array_update_74938[2] = add_74719 == 32'h0000_0002 ? array_update_74936 : array_update_74925[2];
  assign array_update_74938[3] = add_74719 == 32'h0000_0003 ? array_update_74936 : array_update_74925[3];
  assign array_update_74938[4] = add_74719 == 32'h0000_0004 ? array_update_74936 : array_update_74925[4];
  assign array_update_74938[5] = add_74719 == 32'h0000_0005 ? array_update_74936 : array_update_74925[5];
  assign array_update_74938[6] = add_74719 == 32'h0000_0006 ? array_update_74936 : array_update_74925[6];
  assign array_update_74938[7] = add_74719 == 32'h0000_0007 ? array_update_74936 : array_update_74925[7];
  assign array_update_74938[8] = add_74719 == 32'h0000_0008 ? array_update_74936 : array_update_74925[8];
  assign array_update_74938[9] = add_74719 == 32'h0000_0009 ? array_update_74936 : array_update_74925[9];
  assign array_index_74940 = array_update_72021[add_74937 > 32'h0000_0009 ? 4'h9 : add_74937[3:0]];
  assign array_index_74941 = array_update_74938[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_74945 = smul32b_32b_x_32b(array_index_74726[add_74937 > 32'h0000_0009 ? 4'h9 : add_74937[3:0]], array_index_74940[add_74857 > 32'h0000_0009 ? 4'h9 : add_74857[3:0]]);
  assign add_74947 = array_index_74941[add_74857 > 32'h0000_0009 ? 4'h9 : add_74857[3:0]] + smul_74945;
  assign array_update_74949[0] = add_74857 == 32'h0000_0000 ? add_74947 : array_index_74941[0];
  assign array_update_74949[1] = add_74857 == 32'h0000_0001 ? add_74947 : array_index_74941[1];
  assign array_update_74949[2] = add_74857 == 32'h0000_0002 ? add_74947 : array_index_74941[2];
  assign array_update_74949[3] = add_74857 == 32'h0000_0003 ? add_74947 : array_index_74941[3];
  assign array_update_74949[4] = add_74857 == 32'h0000_0004 ? add_74947 : array_index_74941[4];
  assign array_update_74949[5] = add_74857 == 32'h0000_0005 ? add_74947 : array_index_74941[5];
  assign array_update_74949[6] = add_74857 == 32'h0000_0006 ? add_74947 : array_index_74941[6];
  assign array_update_74949[7] = add_74857 == 32'h0000_0007 ? add_74947 : array_index_74941[7];
  assign array_update_74949[8] = add_74857 == 32'h0000_0008 ? add_74947 : array_index_74941[8];
  assign array_update_74949[9] = add_74857 == 32'h0000_0009 ? add_74947 : array_index_74941[9];
  assign add_74950 = add_74937 + 32'h0000_0001;
  assign array_update_74951[0] = add_74719 == 32'h0000_0000 ? array_update_74949 : array_update_74938[0];
  assign array_update_74951[1] = add_74719 == 32'h0000_0001 ? array_update_74949 : array_update_74938[1];
  assign array_update_74951[2] = add_74719 == 32'h0000_0002 ? array_update_74949 : array_update_74938[2];
  assign array_update_74951[3] = add_74719 == 32'h0000_0003 ? array_update_74949 : array_update_74938[3];
  assign array_update_74951[4] = add_74719 == 32'h0000_0004 ? array_update_74949 : array_update_74938[4];
  assign array_update_74951[5] = add_74719 == 32'h0000_0005 ? array_update_74949 : array_update_74938[5];
  assign array_update_74951[6] = add_74719 == 32'h0000_0006 ? array_update_74949 : array_update_74938[6];
  assign array_update_74951[7] = add_74719 == 32'h0000_0007 ? array_update_74949 : array_update_74938[7];
  assign array_update_74951[8] = add_74719 == 32'h0000_0008 ? array_update_74949 : array_update_74938[8];
  assign array_update_74951[9] = add_74719 == 32'h0000_0009 ? array_update_74949 : array_update_74938[9];
  assign array_index_74953 = array_update_72021[add_74950 > 32'h0000_0009 ? 4'h9 : add_74950[3:0]];
  assign array_index_74954 = array_update_74951[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_74958 = smul32b_32b_x_32b(array_index_74726[add_74950 > 32'h0000_0009 ? 4'h9 : add_74950[3:0]], array_index_74953[add_74857 > 32'h0000_0009 ? 4'h9 : add_74857[3:0]]);
  assign add_74960 = array_index_74954[add_74857 > 32'h0000_0009 ? 4'h9 : add_74857[3:0]] + smul_74958;
  assign array_update_74962[0] = add_74857 == 32'h0000_0000 ? add_74960 : array_index_74954[0];
  assign array_update_74962[1] = add_74857 == 32'h0000_0001 ? add_74960 : array_index_74954[1];
  assign array_update_74962[2] = add_74857 == 32'h0000_0002 ? add_74960 : array_index_74954[2];
  assign array_update_74962[3] = add_74857 == 32'h0000_0003 ? add_74960 : array_index_74954[3];
  assign array_update_74962[4] = add_74857 == 32'h0000_0004 ? add_74960 : array_index_74954[4];
  assign array_update_74962[5] = add_74857 == 32'h0000_0005 ? add_74960 : array_index_74954[5];
  assign array_update_74962[6] = add_74857 == 32'h0000_0006 ? add_74960 : array_index_74954[6];
  assign array_update_74962[7] = add_74857 == 32'h0000_0007 ? add_74960 : array_index_74954[7];
  assign array_update_74962[8] = add_74857 == 32'h0000_0008 ? add_74960 : array_index_74954[8];
  assign array_update_74962[9] = add_74857 == 32'h0000_0009 ? add_74960 : array_index_74954[9];
  assign add_74963 = add_74950 + 32'h0000_0001;
  assign array_update_74964[0] = add_74719 == 32'h0000_0000 ? array_update_74962 : array_update_74951[0];
  assign array_update_74964[1] = add_74719 == 32'h0000_0001 ? array_update_74962 : array_update_74951[1];
  assign array_update_74964[2] = add_74719 == 32'h0000_0002 ? array_update_74962 : array_update_74951[2];
  assign array_update_74964[3] = add_74719 == 32'h0000_0003 ? array_update_74962 : array_update_74951[3];
  assign array_update_74964[4] = add_74719 == 32'h0000_0004 ? array_update_74962 : array_update_74951[4];
  assign array_update_74964[5] = add_74719 == 32'h0000_0005 ? array_update_74962 : array_update_74951[5];
  assign array_update_74964[6] = add_74719 == 32'h0000_0006 ? array_update_74962 : array_update_74951[6];
  assign array_update_74964[7] = add_74719 == 32'h0000_0007 ? array_update_74962 : array_update_74951[7];
  assign array_update_74964[8] = add_74719 == 32'h0000_0008 ? array_update_74962 : array_update_74951[8];
  assign array_update_74964[9] = add_74719 == 32'h0000_0009 ? array_update_74962 : array_update_74951[9];
  assign array_index_74966 = array_update_72021[add_74963 > 32'h0000_0009 ? 4'h9 : add_74963[3:0]];
  assign array_index_74967 = array_update_74964[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_74971 = smul32b_32b_x_32b(array_index_74726[add_74963 > 32'h0000_0009 ? 4'h9 : add_74963[3:0]], array_index_74966[add_74857 > 32'h0000_0009 ? 4'h9 : add_74857[3:0]]);
  assign add_74973 = array_index_74967[add_74857 > 32'h0000_0009 ? 4'h9 : add_74857[3:0]] + smul_74971;
  assign array_update_74975[0] = add_74857 == 32'h0000_0000 ? add_74973 : array_index_74967[0];
  assign array_update_74975[1] = add_74857 == 32'h0000_0001 ? add_74973 : array_index_74967[1];
  assign array_update_74975[2] = add_74857 == 32'h0000_0002 ? add_74973 : array_index_74967[2];
  assign array_update_74975[3] = add_74857 == 32'h0000_0003 ? add_74973 : array_index_74967[3];
  assign array_update_74975[4] = add_74857 == 32'h0000_0004 ? add_74973 : array_index_74967[4];
  assign array_update_74975[5] = add_74857 == 32'h0000_0005 ? add_74973 : array_index_74967[5];
  assign array_update_74975[6] = add_74857 == 32'h0000_0006 ? add_74973 : array_index_74967[6];
  assign array_update_74975[7] = add_74857 == 32'h0000_0007 ? add_74973 : array_index_74967[7];
  assign array_update_74975[8] = add_74857 == 32'h0000_0008 ? add_74973 : array_index_74967[8];
  assign array_update_74975[9] = add_74857 == 32'h0000_0009 ? add_74973 : array_index_74967[9];
  assign add_74976 = add_74963 + 32'h0000_0001;
  assign array_update_74977[0] = add_74719 == 32'h0000_0000 ? array_update_74975 : array_update_74964[0];
  assign array_update_74977[1] = add_74719 == 32'h0000_0001 ? array_update_74975 : array_update_74964[1];
  assign array_update_74977[2] = add_74719 == 32'h0000_0002 ? array_update_74975 : array_update_74964[2];
  assign array_update_74977[3] = add_74719 == 32'h0000_0003 ? array_update_74975 : array_update_74964[3];
  assign array_update_74977[4] = add_74719 == 32'h0000_0004 ? array_update_74975 : array_update_74964[4];
  assign array_update_74977[5] = add_74719 == 32'h0000_0005 ? array_update_74975 : array_update_74964[5];
  assign array_update_74977[6] = add_74719 == 32'h0000_0006 ? array_update_74975 : array_update_74964[6];
  assign array_update_74977[7] = add_74719 == 32'h0000_0007 ? array_update_74975 : array_update_74964[7];
  assign array_update_74977[8] = add_74719 == 32'h0000_0008 ? array_update_74975 : array_update_74964[8];
  assign array_update_74977[9] = add_74719 == 32'h0000_0009 ? array_update_74975 : array_update_74964[9];
  assign array_index_74979 = array_update_72021[add_74976 > 32'h0000_0009 ? 4'h9 : add_74976[3:0]];
  assign array_index_74980 = array_update_74977[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_74984 = smul32b_32b_x_32b(array_index_74726[add_74976 > 32'h0000_0009 ? 4'h9 : add_74976[3:0]], array_index_74979[add_74857 > 32'h0000_0009 ? 4'h9 : add_74857[3:0]]);
  assign add_74986 = array_index_74980[add_74857 > 32'h0000_0009 ? 4'h9 : add_74857[3:0]] + smul_74984;
  assign array_update_74987[0] = add_74857 == 32'h0000_0000 ? add_74986 : array_index_74980[0];
  assign array_update_74987[1] = add_74857 == 32'h0000_0001 ? add_74986 : array_index_74980[1];
  assign array_update_74987[2] = add_74857 == 32'h0000_0002 ? add_74986 : array_index_74980[2];
  assign array_update_74987[3] = add_74857 == 32'h0000_0003 ? add_74986 : array_index_74980[3];
  assign array_update_74987[4] = add_74857 == 32'h0000_0004 ? add_74986 : array_index_74980[4];
  assign array_update_74987[5] = add_74857 == 32'h0000_0005 ? add_74986 : array_index_74980[5];
  assign array_update_74987[6] = add_74857 == 32'h0000_0006 ? add_74986 : array_index_74980[6];
  assign array_update_74987[7] = add_74857 == 32'h0000_0007 ? add_74986 : array_index_74980[7];
  assign array_update_74987[8] = add_74857 == 32'h0000_0008 ? add_74986 : array_index_74980[8];
  assign array_update_74987[9] = add_74857 == 32'h0000_0009 ? add_74986 : array_index_74980[9];
  assign array_update_74988[0] = add_74719 == 32'h0000_0000 ? array_update_74987 : array_update_74977[0];
  assign array_update_74988[1] = add_74719 == 32'h0000_0001 ? array_update_74987 : array_update_74977[1];
  assign array_update_74988[2] = add_74719 == 32'h0000_0002 ? array_update_74987 : array_update_74977[2];
  assign array_update_74988[3] = add_74719 == 32'h0000_0003 ? array_update_74987 : array_update_74977[3];
  assign array_update_74988[4] = add_74719 == 32'h0000_0004 ? array_update_74987 : array_update_74977[4];
  assign array_update_74988[5] = add_74719 == 32'h0000_0005 ? array_update_74987 : array_update_74977[5];
  assign array_update_74988[6] = add_74719 == 32'h0000_0006 ? array_update_74987 : array_update_74977[6];
  assign array_update_74988[7] = add_74719 == 32'h0000_0007 ? array_update_74987 : array_update_74977[7];
  assign array_update_74988[8] = add_74719 == 32'h0000_0008 ? array_update_74987 : array_update_74977[8];
  assign array_update_74988[9] = add_74719 == 32'h0000_0009 ? array_update_74987 : array_update_74977[9];
  assign array_index_74990 = array_update_74988[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign add_74992 = add_74857 + 32'h0000_0001;
  assign array_update_74993[0] = add_74992 == 32'h0000_0000 ? 32'h0000_0000 : array_index_74990[0];
  assign array_update_74993[1] = add_74992 == 32'h0000_0001 ? 32'h0000_0000 : array_index_74990[1];
  assign array_update_74993[2] = add_74992 == 32'h0000_0002 ? 32'h0000_0000 : array_index_74990[2];
  assign array_update_74993[3] = add_74992 == 32'h0000_0003 ? 32'h0000_0000 : array_index_74990[3];
  assign array_update_74993[4] = add_74992 == 32'h0000_0004 ? 32'h0000_0000 : array_index_74990[4];
  assign array_update_74993[5] = add_74992 == 32'h0000_0005 ? 32'h0000_0000 : array_index_74990[5];
  assign array_update_74993[6] = add_74992 == 32'h0000_0006 ? 32'h0000_0000 : array_index_74990[6];
  assign array_update_74993[7] = add_74992 == 32'h0000_0007 ? 32'h0000_0000 : array_index_74990[7];
  assign array_update_74993[8] = add_74992 == 32'h0000_0008 ? 32'h0000_0000 : array_index_74990[8];
  assign array_update_74993[9] = add_74992 == 32'h0000_0009 ? 32'h0000_0000 : array_index_74990[9];
  assign literal_74994 = 32'h0000_0000;
  assign array_update_74995[0] = add_74719 == 32'h0000_0000 ? array_update_74993 : array_update_74988[0];
  assign array_update_74995[1] = add_74719 == 32'h0000_0001 ? array_update_74993 : array_update_74988[1];
  assign array_update_74995[2] = add_74719 == 32'h0000_0002 ? array_update_74993 : array_update_74988[2];
  assign array_update_74995[3] = add_74719 == 32'h0000_0003 ? array_update_74993 : array_update_74988[3];
  assign array_update_74995[4] = add_74719 == 32'h0000_0004 ? array_update_74993 : array_update_74988[4];
  assign array_update_74995[5] = add_74719 == 32'h0000_0005 ? array_update_74993 : array_update_74988[5];
  assign array_update_74995[6] = add_74719 == 32'h0000_0006 ? array_update_74993 : array_update_74988[6];
  assign array_update_74995[7] = add_74719 == 32'h0000_0007 ? array_update_74993 : array_update_74988[7];
  assign array_update_74995[8] = add_74719 == 32'h0000_0008 ? array_update_74993 : array_update_74988[8];
  assign array_update_74995[9] = add_74719 == 32'h0000_0009 ? array_update_74993 : array_update_74988[9];
  assign array_index_74997 = array_update_72021[literal_74994 > 32'h0000_0009 ? 4'h9 : literal_74994[3:0]];
  assign array_index_74998 = array_update_74995[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_75002 = smul32b_32b_x_32b(array_index_74726[literal_74994 > 32'h0000_0009 ? 4'h9 : literal_74994[3:0]], array_index_74997[add_74992 > 32'h0000_0009 ? 4'h9 : add_74992[3:0]]);
  assign add_75004 = array_index_74998[add_74992 > 32'h0000_0009 ? 4'h9 : add_74992[3:0]] + smul_75002;
  assign array_update_75006[0] = add_74992 == 32'h0000_0000 ? add_75004 : array_index_74998[0];
  assign array_update_75006[1] = add_74992 == 32'h0000_0001 ? add_75004 : array_index_74998[1];
  assign array_update_75006[2] = add_74992 == 32'h0000_0002 ? add_75004 : array_index_74998[2];
  assign array_update_75006[3] = add_74992 == 32'h0000_0003 ? add_75004 : array_index_74998[3];
  assign array_update_75006[4] = add_74992 == 32'h0000_0004 ? add_75004 : array_index_74998[4];
  assign array_update_75006[5] = add_74992 == 32'h0000_0005 ? add_75004 : array_index_74998[5];
  assign array_update_75006[6] = add_74992 == 32'h0000_0006 ? add_75004 : array_index_74998[6];
  assign array_update_75006[7] = add_74992 == 32'h0000_0007 ? add_75004 : array_index_74998[7];
  assign array_update_75006[8] = add_74992 == 32'h0000_0008 ? add_75004 : array_index_74998[8];
  assign array_update_75006[9] = add_74992 == 32'h0000_0009 ? add_75004 : array_index_74998[9];
  assign add_75007 = literal_74994 + 32'h0000_0001;
  assign array_update_75008[0] = add_74719 == 32'h0000_0000 ? array_update_75006 : array_update_74995[0];
  assign array_update_75008[1] = add_74719 == 32'h0000_0001 ? array_update_75006 : array_update_74995[1];
  assign array_update_75008[2] = add_74719 == 32'h0000_0002 ? array_update_75006 : array_update_74995[2];
  assign array_update_75008[3] = add_74719 == 32'h0000_0003 ? array_update_75006 : array_update_74995[3];
  assign array_update_75008[4] = add_74719 == 32'h0000_0004 ? array_update_75006 : array_update_74995[4];
  assign array_update_75008[5] = add_74719 == 32'h0000_0005 ? array_update_75006 : array_update_74995[5];
  assign array_update_75008[6] = add_74719 == 32'h0000_0006 ? array_update_75006 : array_update_74995[6];
  assign array_update_75008[7] = add_74719 == 32'h0000_0007 ? array_update_75006 : array_update_74995[7];
  assign array_update_75008[8] = add_74719 == 32'h0000_0008 ? array_update_75006 : array_update_74995[8];
  assign array_update_75008[9] = add_74719 == 32'h0000_0009 ? array_update_75006 : array_update_74995[9];
  assign array_index_75010 = array_update_72021[add_75007 > 32'h0000_0009 ? 4'h9 : add_75007[3:0]];
  assign array_index_75011 = array_update_75008[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_75015 = smul32b_32b_x_32b(array_index_74726[add_75007 > 32'h0000_0009 ? 4'h9 : add_75007[3:0]], array_index_75010[add_74992 > 32'h0000_0009 ? 4'h9 : add_74992[3:0]]);
  assign add_75017 = array_index_75011[add_74992 > 32'h0000_0009 ? 4'h9 : add_74992[3:0]] + smul_75015;
  assign array_update_75019[0] = add_74992 == 32'h0000_0000 ? add_75017 : array_index_75011[0];
  assign array_update_75019[1] = add_74992 == 32'h0000_0001 ? add_75017 : array_index_75011[1];
  assign array_update_75019[2] = add_74992 == 32'h0000_0002 ? add_75017 : array_index_75011[2];
  assign array_update_75019[3] = add_74992 == 32'h0000_0003 ? add_75017 : array_index_75011[3];
  assign array_update_75019[4] = add_74992 == 32'h0000_0004 ? add_75017 : array_index_75011[4];
  assign array_update_75019[5] = add_74992 == 32'h0000_0005 ? add_75017 : array_index_75011[5];
  assign array_update_75019[6] = add_74992 == 32'h0000_0006 ? add_75017 : array_index_75011[6];
  assign array_update_75019[7] = add_74992 == 32'h0000_0007 ? add_75017 : array_index_75011[7];
  assign array_update_75019[8] = add_74992 == 32'h0000_0008 ? add_75017 : array_index_75011[8];
  assign array_update_75019[9] = add_74992 == 32'h0000_0009 ? add_75017 : array_index_75011[9];
  assign add_75020 = add_75007 + 32'h0000_0001;
  assign array_update_75021[0] = add_74719 == 32'h0000_0000 ? array_update_75019 : array_update_75008[0];
  assign array_update_75021[1] = add_74719 == 32'h0000_0001 ? array_update_75019 : array_update_75008[1];
  assign array_update_75021[2] = add_74719 == 32'h0000_0002 ? array_update_75019 : array_update_75008[2];
  assign array_update_75021[3] = add_74719 == 32'h0000_0003 ? array_update_75019 : array_update_75008[3];
  assign array_update_75021[4] = add_74719 == 32'h0000_0004 ? array_update_75019 : array_update_75008[4];
  assign array_update_75021[5] = add_74719 == 32'h0000_0005 ? array_update_75019 : array_update_75008[5];
  assign array_update_75021[6] = add_74719 == 32'h0000_0006 ? array_update_75019 : array_update_75008[6];
  assign array_update_75021[7] = add_74719 == 32'h0000_0007 ? array_update_75019 : array_update_75008[7];
  assign array_update_75021[8] = add_74719 == 32'h0000_0008 ? array_update_75019 : array_update_75008[8];
  assign array_update_75021[9] = add_74719 == 32'h0000_0009 ? array_update_75019 : array_update_75008[9];
  assign array_index_75023 = array_update_72021[add_75020 > 32'h0000_0009 ? 4'h9 : add_75020[3:0]];
  assign array_index_75024 = array_update_75021[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_75028 = smul32b_32b_x_32b(array_index_74726[add_75020 > 32'h0000_0009 ? 4'h9 : add_75020[3:0]], array_index_75023[add_74992 > 32'h0000_0009 ? 4'h9 : add_74992[3:0]]);
  assign add_75030 = array_index_75024[add_74992 > 32'h0000_0009 ? 4'h9 : add_74992[3:0]] + smul_75028;
  assign array_update_75032[0] = add_74992 == 32'h0000_0000 ? add_75030 : array_index_75024[0];
  assign array_update_75032[1] = add_74992 == 32'h0000_0001 ? add_75030 : array_index_75024[1];
  assign array_update_75032[2] = add_74992 == 32'h0000_0002 ? add_75030 : array_index_75024[2];
  assign array_update_75032[3] = add_74992 == 32'h0000_0003 ? add_75030 : array_index_75024[3];
  assign array_update_75032[4] = add_74992 == 32'h0000_0004 ? add_75030 : array_index_75024[4];
  assign array_update_75032[5] = add_74992 == 32'h0000_0005 ? add_75030 : array_index_75024[5];
  assign array_update_75032[6] = add_74992 == 32'h0000_0006 ? add_75030 : array_index_75024[6];
  assign array_update_75032[7] = add_74992 == 32'h0000_0007 ? add_75030 : array_index_75024[7];
  assign array_update_75032[8] = add_74992 == 32'h0000_0008 ? add_75030 : array_index_75024[8];
  assign array_update_75032[9] = add_74992 == 32'h0000_0009 ? add_75030 : array_index_75024[9];
  assign add_75033 = add_75020 + 32'h0000_0001;
  assign array_update_75034[0] = add_74719 == 32'h0000_0000 ? array_update_75032 : array_update_75021[0];
  assign array_update_75034[1] = add_74719 == 32'h0000_0001 ? array_update_75032 : array_update_75021[1];
  assign array_update_75034[2] = add_74719 == 32'h0000_0002 ? array_update_75032 : array_update_75021[2];
  assign array_update_75034[3] = add_74719 == 32'h0000_0003 ? array_update_75032 : array_update_75021[3];
  assign array_update_75034[4] = add_74719 == 32'h0000_0004 ? array_update_75032 : array_update_75021[4];
  assign array_update_75034[5] = add_74719 == 32'h0000_0005 ? array_update_75032 : array_update_75021[5];
  assign array_update_75034[6] = add_74719 == 32'h0000_0006 ? array_update_75032 : array_update_75021[6];
  assign array_update_75034[7] = add_74719 == 32'h0000_0007 ? array_update_75032 : array_update_75021[7];
  assign array_update_75034[8] = add_74719 == 32'h0000_0008 ? array_update_75032 : array_update_75021[8];
  assign array_update_75034[9] = add_74719 == 32'h0000_0009 ? array_update_75032 : array_update_75021[9];
  assign array_index_75036 = array_update_72021[add_75033 > 32'h0000_0009 ? 4'h9 : add_75033[3:0]];
  assign array_index_75037 = array_update_75034[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_75041 = smul32b_32b_x_32b(array_index_74726[add_75033 > 32'h0000_0009 ? 4'h9 : add_75033[3:0]], array_index_75036[add_74992 > 32'h0000_0009 ? 4'h9 : add_74992[3:0]]);
  assign add_75043 = array_index_75037[add_74992 > 32'h0000_0009 ? 4'h9 : add_74992[3:0]] + smul_75041;
  assign array_update_75045[0] = add_74992 == 32'h0000_0000 ? add_75043 : array_index_75037[0];
  assign array_update_75045[1] = add_74992 == 32'h0000_0001 ? add_75043 : array_index_75037[1];
  assign array_update_75045[2] = add_74992 == 32'h0000_0002 ? add_75043 : array_index_75037[2];
  assign array_update_75045[3] = add_74992 == 32'h0000_0003 ? add_75043 : array_index_75037[3];
  assign array_update_75045[4] = add_74992 == 32'h0000_0004 ? add_75043 : array_index_75037[4];
  assign array_update_75045[5] = add_74992 == 32'h0000_0005 ? add_75043 : array_index_75037[5];
  assign array_update_75045[6] = add_74992 == 32'h0000_0006 ? add_75043 : array_index_75037[6];
  assign array_update_75045[7] = add_74992 == 32'h0000_0007 ? add_75043 : array_index_75037[7];
  assign array_update_75045[8] = add_74992 == 32'h0000_0008 ? add_75043 : array_index_75037[8];
  assign array_update_75045[9] = add_74992 == 32'h0000_0009 ? add_75043 : array_index_75037[9];
  assign add_75046 = add_75033 + 32'h0000_0001;
  assign array_update_75047[0] = add_74719 == 32'h0000_0000 ? array_update_75045 : array_update_75034[0];
  assign array_update_75047[1] = add_74719 == 32'h0000_0001 ? array_update_75045 : array_update_75034[1];
  assign array_update_75047[2] = add_74719 == 32'h0000_0002 ? array_update_75045 : array_update_75034[2];
  assign array_update_75047[3] = add_74719 == 32'h0000_0003 ? array_update_75045 : array_update_75034[3];
  assign array_update_75047[4] = add_74719 == 32'h0000_0004 ? array_update_75045 : array_update_75034[4];
  assign array_update_75047[5] = add_74719 == 32'h0000_0005 ? array_update_75045 : array_update_75034[5];
  assign array_update_75047[6] = add_74719 == 32'h0000_0006 ? array_update_75045 : array_update_75034[6];
  assign array_update_75047[7] = add_74719 == 32'h0000_0007 ? array_update_75045 : array_update_75034[7];
  assign array_update_75047[8] = add_74719 == 32'h0000_0008 ? array_update_75045 : array_update_75034[8];
  assign array_update_75047[9] = add_74719 == 32'h0000_0009 ? array_update_75045 : array_update_75034[9];
  assign array_index_75049 = array_update_72021[add_75046 > 32'h0000_0009 ? 4'h9 : add_75046[3:0]];
  assign array_index_75050 = array_update_75047[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_75054 = smul32b_32b_x_32b(array_index_74726[add_75046 > 32'h0000_0009 ? 4'h9 : add_75046[3:0]], array_index_75049[add_74992 > 32'h0000_0009 ? 4'h9 : add_74992[3:0]]);
  assign add_75056 = array_index_75050[add_74992 > 32'h0000_0009 ? 4'h9 : add_74992[3:0]] + smul_75054;
  assign array_update_75058[0] = add_74992 == 32'h0000_0000 ? add_75056 : array_index_75050[0];
  assign array_update_75058[1] = add_74992 == 32'h0000_0001 ? add_75056 : array_index_75050[1];
  assign array_update_75058[2] = add_74992 == 32'h0000_0002 ? add_75056 : array_index_75050[2];
  assign array_update_75058[3] = add_74992 == 32'h0000_0003 ? add_75056 : array_index_75050[3];
  assign array_update_75058[4] = add_74992 == 32'h0000_0004 ? add_75056 : array_index_75050[4];
  assign array_update_75058[5] = add_74992 == 32'h0000_0005 ? add_75056 : array_index_75050[5];
  assign array_update_75058[6] = add_74992 == 32'h0000_0006 ? add_75056 : array_index_75050[6];
  assign array_update_75058[7] = add_74992 == 32'h0000_0007 ? add_75056 : array_index_75050[7];
  assign array_update_75058[8] = add_74992 == 32'h0000_0008 ? add_75056 : array_index_75050[8];
  assign array_update_75058[9] = add_74992 == 32'h0000_0009 ? add_75056 : array_index_75050[9];
  assign add_75059 = add_75046 + 32'h0000_0001;
  assign array_update_75060[0] = add_74719 == 32'h0000_0000 ? array_update_75058 : array_update_75047[0];
  assign array_update_75060[1] = add_74719 == 32'h0000_0001 ? array_update_75058 : array_update_75047[1];
  assign array_update_75060[2] = add_74719 == 32'h0000_0002 ? array_update_75058 : array_update_75047[2];
  assign array_update_75060[3] = add_74719 == 32'h0000_0003 ? array_update_75058 : array_update_75047[3];
  assign array_update_75060[4] = add_74719 == 32'h0000_0004 ? array_update_75058 : array_update_75047[4];
  assign array_update_75060[5] = add_74719 == 32'h0000_0005 ? array_update_75058 : array_update_75047[5];
  assign array_update_75060[6] = add_74719 == 32'h0000_0006 ? array_update_75058 : array_update_75047[6];
  assign array_update_75060[7] = add_74719 == 32'h0000_0007 ? array_update_75058 : array_update_75047[7];
  assign array_update_75060[8] = add_74719 == 32'h0000_0008 ? array_update_75058 : array_update_75047[8];
  assign array_update_75060[9] = add_74719 == 32'h0000_0009 ? array_update_75058 : array_update_75047[9];
  assign array_index_75062 = array_update_72021[add_75059 > 32'h0000_0009 ? 4'h9 : add_75059[3:0]];
  assign array_index_75063 = array_update_75060[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_75067 = smul32b_32b_x_32b(array_index_74726[add_75059 > 32'h0000_0009 ? 4'h9 : add_75059[3:0]], array_index_75062[add_74992 > 32'h0000_0009 ? 4'h9 : add_74992[3:0]]);
  assign add_75069 = array_index_75063[add_74992 > 32'h0000_0009 ? 4'h9 : add_74992[3:0]] + smul_75067;
  assign array_update_75071[0] = add_74992 == 32'h0000_0000 ? add_75069 : array_index_75063[0];
  assign array_update_75071[1] = add_74992 == 32'h0000_0001 ? add_75069 : array_index_75063[1];
  assign array_update_75071[2] = add_74992 == 32'h0000_0002 ? add_75069 : array_index_75063[2];
  assign array_update_75071[3] = add_74992 == 32'h0000_0003 ? add_75069 : array_index_75063[3];
  assign array_update_75071[4] = add_74992 == 32'h0000_0004 ? add_75069 : array_index_75063[4];
  assign array_update_75071[5] = add_74992 == 32'h0000_0005 ? add_75069 : array_index_75063[5];
  assign array_update_75071[6] = add_74992 == 32'h0000_0006 ? add_75069 : array_index_75063[6];
  assign array_update_75071[7] = add_74992 == 32'h0000_0007 ? add_75069 : array_index_75063[7];
  assign array_update_75071[8] = add_74992 == 32'h0000_0008 ? add_75069 : array_index_75063[8];
  assign array_update_75071[9] = add_74992 == 32'h0000_0009 ? add_75069 : array_index_75063[9];
  assign add_75072 = add_75059 + 32'h0000_0001;
  assign array_update_75073[0] = add_74719 == 32'h0000_0000 ? array_update_75071 : array_update_75060[0];
  assign array_update_75073[1] = add_74719 == 32'h0000_0001 ? array_update_75071 : array_update_75060[1];
  assign array_update_75073[2] = add_74719 == 32'h0000_0002 ? array_update_75071 : array_update_75060[2];
  assign array_update_75073[3] = add_74719 == 32'h0000_0003 ? array_update_75071 : array_update_75060[3];
  assign array_update_75073[4] = add_74719 == 32'h0000_0004 ? array_update_75071 : array_update_75060[4];
  assign array_update_75073[5] = add_74719 == 32'h0000_0005 ? array_update_75071 : array_update_75060[5];
  assign array_update_75073[6] = add_74719 == 32'h0000_0006 ? array_update_75071 : array_update_75060[6];
  assign array_update_75073[7] = add_74719 == 32'h0000_0007 ? array_update_75071 : array_update_75060[7];
  assign array_update_75073[8] = add_74719 == 32'h0000_0008 ? array_update_75071 : array_update_75060[8];
  assign array_update_75073[9] = add_74719 == 32'h0000_0009 ? array_update_75071 : array_update_75060[9];
  assign array_index_75075 = array_update_72021[add_75072 > 32'h0000_0009 ? 4'h9 : add_75072[3:0]];
  assign array_index_75076 = array_update_75073[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_75080 = smul32b_32b_x_32b(array_index_74726[add_75072 > 32'h0000_0009 ? 4'h9 : add_75072[3:0]], array_index_75075[add_74992 > 32'h0000_0009 ? 4'h9 : add_74992[3:0]]);
  assign add_75082 = array_index_75076[add_74992 > 32'h0000_0009 ? 4'h9 : add_74992[3:0]] + smul_75080;
  assign array_update_75084[0] = add_74992 == 32'h0000_0000 ? add_75082 : array_index_75076[0];
  assign array_update_75084[1] = add_74992 == 32'h0000_0001 ? add_75082 : array_index_75076[1];
  assign array_update_75084[2] = add_74992 == 32'h0000_0002 ? add_75082 : array_index_75076[2];
  assign array_update_75084[3] = add_74992 == 32'h0000_0003 ? add_75082 : array_index_75076[3];
  assign array_update_75084[4] = add_74992 == 32'h0000_0004 ? add_75082 : array_index_75076[4];
  assign array_update_75084[5] = add_74992 == 32'h0000_0005 ? add_75082 : array_index_75076[5];
  assign array_update_75084[6] = add_74992 == 32'h0000_0006 ? add_75082 : array_index_75076[6];
  assign array_update_75084[7] = add_74992 == 32'h0000_0007 ? add_75082 : array_index_75076[7];
  assign array_update_75084[8] = add_74992 == 32'h0000_0008 ? add_75082 : array_index_75076[8];
  assign array_update_75084[9] = add_74992 == 32'h0000_0009 ? add_75082 : array_index_75076[9];
  assign add_75085 = add_75072 + 32'h0000_0001;
  assign array_update_75086[0] = add_74719 == 32'h0000_0000 ? array_update_75084 : array_update_75073[0];
  assign array_update_75086[1] = add_74719 == 32'h0000_0001 ? array_update_75084 : array_update_75073[1];
  assign array_update_75086[2] = add_74719 == 32'h0000_0002 ? array_update_75084 : array_update_75073[2];
  assign array_update_75086[3] = add_74719 == 32'h0000_0003 ? array_update_75084 : array_update_75073[3];
  assign array_update_75086[4] = add_74719 == 32'h0000_0004 ? array_update_75084 : array_update_75073[4];
  assign array_update_75086[5] = add_74719 == 32'h0000_0005 ? array_update_75084 : array_update_75073[5];
  assign array_update_75086[6] = add_74719 == 32'h0000_0006 ? array_update_75084 : array_update_75073[6];
  assign array_update_75086[7] = add_74719 == 32'h0000_0007 ? array_update_75084 : array_update_75073[7];
  assign array_update_75086[8] = add_74719 == 32'h0000_0008 ? array_update_75084 : array_update_75073[8];
  assign array_update_75086[9] = add_74719 == 32'h0000_0009 ? array_update_75084 : array_update_75073[9];
  assign array_index_75088 = array_update_72021[add_75085 > 32'h0000_0009 ? 4'h9 : add_75085[3:0]];
  assign array_index_75089 = array_update_75086[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_75093 = smul32b_32b_x_32b(array_index_74726[add_75085 > 32'h0000_0009 ? 4'h9 : add_75085[3:0]], array_index_75088[add_74992 > 32'h0000_0009 ? 4'h9 : add_74992[3:0]]);
  assign add_75095 = array_index_75089[add_74992 > 32'h0000_0009 ? 4'h9 : add_74992[3:0]] + smul_75093;
  assign array_update_75097[0] = add_74992 == 32'h0000_0000 ? add_75095 : array_index_75089[0];
  assign array_update_75097[1] = add_74992 == 32'h0000_0001 ? add_75095 : array_index_75089[1];
  assign array_update_75097[2] = add_74992 == 32'h0000_0002 ? add_75095 : array_index_75089[2];
  assign array_update_75097[3] = add_74992 == 32'h0000_0003 ? add_75095 : array_index_75089[3];
  assign array_update_75097[4] = add_74992 == 32'h0000_0004 ? add_75095 : array_index_75089[4];
  assign array_update_75097[5] = add_74992 == 32'h0000_0005 ? add_75095 : array_index_75089[5];
  assign array_update_75097[6] = add_74992 == 32'h0000_0006 ? add_75095 : array_index_75089[6];
  assign array_update_75097[7] = add_74992 == 32'h0000_0007 ? add_75095 : array_index_75089[7];
  assign array_update_75097[8] = add_74992 == 32'h0000_0008 ? add_75095 : array_index_75089[8];
  assign array_update_75097[9] = add_74992 == 32'h0000_0009 ? add_75095 : array_index_75089[9];
  assign add_75098 = add_75085 + 32'h0000_0001;
  assign array_update_75099[0] = add_74719 == 32'h0000_0000 ? array_update_75097 : array_update_75086[0];
  assign array_update_75099[1] = add_74719 == 32'h0000_0001 ? array_update_75097 : array_update_75086[1];
  assign array_update_75099[2] = add_74719 == 32'h0000_0002 ? array_update_75097 : array_update_75086[2];
  assign array_update_75099[3] = add_74719 == 32'h0000_0003 ? array_update_75097 : array_update_75086[3];
  assign array_update_75099[4] = add_74719 == 32'h0000_0004 ? array_update_75097 : array_update_75086[4];
  assign array_update_75099[5] = add_74719 == 32'h0000_0005 ? array_update_75097 : array_update_75086[5];
  assign array_update_75099[6] = add_74719 == 32'h0000_0006 ? array_update_75097 : array_update_75086[6];
  assign array_update_75099[7] = add_74719 == 32'h0000_0007 ? array_update_75097 : array_update_75086[7];
  assign array_update_75099[8] = add_74719 == 32'h0000_0008 ? array_update_75097 : array_update_75086[8];
  assign array_update_75099[9] = add_74719 == 32'h0000_0009 ? array_update_75097 : array_update_75086[9];
  assign array_index_75101 = array_update_72021[add_75098 > 32'h0000_0009 ? 4'h9 : add_75098[3:0]];
  assign array_index_75102 = array_update_75099[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_75106 = smul32b_32b_x_32b(array_index_74726[add_75098 > 32'h0000_0009 ? 4'h9 : add_75098[3:0]], array_index_75101[add_74992 > 32'h0000_0009 ? 4'h9 : add_74992[3:0]]);
  assign add_75108 = array_index_75102[add_74992 > 32'h0000_0009 ? 4'h9 : add_74992[3:0]] + smul_75106;
  assign array_update_75110[0] = add_74992 == 32'h0000_0000 ? add_75108 : array_index_75102[0];
  assign array_update_75110[1] = add_74992 == 32'h0000_0001 ? add_75108 : array_index_75102[1];
  assign array_update_75110[2] = add_74992 == 32'h0000_0002 ? add_75108 : array_index_75102[2];
  assign array_update_75110[3] = add_74992 == 32'h0000_0003 ? add_75108 : array_index_75102[3];
  assign array_update_75110[4] = add_74992 == 32'h0000_0004 ? add_75108 : array_index_75102[4];
  assign array_update_75110[5] = add_74992 == 32'h0000_0005 ? add_75108 : array_index_75102[5];
  assign array_update_75110[6] = add_74992 == 32'h0000_0006 ? add_75108 : array_index_75102[6];
  assign array_update_75110[7] = add_74992 == 32'h0000_0007 ? add_75108 : array_index_75102[7];
  assign array_update_75110[8] = add_74992 == 32'h0000_0008 ? add_75108 : array_index_75102[8];
  assign array_update_75110[9] = add_74992 == 32'h0000_0009 ? add_75108 : array_index_75102[9];
  assign add_75111 = add_75098 + 32'h0000_0001;
  assign array_update_75112[0] = add_74719 == 32'h0000_0000 ? array_update_75110 : array_update_75099[0];
  assign array_update_75112[1] = add_74719 == 32'h0000_0001 ? array_update_75110 : array_update_75099[1];
  assign array_update_75112[2] = add_74719 == 32'h0000_0002 ? array_update_75110 : array_update_75099[2];
  assign array_update_75112[3] = add_74719 == 32'h0000_0003 ? array_update_75110 : array_update_75099[3];
  assign array_update_75112[4] = add_74719 == 32'h0000_0004 ? array_update_75110 : array_update_75099[4];
  assign array_update_75112[5] = add_74719 == 32'h0000_0005 ? array_update_75110 : array_update_75099[5];
  assign array_update_75112[6] = add_74719 == 32'h0000_0006 ? array_update_75110 : array_update_75099[6];
  assign array_update_75112[7] = add_74719 == 32'h0000_0007 ? array_update_75110 : array_update_75099[7];
  assign array_update_75112[8] = add_74719 == 32'h0000_0008 ? array_update_75110 : array_update_75099[8];
  assign array_update_75112[9] = add_74719 == 32'h0000_0009 ? array_update_75110 : array_update_75099[9];
  assign array_index_75114 = array_update_72021[add_75111 > 32'h0000_0009 ? 4'h9 : add_75111[3:0]];
  assign array_index_75115 = array_update_75112[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_75119 = smul32b_32b_x_32b(array_index_74726[add_75111 > 32'h0000_0009 ? 4'h9 : add_75111[3:0]], array_index_75114[add_74992 > 32'h0000_0009 ? 4'h9 : add_74992[3:0]]);
  assign add_75121 = array_index_75115[add_74992 > 32'h0000_0009 ? 4'h9 : add_74992[3:0]] + smul_75119;
  assign array_update_75122[0] = add_74992 == 32'h0000_0000 ? add_75121 : array_index_75115[0];
  assign array_update_75122[1] = add_74992 == 32'h0000_0001 ? add_75121 : array_index_75115[1];
  assign array_update_75122[2] = add_74992 == 32'h0000_0002 ? add_75121 : array_index_75115[2];
  assign array_update_75122[3] = add_74992 == 32'h0000_0003 ? add_75121 : array_index_75115[3];
  assign array_update_75122[4] = add_74992 == 32'h0000_0004 ? add_75121 : array_index_75115[4];
  assign array_update_75122[5] = add_74992 == 32'h0000_0005 ? add_75121 : array_index_75115[5];
  assign array_update_75122[6] = add_74992 == 32'h0000_0006 ? add_75121 : array_index_75115[6];
  assign array_update_75122[7] = add_74992 == 32'h0000_0007 ? add_75121 : array_index_75115[7];
  assign array_update_75122[8] = add_74992 == 32'h0000_0008 ? add_75121 : array_index_75115[8];
  assign array_update_75122[9] = add_74992 == 32'h0000_0009 ? add_75121 : array_index_75115[9];
  assign array_update_75123[0] = add_74719 == 32'h0000_0000 ? array_update_75122 : array_update_75112[0];
  assign array_update_75123[1] = add_74719 == 32'h0000_0001 ? array_update_75122 : array_update_75112[1];
  assign array_update_75123[2] = add_74719 == 32'h0000_0002 ? array_update_75122 : array_update_75112[2];
  assign array_update_75123[3] = add_74719 == 32'h0000_0003 ? array_update_75122 : array_update_75112[3];
  assign array_update_75123[4] = add_74719 == 32'h0000_0004 ? array_update_75122 : array_update_75112[4];
  assign array_update_75123[5] = add_74719 == 32'h0000_0005 ? array_update_75122 : array_update_75112[5];
  assign array_update_75123[6] = add_74719 == 32'h0000_0006 ? array_update_75122 : array_update_75112[6];
  assign array_update_75123[7] = add_74719 == 32'h0000_0007 ? array_update_75122 : array_update_75112[7];
  assign array_update_75123[8] = add_74719 == 32'h0000_0008 ? array_update_75122 : array_update_75112[8];
  assign array_update_75123[9] = add_74719 == 32'h0000_0009 ? array_update_75122 : array_update_75112[9];
  assign array_index_75125 = array_update_75123[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign add_75127 = add_74992 + 32'h0000_0001;
  assign array_update_75128[0] = add_75127 == 32'h0000_0000 ? 32'h0000_0000 : array_index_75125[0];
  assign array_update_75128[1] = add_75127 == 32'h0000_0001 ? 32'h0000_0000 : array_index_75125[1];
  assign array_update_75128[2] = add_75127 == 32'h0000_0002 ? 32'h0000_0000 : array_index_75125[2];
  assign array_update_75128[3] = add_75127 == 32'h0000_0003 ? 32'h0000_0000 : array_index_75125[3];
  assign array_update_75128[4] = add_75127 == 32'h0000_0004 ? 32'h0000_0000 : array_index_75125[4];
  assign array_update_75128[5] = add_75127 == 32'h0000_0005 ? 32'h0000_0000 : array_index_75125[5];
  assign array_update_75128[6] = add_75127 == 32'h0000_0006 ? 32'h0000_0000 : array_index_75125[6];
  assign array_update_75128[7] = add_75127 == 32'h0000_0007 ? 32'h0000_0000 : array_index_75125[7];
  assign array_update_75128[8] = add_75127 == 32'h0000_0008 ? 32'h0000_0000 : array_index_75125[8];
  assign array_update_75128[9] = add_75127 == 32'h0000_0009 ? 32'h0000_0000 : array_index_75125[9];
  assign literal_75129 = 32'h0000_0000;
  assign array_update_75130[0] = add_74719 == 32'h0000_0000 ? array_update_75128 : array_update_75123[0];
  assign array_update_75130[1] = add_74719 == 32'h0000_0001 ? array_update_75128 : array_update_75123[1];
  assign array_update_75130[2] = add_74719 == 32'h0000_0002 ? array_update_75128 : array_update_75123[2];
  assign array_update_75130[3] = add_74719 == 32'h0000_0003 ? array_update_75128 : array_update_75123[3];
  assign array_update_75130[4] = add_74719 == 32'h0000_0004 ? array_update_75128 : array_update_75123[4];
  assign array_update_75130[5] = add_74719 == 32'h0000_0005 ? array_update_75128 : array_update_75123[5];
  assign array_update_75130[6] = add_74719 == 32'h0000_0006 ? array_update_75128 : array_update_75123[6];
  assign array_update_75130[7] = add_74719 == 32'h0000_0007 ? array_update_75128 : array_update_75123[7];
  assign array_update_75130[8] = add_74719 == 32'h0000_0008 ? array_update_75128 : array_update_75123[8];
  assign array_update_75130[9] = add_74719 == 32'h0000_0009 ? array_update_75128 : array_update_75123[9];
  assign array_index_75132 = array_update_72021[literal_75129 > 32'h0000_0009 ? 4'h9 : literal_75129[3:0]];
  assign array_index_75133 = array_update_75130[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_75137 = smul32b_32b_x_32b(array_index_74726[literal_75129 > 32'h0000_0009 ? 4'h9 : literal_75129[3:0]], array_index_75132[add_75127 > 32'h0000_0009 ? 4'h9 : add_75127[3:0]]);
  assign add_75139 = array_index_75133[add_75127 > 32'h0000_0009 ? 4'h9 : add_75127[3:0]] + smul_75137;
  assign array_update_75141[0] = add_75127 == 32'h0000_0000 ? add_75139 : array_index_75133[0];
  assign array_update_75141[1] = add_75127 == 32'h0000_0001 ? add_75139 : array_index_75133[1];
  assign array_update_75141[2] = add_75127 == 32'h0000_0002 ? add_75139 : array_index_75133[2];
  assign array_update_75141[3] = add_75127 == 32'h0000_0003 ? add_75139 : array_index_75133[3];
  assign array_update_75141[4] = add_75127 == 32'h0000_0004 ? add_75139 : array_index_75133[4];
  assign array_update_75141[5] = add_75127 == 32'h0000_0005 ? add_75139 : array_index_75133[5];
  assign array_update_75141[6] = add_75127 == 32'h0000_0006 ? add_75139 : array_index_75133[6];
  assign array_update_75141[7] = add_75127 == 32'h0000_0007 ? add_75139 : array_index_75133[7];
  assign array_update_75141[8] = add_75127 == 32'h0000_0008 ? add_75139 : array_index_75133[8];
  assign array_update_75141[9] = add_75127 == 32'h0000_0009 ? add_75139 : array_index_75133[9];
  assign add_75142 = literal_75129 + 32'h0000_0001;
  assign array_update_75143[0] = add_74719 == 32'h0000_0000 ? array_update_75141 : array_update_75130[0];
  assign array_update_75143[1] = add_74719 == 32'h0000_0001 ? array_update_75141 : array_update_75130[1];
  assign array_update_75143[2] = add_74719 == 32'h0000_0002 ? array_update_75141 : array_update_75130[2];
  assign array_update_75143[3] = add_74719 == 32'h0000_0003 ? array_update_75141 : array_update_75130[3];
  assign array_update_75143[4] = add_74719 == 32'h0000_0004 ? array_update_75141 : array_update_75130[4];
  assign array_update_75143[5] = add_74719 == 32'h0000_0005 ? array_update_75141 : array_update_75130[5];
  assign array_update_75143[6] = add_74719 == 32'h0000_0006 ? array_update_75141 : array_update_75130[6];
  assign array_update_75143[7] = add_74719 == 32'h0000_0007 ? array_update_75141 : array_update_75130[7];
  assign array_update_75143[8] = add_74719 == 32'h0000_0008 ? array_update_75141 : array_update_75130[8];
  assign array_update_75143[9] = add_74719 == 32'h0000_0009 ? array_update_75141 : array_update_75130[9];
  assign array_index_75145 = array_update_72021[add_75142 > 32'h0000_0009 ? 4'h9 : add_75142[3:0]];
  assign array_index_75146 = array_update_75143[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_75150 = smul32b_32b_x_32b(array_index_74726[add_75142 > 32'h0000_0009 ? 4'h9 : add_75142[3:0]], array_index_75145[add_75127 > 32'h0000_0009 ? 4'h9 : add_75127[3:0]]);
  assign add_75152 = array_index_75146[add_75127 > 32'h0000_0009 ? 4'h9 : add_75127[3:0]] + smul_75150;
  assign array_update_75154[0] = add_75127 == 32'h0000_0000 ? add_75152 : array_index_75146[0];
  assign array_update_75154[1] = add_75127 == 32'h0000_0001 ? add_75152 : array_index_75146[1];
  assign array_update_75154[2] = add_75127 == 32'h0000_0002 ? add_75152 : array_index_75146[2];
  assign array_update_75154[3] = add_75127 == 32'h0000_0003 ? add_75152 : array_index_75146[3];
  assign array_update_75154[4] = add_75127 == 32'h0000_0004 ? add_75152 : array_index_75146[4];
  assign array_update_75154[5] = add_75127 == 32'h0000_0005 ? add_75152 : array_index_75146[5];
  assign array_update_75154[6] = add_75127 == 32'h0000_0006 ? add_75152 : array_index_75146[6];
  assign array_update_75154[7] = add_75127 == 32'h0000_0007 ? add_75152 : array_index_75146[7];
  assign array_update_75154[8] = add_75127 == 32'h0000_0008 ? add_75152 : array_index_75146[8];
  assign array_update_75154[9] = add_75127 == 32'h0000_0009 ? add_75152 : array_index_75146[9];
  assign add_75155 = add_75142 + 32'h0000_0001;
  assign array_update_75156[0] = add_74719 == 32'h0000_0000 ? array_update_75154 : array_update_75143[0];
  assign array_update_75156[1] = add_74719 == 32'h0000_0001 ? array_update_75154 : array_update_75143[1];
  assign array_update_75156[2] = add_74719 == 32'h0000_0002 ? array_update_75154 : array_update_75143[2];
  assign array_update_75156[3] = add_74719 == 32'h0000_0003 ? array_update_75154 : array_update_75143[3];
  assign array_update_75156[4] = add_74719 == 32'h0000_0004 ? array_update_75154 : array_update_75143[4];
  assign array_update_75156[5] = add_74719 == 32'h0000_0005 ? array_update_75154 : array_update_75143[5];
  assign array_update_75156[6] = add_74719 == 32'h0000_0006 ? array_update_75154 : array_update_75143[6];
  assign array_update_75156[7] = add_74719 == 32'h0000_0007 ? array_update_75154 : array_update_75143[7];
  assign array_update_75156[8] = add_74719 == 32'h0000_0008 ? array_update_75154 : array_update_75143[8];
  assign array_update_75156[9] = add_74719 == 32'h0000_0009 ? array_update_75154 : array_update_75143[9];
  assign array_index_75158 = array_update_72021[add_75155 > 32'h0000_0009 ? 4'h9 : add_75155[3:0]];
  assign array_index_75159 = array_update_75156[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_75163 = smul32b_32b_x_32b(array_index_74726[add_75155 > 32'h0000_0009 ? 4'h9 : add_75155[3:0]], array_index_75158[add_75127 > 32'h0000_0009 ? 4'h9 : add_75127[3:0]]);
  assign add_75165 = array_index_75159[add_75127 > 32'h0000_0009 ? 4'h9 : add_75127[3:0]] + smul_75163;
  assign array_update_75167[0] = add_75127 == 32'h0000_0000 ? add_75165 : array_index_75159[0];
  assign array_update_75167[1] = add_75127 == 32'h0000_0001 ? add_75165 : array_index_75159[1];
  assign array_update_75167[2] = add_75127 == 32'h0000_0002 ? add_75165 : array_index_75159[2];
  assign array_update_75167[3] = add_75127 == 32'h0000_0003 ? add_75165 : array_index_75159[3];
  assign array_update_75167[4] = add_75127 == 32'h0000_0004 ? add_75165 : array_index_75159[4];
  assign array_update_75167[5] = add_75127 == 32'h0000_0005 ? add_75165 : array_index_75159[5];
  assign array_update_75167[6] = add_75127 == 32'h0000_0006 ? add_75165 : array_index_75159[6];
  assign array_update_75167[7] = add_75127 == 32'h0000_0007 ? add_75165 : array_index_75159[7];
  assign array_update_75167[8] = add_75127 == 32'h0000_0008 ? add_75165 : array_index_75159[8];
  assign array_update_75167[9] = add_75127 == 32'h0000_0009 ? add_75165 : array_index_75159[9];
  assign add_75168 = add_75155 + 32'h0000_0001;
  assign array_update_75169[0] = add_74719 == 32'h0000_0000 ? array_update_75167 : array_update_75156[0];
  assign array_update_75169[1] = add_74719 == 32'h0000_0001 ? array_update_75167 : array_update_75156[1];
  assign array_update_75169[2] = add_74719 == 32'h0000_0002 ? array_update_75167 : array_update_75156[2];
  assign array_update_75169[3] = add_74719 == 32'h0000_0003 ? array_update_75167 : array_update_75156[3];
  assign array_update_75169[4] = add_74719 == 32'h0000_0004 ? array_update_75167 : array_update_75156[4];
  assign array_update_75169[5] = add_74719 == 32'h0000_0005 ? array_update_75167 : array_update_75156[5];
  assign array_update_75169[6] = add_74719 == 32'h0000_0006 ? array_update_75167 : array_update_75156[6];
  assign array_update_75169[7] = add_74719 == 32'h0000_0007 ? array_update_75167 : array_update_75156[7];
  assign array_update_75169[8] = add_74719 == 32'h0000_0008 ? array_update_75167 : array_update_75156[8];
  assign array_update_75169[9] = add_74719 == 32'h0000_0009 ? array_update_75167 : array_update_75156[9];
  assign array_index_75171 = array_update_72021[add_75168 > 32'h0000_0009 ? 4'h9 : add_75168[3:0]];
  assign array_index_75172 = array_update_75169[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_75176 = smul32b_32b_x_32b(array_index_74726[add_75168 > 32'h0000_0009 ? 4'h9 : add_75168[3:0]], array_index_75171[add_75127 > 32'h0000_0009 ? 4'h9 : add_75127[3:0]]);
  assign add_75178 = array_index_75172[add_75127 > 32'h0000_0009 ? 4'h9 : add_75127[3:0]] + smul_75176;
  assign array_update_75180[0] = add_75127 == 32'h0000_0000 ? add_75178 : array_index_75172[0];
  assign array_update_75180[1] = add_75127 == 32'h0000_0001 ? add_75178 : array_index_75172[1];
  assign array_update_75180[2] = add_75127 == 32'h0000_0002 ? add_75178 : array_index_75172[2];
  assign array_update_75180[3] = add_75127 == 32'h0000_0003 ? add_75178 : array_index_75172[3];
  assign array_update_75180[4] = add_75127 == 32'h0000_0004 ? add_75178 : array_index_75172[4];
  assign array_update_75180[5] = add_75127 == 32'h0000_0005 ? add_75178 : array_index_75172[5];
  assign array_update_75180[6] = add_75127 == 32'h0000_0006 ? add_75178 : array_index_75172[6];
  assign array_update_75180[7] = add_75127 == 32'h0000_0007 ? add_75178 : array_index_75172[7];
  assign array_update_75180[8] = add_75127 == 32'h0000_0008 ? add_75178 : array_index_75172[8];
  assign array_update_75180[9] = add_75127 == 32'h0000_0009 ? add_75178 : array_index_75172[9];
  assign add_75181 = add_75168 + 32'h0000_0001;
  assign array_update_75182[0] = add_74719 == 32'h0000_0000 ? array_update_75180 : array_update_75169[0];
  assign array_update_75182[1] = add_74719 == 32'h0000_0001 ? array_update_75180 : array_update_75169[1];
  assign array_update_75182[2] = add_74719 == 32'h0000_0002 ? array_update_75180 : array_update_75169[2];
  assign array_update_75182[3] = add_74719 == 32'h0000_0003 ? array_update_75180 : array_update_75169[3];
  assign array_update_75182[4] = add_74719 == 32'h0000_0004 ? array_update_75180 : array_update_75169[4];
  assign array_update_75182[5] = add_74719 == 32'h0000_0005 ? array_update_75180 : array_update_75169[5];
  assign array_update_75182[6] = add_74719 == 32'h0000_0006 ? array_update_75180 : array_update_75169[6];
  assign array_update_75182[7] = add_74719 == 32'h0000_0007 ? array_update_75180 : array_update_75169[7];
  assign array_update_75182[8] = add_74719 == 32'h0000_0008 ? array_update_75180 : array_update_75169[8];
  assign array_update_75182[9] = add_74719 == 32'h0000_0009 ? array_update_75180 : array_update_75169[9];
  assign array_index_75184 = array_update_72021[add_75181 > 32'h0000_0009 ? 4'h9 : add_75181[3:0]];
  assign array_index_75185 = array_update_75182[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_75189 = smul32b_32b_x_32b(array_index_74726[add_75181 > 32'h0000_0009 ? 4'h9 : add_75181[3:0]], array_index_75184[add_75127 > 32'h0000_0009 ? 4'h9 : add_75127[3:0]]);
  assign add_75191 = array_index_75185[add_75127 > 32'h0000_0009 ? 4'h9 : add_75127[3:0]] + smul_75189;
  assign array_update_75193[0] = add_75127 == 32'h0000_0000 ? add_75191 : array_index_75185[0];
  assign array_update_75193[1] = add_75127 == 32'h0000_0001 ? add_75191 : array_index_75185[1];
  assign array_update_75193[2] = add_75127 == 32'h0000_0002 ? add_75191 : array_index_75185[2];
  assign array_update_75193[3] = add_75127 == 32'h0000_0003 ? add_75191 : array_index_75185[3];
  assign array_update_75193[4] = add_75127 == 32'h0000_0004 ? add_75191 : array_index_75185[4];
  assign array_update_75193[5] = add_75127 == 32'h0000_0005 ? add_75191 : array_index_75185[5];
  assign array_update_75193[6] = add_75127 == 32'h0000_0006 ? add_75191 : array_index_75185[6];
  assign array_update_75193[7] = add_75127 == 32'h0000_0007 ? add_75191 : array_index_75185[7];
  assign array_update_75193[8] = add_75127 == 32'h0000_0008 ? add_75191 : array_index_75185[8];
  assign array_update_75193[9] = add_75127 == 32'h0000_0009 ? add_75191 : array_index_75185[9];
  assign add_75194 = add_75181 + 32'h0000_0001;
  assign array_update_75195[0] = add_74719 == 32'h0000_0000 ? array_update_75193 : array_update_75182[0];
  assign array_update_75195[1] = add_74719 == 32'h0000_0001 ? array_update_75193 : array_update_75182[1];
  assign array_update_75195[2] = add_74719 == 32'h0000_0002 ? array_update_75193 : array_update_75182[2];
  assign array_update_75195[3] = add_74719 == 32'h0000_0003 ? array_update_75193 : array_update_75182[3];
  assign array_update_75195[4] = add_74719 == 32'h0000_0004 ? array_update_75193 : array_update_75182[4];
  assign array_update_75195[5] = add_74719 == 32'h0000_0005 ? array_update_75193 : array_update_75182[5];
  assign array_update_75195[6] = add_74719 == 32'h0000_0006 ? array_update_75193 : array_update_75182[6];
  assign array_update_75195[7] = add_74719 == 32'h0000_0007 ? array_update_75193 : array_update_75182[7];
  assign array_update_75195[8] = add_74719 == 32'h0000_0008 ? array_update_75193 : array_update_75182[8];
  assign array_update_75195[9] = add_74719 == 32'h0000_0009 ? array_update_75193 : array_update_75182[9];
  assign array_index_75197 = array_update_72021[add_75194 > 32'h0000_0009 ? 4'h9 : add_75194[3:0]];
  assign array_index_75198 = array_update_75195[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_75202 = smul32b_32b_x_32b(array_index_74726[add_75194 > 32'h0000_0009 ? 4'h9 : add_75194[3:0]], array_index_75197[add_75127 > 32'h0000_0009 ? 4'h9 : add_75127[3:0]]);
  assign add_75204 = array_index_75198[add_75127 > 32'h0000_0009 ? 4'h9 : add_75127[3:0]] + smul_75202;
  assign array_update_75206[0] = add_75127 == 32'h0000_0000 ? add_75204 : array_index_75198[0];
  assign array_update_75206[1] = add_75127 == 32'h0000_0001 ? add_75204 : array_index_75198[1];
  assign array_update_75206[2] = add_75127 == 32'h0000_0002 ? add_75204 : array_index_75198[2];
  assign array_update_75206[3] = add_75127 == 32'h0000_0003 ? add_75204 : array_index_75198[3];
  assign array_update_75206[4] = add_75127 == 32'h0000_0004 ? add_75204 : array_index_75198[4];
  assign array_update_75206[5] = add_75127 == 32'h0000_0005 ? add_75204 : array_index_75198[5];
  assign array_update_75206[6] = add_75127 == 32'h0000_0006 ? add_75204 : array_index_75198[6];
  assign array_update_75206[7] = add_75127 == 32'h0000_0007 ? add_75204 : array_index_75198[7];
  assign array_update_75206[8] = add_75127 == 32'h0000_0008 ? add_75204 : array_index_75198[8];
  assign array_update_75206[9] = add_75127 == 32'h0000_0009 ? add_75204 : array_index_75198[9];
  assign add_75207 = add_75194 + 32'h0000_0001;
  assign array_update_75208[0] = add_74719 == 32'h0000_0000 ? array_update_75206 : array_update_75195[0];
  assign array_update_75208[1] = add_74719 == 32'h0000_0001 ? array_update_75206 : array_update_75195[1];
  assign array_update_75208[2] = add_74719 == 32'h0000_0002 ? array_update_75206 : array_update_75195[2];
  assign array_update_75208[3] = add_74719 == 32'h0000_0003 ? array_update_75206 : array_update_75195[3];
  assign array_update_75208[4] = add_74719 == 32'h0000_0004 ? array_update_75206 : array_update_75195[4];
  assign array_update_75208[5] = add_74719 == 32'h0000_0005 ? array_update_75206 : array_update_75195[5];
  assign array_update_75208[6] = add_74719 == 32'h0000_0006 ? array_update_75206 : array_update_75195[6];
  assign array_update_75208[7] = add_74719 == 32'h0000_0007 ? array_update_75206 : array_update_75195[7];
  assign array_update_75208[8] = add_74719 == 32'h0000_0008 ? array_update_75206 : array_update_75195[8];
  assign array_update_75208[9] = add_74719 == 32'h0000_0009 ? array_update_75206 : array_update_75195[9];
  assign array_index_75210 = array_update_72021[add_75207 > 32'h0000_0009 ? 4'h9 : add_75207[3:0]];
  assign array_index_75211 = array_update_75208[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_75215 = smul32b_32b_x_32b(array_index_74726[add_75207 > 32'h0000_0009 ? 4'h9 : add_75207[3:0]], array_index_75210[add_75127 > 32'h0000_0009 ? 4'h9 : add_75127[3:0]]);
  assign add_75217 = array_index_75211[add_75127 > 32'h0000_0009 ? 4'h9 : add_75127[3:0]] + smul_75215;
  assign array_update_75219[0] = add_75127 == 32'h0000_0000 ? add_75217 : array_index_75211[0];
  assign array_update_75219[1] = add_75127 == 32'h0000_0001 ? add_75217 : array_index_75211[1];
  assign array_update_75219[2] = add_75127 == 32'h0000_0002 ? add_75217 : array_index_75211[2];
  assign array_update_75219[3] = add_75127 == 32'h0000_0003 ? add_75217 : array_index_75211[3];
  assign array_update_75219[4] = add_75127 == 32'h0000_0004 ? add_75217 : array_index_75211[4];
  assign array_update_75219[5] = add_75127 == 32'h0000_0005 ? add_75217 : array_index_75211[5];
  assign array_update_75219[6] = add_75127 == 32'h0000_0006 ? add_75217 : array_index_75211[6];
  assign array_update_75219[7] = add_75127 == 32'h0000_0007 ? add_75217 : array_index_75211[7];
  assign array_update_75219[8] = add_75127 == 32'h0000_0008 ? add_75217 : array_index_75211[8];
  assign array_update_75219[9] = add_75127 == 32'h0000_0009 ? add_75217 : array_index_75211[9];
  assign add_75220 = add_75207 + 32'h0000_0001;
  assign array_update_75221[0] = add_74719 == 32'h0000_0000 ? array_update_75219 : array_update_75208[0];
  assign array_update_75221[1] = add_74719 == 32'h0000_0001 ? array_update_75219 : array_update_75208[1];
  assign array_update_75221[2] = add_74719 == 32'h0000_0002 ? array_update_75219 : array_update_75208[2];
  assign array_update_75221[3] = add_74719 == 32'h0000_0003 ? array_update_75219 : array_update_75208[3];
  assign array_update_75221[4] = add_74719 == 32'h0000_0004 ? array_update_75219 : array_update_75208[4];
  assign array_update_75221[5] = add_74719 == 32'h0000_0005 ? array_update_75219 : array_update_75208[5];
  assign array_update_75221[6] = add_74719 == 32'h0000_0006 ? array_update_75219 : array_update_75208[6];
  assign array_update_75221[7] = add_74719 == 32'h0000_0007 ? array_update_75219 : array_update_75208[7];
  assign array_update_75221[8] = add_74719 == 32'h0000_0008 ? array_update_75219 : array_update_75208[8];
  assign array_update_75221[9] = add_74719 == 32'h0000_0009 ? array_update_75219 : array_update_75208[9];
  assign array_index_75223 = array_update_72021[add_75220 > 32'h0000_0009 ? 4'h9 : add_75220[3:0]];
  assign array_index_75224 = array_update_75221[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_75228 = smul32b_32b_x_32b(array_index_74726[add_75220 > 32'h0000_0009 ? 4'h9 : add_75220[3:0]], array_index_75223[add_75127 > 32'h0000_0009 ? 4'h9 : add_75127[3:0]]);
  assign add_75230 = array_index_75224[add_75127 > 32'h0000_0009 ? 4'h9 : add_75127[3:0]] + smul_75228;
  assign array_update_75232[0] = add_75127 == 32'h0000_0000 ? add_75230 : array_index_75224[0];
  assign array_update_75232[1] = add_75127 == 32'h0000_0001 ? add_75230 : array_index_75224[1];
  assign array_update_75232[2] = add_75127 == 32'h0000_0002 ? add_75230 : array_index_75224[2];
  assign array_update_75232[3] = add_75127 == 32'h0000_0003 ? add_75230 : array_index_75224[3];
  assign array_update_75232[4] = add_75127 == 32'h0000_0004 ? add_75230 : array_index_75224[4];
  assign array_update_75232[5] = add_75127 == 32'h0000_0005 ? add_75230 : array_index_75224[5];
  assign array_update_75232[6] = add_75127 == 32'h0000_0006 ? add_75230 : array_index_75224[6];
  assign array_update_75232[7] = add_75127 == 32'h0000_0007 ? add_75230 : array_index_75224[7];
  assign array_update_75232[8] = add_75127 == 32'h0000_0008 ? add_75230 : array_index_75224[8];
  assign array_update_75232[9] = add_75127 == 32'h0000_0009 ? add_75230 : array_index_75224[9];
  assign add_75233 = add_75220 + 32'h0000_0001;
  assign array_update_75234[0] = add_74719 == 32'h0000_0000 ? array_update_75232 : array_update_75221[0];
  assign array_update_75234[1] = add_74719 == 32'h0000_0001 ? array_update_75232 : array_update_75221[1];
  assign array_update_75234[2] = add_74719 == 32'h0000_0002 ? array_update_75232 : array_update_75221[2];
  assign array_update_75234[3] = add_74719 == 32'h0000_0003 ? array_update_75232 : array_update_75221[3];
  assign array_update_75234[4] = add_74719 == 32'h0000_0004 ? array_update_75232 : array_update_75221[4];
  assign array_update_75234[5] = add_74719 == 32'h0000_0005 ? array_update_75232 : array_update_75221[5];
  assign array_update_75234[6] = add_74719 == 32'h0000_0006 ? array_update_75232 : array_update_75221[6];
  assign array_update_75234[7] = add_74719 == 32'h0000_0007 ? array_update_75232 : array_update_75221[7];
  assign array_update_75234[8] = add_74719 == 32'h0000_0008 ? array_update_75232 : array_update_75221[8];
  assign array_update_75234[9] = add_74719 == 32'h0000_0009 ? array_update_75232 : array_update_75221[9];
  assign array_index_75236 = array_update_72021[add_75233 > 32'h0000_0009 ? 4'h9 : add_75233[3:0]];
  assign array_index_75237 = array_update_75234[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_75241 = smul32b_32b_x_32b(array_index_74726[add_75233 > 32'h0000_0009 ? 4'h9 : add_75233[3:0]], array_index_75236[add_75127 > 32'h0000_0009 ? 4'h9 : add_75127[3:0]]);
  assign add_75243 = array_index_75237[add_75127 > 32'h0000_0009 ? 4'h9 : add_75127[3:0]] + smul_75241;
  assign array_update_75245[0] = add_75127 == 32'h0000_0000 ? add_75243 : array_index_75237[0];
  assign array_update_75245[1] = add_75127 == 32'h0000_0001 ? add_75243 : array_index_75237[1];
  assign array_update_75245[2] = add_75127 == 32'h0000_0002 ? add_75243 : array_index_75237[2];
  assign array_update_75245[3] = add_75127 == 32'h0000_0003 ? add_75243 : array_index_75237[3];
  assign array_update_75245[4] = add_75127 == 32'h0000_0004 ? add_75243 : array_index_75237[4];
  assign array_update_75245[5] = add_75127 == 32'h0000_0005 ? add_75243 : array_index_75237[5];
  assign array_update_75245[6] = add_75127 == 32'h0000_0006 ? add_75243 : array_index_75237[6];
  assign array_update_75245[7] = add_75127 == 32'h0000_0007 ? add_75243 : array_index_75237[7];
  assign array_update_75245[8] = add_75127 == 32'h0000_0008 ? add_75243 : array_index_75237[8];
  assign array_update_75245[9] = add_75127 == 32'h0000_0009 ? add_75243 : array_index_75237[9];
  assign add_75246 = add_75233 + 32'h0000_0001;
  assign array_update_75247[0] = add_74719 == 32'h0000_0000 ? array_update_75245 : array_update_75234[0];
  assign array_update_75247[1] = add_74719 == 32'h0000_0001 ? array_update_75245 : array_update_75234[1];
  assign array_update_75247[2] = add_74719 == 32'h0000_0002 ? array_update_75245 : array_update_75234[2];
  assign array_update_75247[3] = add_74719 == 32'h0000_0003 ? array_update_75245 : array_update_75234[3];
  assign array_update_75247[4] = add_74719 == 32'h0000_0004 ? array_update_75245 : array_update_75234[4];
  assign array_update_75247[5] = add_74719 == 32'h0000_0005 ? array_update_75245 : array_update_75234[5];
  assign array_update_75247[6] = add_74719 == 32'h0000_0006 ? array_update_75245 : array_update_75234[6];
  assign array_update_75247[7] = add_74719 == 32'h0000_0007 ? array_update_75245 : array_update_75234[7];
  assign array_update_75247[8] = add_74719 == 32'h0000_0008 ? array_update_75245 : array_update_75234[8];
  assign array_update_75247[9] = add_74719 == 32'h0000_0009 ? array_update_75245 : array_update_75234[9];
  assign array_index_75249 = array_update_72021[add_75246 > 32'h0000_0009 ? 4'h9 : add_75246[3:0]];
  assign array_index_75250 = array_update_75247[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_75254 = smul32b_32b_x_32b(array_index_74726[add_75246 > 32'h0000_0009 ? 4'h9 : add_75246[3:0]], array_index_75249[add_75127 > 32'h0000_0009 ? 4'h9 : add_75127[3:0]]);
  assign add_75256 = array_index_75250[add_75127 > 32'h0000_0009 ? 4'h9 : add_75127[3:0]] + smul_75254;
  assign array_update_75257[0] = add_75127 == 32'h0000_0000 ? add_75256 : array_index_75250[0];
  assign array_update_75257[1] = add_75127 == 32'h0000_0001 ? add_75256 : array_index_75250[1];
  assign array_update_75257[2] = add_75127 == 32'h0000_0002 ? add_75256 : array_index_75250[2];
  assign array_update_75257[3] = add_75127 == 32'h0000_0003 ? add_75256 : array_index_75250[3];
  assign array_update_75257[4] = add_75127 == 32'h0000_0004 ? add_75256 : array_index_75250[4];
  assign array_update_75257[5] = add_75127 == 32'h0000_0005 ? add_75256 : array_index_75250[5];
  assign array_update_75257[6] = add_75127 == 32'h0000_0006 ? add_75256 : array_index_75250[6];
  assign array_update_75257[7] = add_75127 == 32'h0000_0007 ? add_75256 : array_index_75250[7];
  assign array_update_75257[8] = add_75127 == 32'h0000_0008 ? add_75256 : array_index_75250[8];
  assign array_update_75257[9] = add_75127 == 32'h0000_0009 ? add_75256 : array_index_75250[9];
  assign array_update_75258[0] = add_74719 == 32'h0000_0000 ? array_update_75257 : array_update_75247[0];
  assign array_update_75258[1] = add_74719 == 32'h0000_0001 ? array_update_75257 : array_update_75247[1];
  assign array_update_75258[2] = add_74719 == 32'h0000_0002 ? array_update_75257 : array_update_75247[2];
  assign array_update_75258[3] = add_74719 == 32'h0000_0003 ? array_update_75257 : array_update_75247[3];
  assign array_update_75258[4] = add_74719 == 32'h0000_0004 ? array_update_75257 : array_update_75247[4];
  assign array_update_75258[5] = add_74719 == 32'h0000_0005 ? array_update_75257 : array_update_75247[5];
  assign array_update_75258[6] = add_74719 == 32'h0000_0006 ? array_update_75257 : array_update_75247[6];
  assign array_update_75258[7] = add_74719 == 32'h0000_0007 ? array_update_75257 : array_update_75247[7];
  assign array_update_75258[8] = add_74719 == 32'h0000_0008 ? array_update_75257 : array_update_75247[8];
  assign array_update_75258[9] = add_74719 == 32'h0000_0009 ? array_update_75257 : array_update_75247[9];
  assign array_index_75260 = array_update_75258[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign add_75262 = add_75127 + 32'h0000_0001;
  assign array_update_75263[0] = add_75262 == 32'h0000_0000 ? 32'h0000_0000 : array_index_75260[0];
  assign array_update_75263[1] = add_75262 == 32'h0000_0001 ? 32'h0000_0000 : array_index_75260[1];
  assign array_update_75263[2] = add_75262 == 32'h0000_0002 ? 32'h0000_0000 : array_index_75260[2];
  assign array_update_75263[3] = add_75262 == 32'h0000_0003 ? 32'h0000_0000 : array_index_75260[3];
  assign array_update_75263[4] = add_75262 == 32'h0000_0004 ? 32'h0000_0000 : array_index_75260[4];
  assign array_update_75263[5] = add_75262 == 32'h0000_0005 ? 32'h0000_0000 : array_index_75260[5];
  assign array_update_75263[6] = add_75262 == 32'h0000_0006 ? 32'h0000_0000 : array_index_75260[6];
  assign array_update_75263[7] = add_75262 == 32'h0000_0007 ? 32'h0000_0000 : array_index_75260[7];
  assign array_update_75263[8] = add_75262 == 32'h0000_0008 ? 32'h0000_0000 : array_index_75260[8];
  assign array_update_75263[9] = add_75262 == 32'h0000_0009 ? 32'h0000_0000 : array_index_75260[9];
  assign literal_75264 = 32'h0000_0000;
  assign array_update_75265[0] = add_74719 == 32'h0000_0000 ? array_update_75263 : array_update_75258[0];
  assign array_update_75265[1] = add_74719 == 32'h0000_0001 ? array_update_75263 : array_update_75258[1];
  assign array_update_75265[2] = add_74719 == 32'h0000_0002 ? array_update_75263 : array_update_75258[2];
  assign array_update_75265[3] = add_74719 == 32'h0000_0003 ? array_update_75263 : array_update_75258[3];
  assign array_update_75265[4] = add_74719 == 32'h0000_0004 ? array_update_75263 : array_update_75258[4];
  assign array_update_75265[5] = add_74719 == 32'h0000_0005 ? array_update_75263 : array_update_75258[5];
  assign array_update_75265[6] = add_74719 == 32'h0000_0006 ? array_update_75263 : array_update_75258[6];
  assign array_update_75265[7] = add_74719 == 32'h0000_0007 ? array_update_75263 : array_update_75258[7];
  assign array_update_75265[8] = add_74719 == 32'h0000_0008 ? array_update_75263 : array_update_75258[8];
  assign array_update_75265[9] = add_74719 == 32'h0000_0009 ? array_update_75263 : array_update_75258[9];
  assign array_index_75267 = array_update_72021[literal_75264 > 32'h0000_0009 ? 4'h9 : literal_75264[3:0]];
  assign array_index_75268 = array_update_75265[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_75272 = smul32b_32b_x_32b(array_index_74726[literal_75264 > 32'h0000_0009 ? 4'h9 : literal_75264[3:0]], array_index_75267[add_75262 > 32'h0000_0009 ? 4'h9 : add_75262[3:0]]);
  assign add_75274 = array_index_75268[add_75262 > 32'h0000_0009 ? 4'h9 : add_75262[3:0]] + smul_75272;
  assign array_update_75276[0] = add_75262 == 32'h0000_0000 ? add_75274 : array_index_75268[0];
  assign array_update_75276[1] = add_75262 == 32'h0000_0001 ? add_75274 : array_index_75268[1];
  assign array_update_75276[2] = add_75262 == 32'h0000_0002 ? add_75274 : array_index_75268[2];
  assign array_update_75276[3] = add_75262 == 32'h0000_0003 ? add_75274 : array_index_75268[3];
  assign array_update_75276[4] = add_75262 == 32'h0000_0004 ? add_75274 : array_index_75268[4];
  assign array_update_75276[5] = add_75262 == 32'h0000_0005 ? add_75274 : array_index_75268[5];
  assign array_update_75276[6] = add_75262 == 32'h0000_0006 ? add_75274 : array_index_75268[6];
  assign array_update_75276[7] = add_75262 == 32'h0000_0007 ? add_75274 : array_index_75268[7];
  assign array_update_75276[8] = add_75262 == 32'h0000_0008 ? add_75274 : array_index_75268[8];
  assign array_update_75276[9] = add_75262 == 32'h0000_0009 ? add_75274 : array_index_75268[9];
  assign add_75277 = literal_75264 + 32'h0000_0001;
  assign array_update_75278[0] = add_74719 == 32'h0000_0000 ? array_update_75276 : array_update_75265[0];
  assign array_update_75278[1] = add_74719 == 32'h0000_0001 ? array_update_75276 : array_update_75265[1];
  assign array_update_75278[2] = add_74719 == 32'h0000_0002 ? array_update_75276 : array_update_75265[2];
  assign array_update_75278[3] = add_74719 == 32'h0000_0003 ? array_update_75276 : array_update_75265[3];
  assign array_update_75278[4] = add_74719 == 32'h0000_0004 ? array_update_75276 : array_update_75265[4];
  assign array_update_75278[5] = add_74719 == 32'h0000_0005 ? array_update_75276 : array_update_75265[5];
  assign array_update_75278[6] = add_74719 == 32'h0000_0006 ? array_update_75276 : array_update_75265[6];
  assign array_update_75278[7] = add_74719 == 32'h0000_0007 ? array_update_75276 : array_update_75265[7];
  assign array_update_75278[8] = add_74719 == 32'h0000_0008 ? array_update_75276 : array_update_75265[8];
  assign array_update_75278[9] = add_74719 == 32'h0000_0009 ? array_update_75276 : array_update_75265[9];
  assign array_index_75280 = array_update_72021[add_75277 > 32'h0000_0009 ? 4'h9 : add_75277[3:0]];
  assign array_index_75281 = array_update_75278[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_75285 = smul32b_32b_x_32b(array_index_74726[add_75277 > 32'h0000_0009 ? 4'h9 : add_75277[3:0]], array_index_75280[add_75262 > 32'h0000_0009 ? 4'h9 : add_75262[3:0]]);
  assign add_75287 = array_index_75281[add_75262 > 32'h0000_0009 ? 4'h9 : add_75262[3:0]] + smul_75285;
  assign array_update_75289[0] = add_75262 == 32'h0000_0000 ? add_75287 : array_index_75281[0];
  assign array_update_75289[1] = add_75262 == 32'h0000_0001 ? add_75287 : array_index_75281[1];
  assign array_update_75289[2] = add_75262 == 32'h0000_0002 ? add_75287 : array_index_75281[2];
  assign array_update_75289[3] = add_75262 == 32'h0000_0003 ? add_75287 : array_index_75281[3];
  assign array_update_75289[4] = add_75262 == 32'h0000_0004 ? add_75287 : array_index_75281[4];
  assign array_update_75289[5] = add_75262 == 32'h0000_0005 ? add_75287 : array_index_75281[5];
  assign array_update_75289[6] = add_75262 == 32'h0000_0006 ? add_75287 : array_index_75281[6];
  assign array_update_75289[7] = add_75262 == 32'h0000_0007 ? add_75287 : array_index_75281[7];
  assign array_update_75289[8] = add_75262 == 32'h0000_0008 ? add_75287 : array_index_75281[8];
  assign array_update_75289[9] = add_75262 == 32'h0000_0009 ? add_75287 : array_index_75281[9];
  assign add_75290 = add_75277 + 32'h0000_0001;
  assign array_update_75291[0] = add_74719 == 32'h0000_0000 ? array_update_75289 : array_update_75278[0];
  assign array_update_75291[1] = add_74719 == 32'h0000_0001 ? array_update_75289 : array_update_75278[1];
  assign array_update_75291[2] = add_74719 == 32'h0000_0002 ? array_update_75289 : array_update_75278[2];
  assign array_update_75291[3] = add_74719 == 32'h0000_0003 ? array_update_75289 : array_update_75278[3];
  assign array_update_75291[4] = add_74719 == 32'h0000_0004 ? array_update_75289 : array_update_75278[4];
  assign array_update_75291[5] = add_74719 == 32'h0000_0005 ? array_update_75289 : array_update_75278[5];
  assign array_update_75291[6] = add_74719 == 32'h0000_0006 ? array_update_75289 : array_update_75278[6];
  assign array_update_75291[7] = add_74719 == 32'h0000_0007 ? array_update_75289 : array_update_75278[7];
  assign array_update_75291[8] = add_74719 == 32'h0000_0008 ? array_update_75289 : array_update_75278[8];
  assign array_update_75291[9] = add_74719 == 32'h0000_0009 ? array_update_75289 : array_update_75278[9];
  assign array_index_75293 = array_update_72021[add_75290 > 32'h0000_0009 ? 4'h9 : add_75290[3:0]];
  assign array_index_75294 = array_update_75291[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_75298 = smul32b_32b_x_32b(array_index_74726[add_75290 > 32'h0000_0009 ? 4'h9 : add_75290[3:0]], array_index_75293[add_75262 > 32'h0000_0009 ? 4'h9 : add_75262[3:0]]);
  assign add_75300 = array_index_75294[add_75262 > 32'h0000_0009 ? 4'h9 : add_75262[3:0]] + smul_75298;
  assign array_update_75302[0] = add_75262 == 32'h0000_0000 ? add_75300 : array_index_75294[0];
  assign array_update_75302[1] = add_75262 == 32'h0000_0001 ? add_75300 : array_index_75294[1];
  assign array_update_75302[2] = add_75262 == 32'h0000_0002 ? add_75300 : array_index_75294[2];
  assign array_update_75302[3] = add_75262 == 32'h0000_0003 ? add_75300 : array_index_75294[3];
  assign array_update_75302[4] = add_75262 == 32'h0000_0004 ? add_75300 : array_index_75294[4];
  assign array_update_75302[5] = add_75262 == 32'h0000_0005 ? add_75300 : array_index_75294[5];
  assign array_update_75302[6] = add_75262 == 32'h0000_0006 ? add_75300 : array_index_75294[6];
  assign array_update_75302[7] = add_75262 == 32'h0000_0007 ? add_75300 : array_index_75294[7];
  assign array_update_75302[8] = add_75262 == 32'h0000_0008 ? add_75300 : array_index_75294[8];
  assign array_update_75302[9] = add_75262 == 32'h0000_0009 ? add_75300 : array_index_75294[9];
  assign add_75303 = add_75290 + 32'h0000_0001;
  assign array_update_75304[0] = add_74719 == 32'h0000_0000 ? array_update_75302 : array_update_75291[0];
  assign array_update_75304[1] = add_74719 == 32'h0000_0001 ? array_update_75302 : array_update_75291[1];
  assign array_update_75304[2] = add_74719 == 32'h0000_0002 ? array_update_75302 : array_update_75291[2];
  assign array_update_75304[3] = add_74719 == 32'h0000_0003 ? array_update_75302 : array_update_75291[3];
  assign array_update_75304[4] = add_74719 == 32'h0000_0004 ? array_update_75302 : array_update_75291[4];
  assign array_update_75304[5] = add_74719 == 32'h0000_0005 ? array_update_75302 : array_update_75291[5];
  assign array_update_75304[6] = add_74719 == 32'h0000_0006 ? array_update_75302 : array_update_75291[6];
  assign array_update_75304[7] = add_74719 == 32'h0000_0007 ? array_update_75302 : array_update_75291[7];
  assign array_update_75304[8] = add_74719 == 32'h0000_0008 ? array_update_75302 : array_update_75291[8];
  assign array_update_75304[9] = add_74719 == 32'h0000_0009 ? array_update_75302 : array_update_75291[9];
  assign array_index_75306 = array_update_72021[add_75303 > 32'h0000_0009 ? 4'h9 : add_75303[3:0]];
  assign array_index_75307 = array_update_75304[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_75311 = smul32b_32b_x_32b(array_index_74726[add_75303 > 32'h0000_0009 ? 4'h9 : add_75303[3:0]], array_index_75306[add_75262 > 32'h0000_0009 ? 4'h9 : add_75262[3:0]]);
  assign add_75313 = array_index_75307[add_75262 > 32'h0000_0009 ? 4'h9 : add_75262[3:0]] + smul_75311;
  assign array_update_75315[0] = add_75262 == 32'h0000_0000 ? add_75313 : array_index_75307[0];
  assign array_update_75315[1] = add_75262 == 32'h0000_0001 ? add_75313 : array_index_75307[1];
  assign array_update_75315[2] = add_75262 == 32'h0000_0002 ? add_75313 : array_index_75307[2];
  assign array_update_75315[3] = add_75262 == 32'h0000_0003 ? add_75313 : array_index_75307[3];
  assign array_update_75315[4] = add_75262 == 32'h0000_0004 ? add_75313 : array_index_75307[4];
  assign array_update_75315[5] = add_75262 == 32'h0000_0005 ? add_75313 : array_index_75307[5];
  assign array_update_75315[6] = add_75262 == 32'h0000_0006 ? add_75313 : array_index_75307[6];
  assign array_update_75315[7] = add_75262 == 32'h0000_0007 ? add_75313 : array_index_75307[7];
  assign array_update_75315[8] = add_75262 == 32'h0000_0008 ? add_75313 : array_index_75307[8];
  assign array_update_75315[9] = add_75262 == 32'h0000_0009 ? add_75313 : array_index_75307[9];
  assign add_75316 = add_75303 + 32'h0000_0001;
  assign array_update_75317[0] = add_74719 == 32'h0000_0000 ? array_update_75315 : array_update_75304[0];
  assign array_update_75317[1] = add_74719 == 32'h0000_0001 ? array_update_75315 : array_update_75304[1];
  assign array_update_75317[2] = add_74719 == 32'h0000_0002 ? array_update_75315 : array_update_75304[2];
  assign array_update_75317[3] = add_74719 == 32'h0000_0003 ? array_update_75315 : array_update_75304[3];
  assign array_update_75317[4] = add_74719 == 32'h0000_0004 ? array_update_75315 : array_update_75304[4];
  assign array_update_75317[5] = add_74719 == 32'h0000_0005 ? array_update_75315 : array_update_75304[5];
  assign array_update_75317[6] = add_74719 == 32'h0000_0006 ? array_update_75315 : array_update_75304[6];
  assign array_update_75317[7] = add_74719 == 32'h0000_0007 ? array_update_75315 : array_update_75304[7];
  assign array_update_75317[8] = add_74719 == 32'h0000_0008 ? array_update_75315 : array_update_75304[8];
  assign array_update_75317[9] = add_74719 == 32'h0000_0009 ? array_update_75315 : array_update_75304[9];
  assign array_index_75319 = array_update_72021[add_75316 > 32'h0000_0009 ? 4'h9 : add_75316[3:0]];
  assign array_index_75320 = array_update_75317[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_75324 = smul32b_32b_x_32b(array_index_74726[add_75316 > 32'h0000_0009 ? 4'h9 : add_75316[3:0]], array_index_75319[add_75262 > 32'h0000_0009 ? 4'h9 : add_75262[3:0]]);
  assign add_75326 = array_index_75320[add_75262 > 32'h0000_0009 ? 4'h9 : add_75262[3:0]] + smul_75324;
  assign array_update_75328[0] = add_75262 == 32'h0000_0000 ? add_75326 : array_index_75320[0];
  assign array_update_75328[1] = add_75262 == 32'h0000_0001 ? add_75326 : array_index_75320[1];
  assign array_update_75328[2] = add_75262 == 32'h0000_0002 ? add_75326 : array_index_75320[2];
  assign array_update_75328[3] = add_75262 == 32'h0000_0003 ? add_75326 : array_index_75320[3];
  assign array_update_75328[4] = add_75262 == 32'h0000_0004 ? add_75326 : array_index_75320[4];
  assign array_update_75328[5] = add_75262 == 32'h0000_0005 ? add_75326 : array_index_75320[5];
  assign array_update_75328[6] = add_75262 == 32'h0000_0006 ? add_75326 : array_index_75320[6];
  assign array_update_75328[7] = add_75262 == 32'h0000_0007 ? add_75326 : array_index_75320[7];
  assign array_update_75328[8] = add_75262 == 32'h0000_0008 ? add_75326 : array_index_75320[8];
  assign array_update_75328[9] = add_75262 == 32'h0000_0009 ? add_75326 : array_index_75320[9];
  assign add_75329 = add_75316 + 32'h0000_0001;
  assign array_update_75330[0] = add_74719 == 32'h0000_0000 ? array_update_75328 : array_update_75317[0];
  assign array_update_75330[1] = add_74719 == 32'h0000_0001 ? array_update_75328 : array_update_75317[1];
  assign array_update_75330[2] = add_74719 == 32'h0000_0002 ? array_update_75328 : array_update_75317[2];
  assign array_update_75330[3] = add_74719 == 32'h0000_0003 ? array_update_75328 : array_update_75317[3];
  assign array_update_75330[4] = add_74719 == 32'h0000_0004 ? array_update_75328 : array_update_75317[4];
  assign array_update_75330[5] = add_74719 == 32'h0000_0005 ? array_update_75328 : array_update_75317[5];
  assign array_update_75330[6] = add_74719 == 32'h0000_0006 ? array_update_75328 : array_update_75317[6];
  assign array_update_75330[7] = add_74719 == 32'h0000_0007 ? array_update_75328 : array_update_75317[7];
  assign array_update_75330[8] = add_74719 == 32'h0000_0008 ? array_update_75328 : array_update_75317[8];
  assign array_update_75330[9] = add_74719 == 32'h0000_0009 ? array_update_75328 : array_update_75317[9];
  assign array_index_75332 = array_update_72021[add_75329 > 32'h0000_0009 ? 4'h9 : add_75329[3:0]];
  assign array_index_75333 = array_update_75330[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_75337 = smul32b_32b_x_32b(array_index_74726[add_75329 > 32'h0000_0009 ? 4'h9 : add_75329[3:0]], array_index_75332[add_75262 > 32'h0000_0009 ? 4'h9 : add_75262[3:0]]);
  assign add_75339 = array_index_75333[add_75262 > 32'h0000_0009 ? 4'h9 : add_75262[3:0]] + smul_75337;
  assign array_update_75341[0] = add_75262 == 32'h0000_0000 ? add_75339 : array_index_75333[0];
  assign array_update_75341[1] = add_75262 == 32'h0000_0001 ? add_75339 : array_index_75333[1];
  assign array_update_75341[2] = add_75262 == 32'h0000_0002 ? add_75339 : array_index_75333[2];
  assign array_update_75341[3] = add_75262 == 32'h0000_0003 ? add_75339 : array_index_75333[3];
  assign array_update_75341[4] = add_75262 == 32'h0000_0004 ? add_75339 : array_index_75333[4];
  assign array_update_75341[5] = add_75262 == 32'h0000_0005 ? add_75339 : array_index_75333[5];
  assign array_update_75341[6] = add_75262 == 32'h0000_0006 ? add_75339 : array_index_75333[6];
  assign array_update_75341[7] = add_75262 == 32'h0000_0007 ? add_75339 : array_index_75333[7];
  assign array_update_75341[8] = add_75262 == 32'h0000_0008 ? add_75339 : array_index_75333[8];
  assign array_update_75341[9] = add_75262 == 32'h0000_0009 ? add_75339 : array_index_75333[9];
  assign add_75342 = add_75329 + 32'h0000_0001;
  assign array_update_75343[0] = add_74719 == 32'h0000_0000 ? array_update_75341 : array_update_75330[0];
  assign array_update_75343[1] = add_74719 == 32'h0000_0001 ? array_update_75341 : array_update_75330[1];
  assign array_update_75343[2] = add_74719 == 32'h0000_0002 ? array_update_75341 : array_update_75330[2];
  assign array_update_75343[3] = add_74719 == 32'h0000_0003 ? array_update_75341 : array_update_75330[3];
  assign array_update_75343[4] = add_74719 == 32'h0000_0004 ? array_update_75341 : array_update_75330[4];
  assign array_update_75343[5] = add_74719 == 32'h0000_0005 ? array_update_75341 : array_update_75330[5];
  assign array_update_75343[6] = add_74719 == 32'h0000_0006 ? array_update_75341 : array_update_75330[6];
  assign array_update_75343[7] = add_74719 == 32'h0000_0007 ? array_update_75341 : array_update_75330[7];
  assign array_update_75343[8] = add_74719 == 32'h0000_0008 ? array_update_75341 : array_update_75330[8];
  assign array_update_75343[9] = add_74719 == 32'h0000_0009 ? array_update_75341 : array_update_75330[9];
  assign array_index_75345 = array_update_72021[add_75342 > 32'h0000_0009 ? 4'h9 : add_75342[3:0]];
  assign array_index_75346 = array_update_75343[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_75350 = smul32b_32b_x_32b(array_index_74726[add_75342 > 32'h0000_0009 ? 4'h9 : add_75342[3:0]], array_index_75345[add_75262 > 32'h0000_0009 ? 4'h9 : add_75262[3:0]]);
  assign add_75352 = array_index_75346[add_75262 > 32'h0000_0009 ? 4'h9 : add_75262[3:0]] + smul_75350;
  assign array_update_75354[0] = add_75262 == 32'h0000_0000 ? add_75352 : array_index_75346[0];
  assign array_update_75354[1] = add_75262 == 32'h0000_0001 ? add_75352 : array_index_75346[1];
  assign array_update_75354[2] = add_75262 == 32'h0000_0002 ? add_75352 : array_index_75346[2];
  assign array_update_75354[3] = add_75262 == 32'h0000_0003 ? add_75352 : array_index_75346[3];
  assign array_update_75354[4] = add_75262 == 32'h0000_0004 ? add_75352 : array_index_75346[4];
  assign array_update_75354[5] = add_75262 == 32'h0000_0005 ? add_75352 : array_index_75346[5];
  assign array_update_75354[6] = add_75262 == 32'h0000_0006 ? add_75352 : array_index_75346[6];
  assign array_update_75354[7] = add_75262 == 32'h0000_0007 ? add_75352 : array_index_75346[7];
  assign array_update_75354[8] = add_75262 == 32'h0000_0008 ? add_75352 : array_index_75346[8];
  assign array_update_75354[9] = add_75262 == 32'h0000_0009 ? add_75352 : array_index_75346[9];
  assign add_75355 = add_75342 + 32'h0000_0001;
  assign array_update_75356[0] = add_74719 == 32'h0000_0000 ? array_update_75354 : array_update_75343[0];
  assign array_update_75356[1] = add_74719 == 32'h0000_0001 ? array_update_75354 : array_update_75343[1];
  assign array_update_75356[2] = add_74719 == 32'h0000_0002 ? array_update_75354 : array_update_75343[2];
  assign array_update_75356[3] = add_74719 == 32'h0000_0003 ? array_update_75354 : array_update_75343[3];
  assign array_update_75356[4] = add_74719 == 32'h0000_0004 ? array_update_75354 : array_update_75343[4];
  assign array_update_75356[5] = add_74719 == 32'h0000_0005 ? array_update_75354 : array_update_75343[5];
  assign array_update_75356[6] = add_74719 == 32'h0000_0006 ? array_update_75354 : array_update_75343[6];
  assign array_update_75356[7] = add_74719 == 32'h0000_0007 ? array_update_75354 : array_update_75343[7];
  assign array_update_75356[8] = add_74719 == 32'h0000_0008 ? array_update_75354 : array_update_75343[8];
  assign array_update_75356[9] = add_74719 == 32'h0000_0009 ? array_update_75354 : array_update_75343[9];
  assign array_index_75358 = array_update_72021[add_75355 > 32'h0000_0009 ? 4'h9 : add_75355[3:0]];
  assign array_index_75359 = array_update_75356[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_75363 = smul32b_32b_x_32b(array_index_74726[add_75355 > 32'h0000_0009 ? 4'h9 : add_75355[3:0]], array_index_75358[add_75262 > 32'h0000_0009 ? 4'h9 : add_75262[3:0]]);
  assign add_75365 = array_index_75359[add_75262 > 32'h0000_0009 ? 4'h9 : add_75262[3:0]] + smul_75363;
  assign array_update_75367[0] = add_75262 == 32'h0000_0000 ? add_75365 : array_index_75359[0];
  assign array_update_75367[1] = add_75262 == 32'h0000_0001 ? add_75365 : array_index_75359[1];
  assign array_update_75367[2] = add_75262 == 32'h0000_0002 ? add_75365 : array_index_75359[2];
  assign array_update_75367[3] = add_75262 == 32'h0000_0003 ? add_75365 : array_index_75359[3];
  assign array_update_75367[4] = add_75262 == 32'h0000_0004 ? add_75365 : array_index_75359[4];
  assign array_update_75367[5] = add_75262 == 32'h0000_0005 ? add_75365 : array_index_75359[5];
  assign array_update_75367[6] = add_75262 == 32'h0000_0006 ? add_75365 : array_index_75359[6];
  assign array_update_75367[7] = add_75262 == 32'h0000_0007 ? add_75365 : array_index_75359[7];
  assign array_update_75367[8] = add_75262 == 32'h0000_0008 ? add_75365 : array_index_75359[8];
  assign array_update_75367[9] = add_75262 == 32'h0000_0009 ? add_75365 : array_index_75359[9];
  assign add_75368 = add_75355 + 32'h0000_0001;
  assign array_update_75369[0] = add_74719 == 32'h0000_0000 ? array_update_75367 : array_update_75356[0];
  assign array_update_75369[1] = add_74719 == 32'h0000_0001 ? array_update_75367 : array_update_75356[1];
  assign array_update_75369[2] = add_74719 == 32'h0000_0002 ? array_update_75367 : array_update_75356[2];
  assign array_update_75369[3] = add_74719 == 32'h0000_0003 ? array_update_75367 : array_update_75356[3];
  assign array_update_75369[4] = add_74719 == 32'h0000_0004 ? array_update_75367 : array_update_75356[4];
  assign array_update_75369[5] = add_74719 == 32'h0000_0005 ? array_update_75367 : array_update_75356[5];
  assign array_update_75369[6] = add_74719 == 32'h0000_0006 ? array_update_75367 : array_update_75356[6];
  assign array_update_75369[7] = add_74719 == 32'h0000_0007 ? array_update_75367 : array_update_75356[7];
  assign array_update_75369[8] = add_74719 == 32'h0000_0008 ? array_update_75367 : array_update_75356[8];
  assign array_update_75369[9] = add_74719 == 32'h0000_0009 ? array_update_75367 : array_update_75356[9];
  assign array_index_75371 = array_update_72021[add_75368 > 32'h0000_0009 ? 4'h9 : add_75368[3:0]];
  assign array_index_75372 = array_update_75369[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_75376 = smul32b_32b_x_32b(array_index_74726[add_75368 > 32'h0000_0009 ? 4'h9 : add_75368[3:0]], array_index_75371[add_75262 > 32'h0000_0009 ? 4'h9 : add_75262[3:0]]);
  assign add_75378 = array_index_75372[add_75262 > 32'h0000_0009 ? 4'h9 : add_75262[3:0]] + smul_75376;
  assign array_update_75380[0] = add_75262 == 32'h0000_0000 ? add_75378 : array_index_75372[0];
  assign array_update_75380[1] = add_75262 == 32'h0000_0001 ? add_75378 : array_index_75372[1];
  assign array_update_75380[2] = add_75262 == 32'h0000_0002 ? add_75378 : array_index_75372[2];
  assign array_update_75380[3] = add_75262 == 32'h0000_0003 ? add_75378 : array_index_75372[3];
  assign array_update_75380[4] = add_75262 == 32'h0000_0004 ? add_75378 : array_index_75372[4];
  assign array_update_75380[5] = add_75262 == 32'h0000_0005 ? add_75378 : array_index_75372[5];
  assign array_update_75380[6] = add_75262 == 32'h0000_0006 ? add_75378 : array_index_75372[6];
  assign array_update_75380[7] = add_75262 == 32'h0000_0007 ? add_75378 : array_index_75372[7];
  assign array_update_75380[8] = add_75262 == 32'h0000_0008 ? add_75378 : array_index_75372[8];
  assign array_update_75380[9] = add_75262 == 32'h0000_0009 ? add_75378 : array_index_75372[9];
  assign add_75381 = add_75368 + 32'h0000_0001;
  assign array_update_75382[0] = add_74719 == 32'h0000_0000 ? array_update_75380 : array_update_75369[0];
  assign array_update_75382[1] = add_74719 == 32'h0000_0001 ? array_update_75380 : array_update_75369[1];
  assign array_update_75382[2] = add_74719 == 32'h0000_0002 ? array_update_75380 : array_update_75369[2];
  assign array_update_75382[3] = add_74719 == 32'h0000_0003 ? array_update_75380 : array_update_75369[3];
  assign array_update_75382[4] = add_74719 == 32'h0000_0004 ? array_update_75380 : array_update_75369[4];
  assign array_update_75382[5] = add_74719 == 32'h0000_0005 ? array_update_75380 : array_update_75369[5];
  assign array_update_75382[6] = add_74719 == 32'h0000_0006 ? array_update_75380 : array_update_75369[6];
  assign array_update_75382[7] = add_74719 == 32'h0000_0007 ? array_update_75380 : array_update_75369[7];
  assign array_update_75382[8] = add_74719 == 32'h0000_0008 ? array_update_75380 : array_update_75369[8];
  assign array_update_75382[9] = add_74719 == 32'h0000_0009 ? array_update_75380 : array_update_75369[9];
  assign array_index_75384 = array_update_72021[add_75381 > 32'h0000_0009 ? 4'h9 : add_75381[3:0]];
  assign array_index_75385 = array_update_75382[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_75389 = smul32b_32b_x_32b(array_index_74726[add_75381 > 32'h0000_0009 ? 4'h9 : add_75381[3:0]], array_index_75384[add_75262 > 32'h0000_0009 ? 4'h9 : add_75262[3:0]]);
  assign add_75391 = array_index_75385[add_75262 > 32'h0000_0009 ? 4'h9 : add_75262[3:0]] + smul_75389;
  assign array_update_75392[0] = add_75262 == 32'h0000_0000 ? add_75391 : array_index_75385[0];
  assign array_update_75392[1] = add_75262 == 32'h0000_0001 ? add_75391 : array_index_75385[1];
  assign array_update_75392[2] = add_75262 == 32'h0000_0002 ? add_75391 : array_index_75385[2];
  assign array_update_75392[3] = add_75262 == 32'h0000_0003 ? add_75391 : array_index_75385[3];
  assign array_update_75392[4] = add_75262 == 32'h0000_0004 ? add_75391 : array_index_75385[4];
  assign array_update_75392[5] = add_75262 == 32'h0000_0005 ? add_75391 : array_index_75385[5];
  assign array_update_75392[6] = add_75262 == 32'h0000_0006 ? add_75391 : array_index_75385[6];
  assign array_update_75392[7] = add_75262 == 32'h0000_0007 ? add_75391 : array_index_75385[7];
  assign array_update_75392[8] = add_75262 == 32'h0000_0008 ? add_75391 : array_index_75385[8];
  assign array_update_75392[9] = add_75262 == 32'h0000_0009 ? add_75391 : array_index_75385[9];
  assign array_update_75393[0] = add_74719 == 32'h0000_0000 ? array_update_75392 : array_update_75382[0];
  assign array_update_75393[1] = add_74719 == 32'h0000_0001 ? array_update_75392 : array_update_75382[1];
  assign array_update_75393[2] = add_74719 == 32'h0000_0002 ? array_update_75392 : array_update_75382[2];
  assign array_update_75393[3] = add_74719 == 32'h0000_0003 ? array_update_75392 : array_update_75382[3];
  assign array_update_75393[4] = add_74719 == 32'h0000_0004 ? array_update_75392 : array_update_75382[4];
  assign array_update_75393[5] = add_74719 == 32'h0000_0005 ? array_update_75392 : array_update_75382[5];
  assign array_update_75393[6] = add_74719 == 32'h0000_0006 ? array_update_75392 : array_update_75382[6];
  assign array_update_75393[7] = add_74719 == 32'h0000_0007 ? array_update_75392 : array_update_75382[7];
  assign array_update_75393[8] = add_74719 == 32'h0000_0008 ? array_update_75392 : array_update_75382[8];
  assign array_update_75393[9] = add_74719 == 32'h0000_0009 ? array_update_75392 : array_update_75382[9];
  assign array_index_75395 = array_update_75393[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign add_75397 = add_75262 + 32'h0000_0001;
  assign array_update_75398[0] = add_75397 == 32'h0000_0000 ? 32'h0000_0000 : array_index_75395[0];
  assign array_update_75398[1] = add_75397 == 32'h0000_0001 ? 32'h0000_0000 : array_index_75395[1];
  assign array_update_75398[2] = add_75397 == 32'h0000_0002 ? 32'h0000_0000 : array_index_75395[2];
  assign array_update_75398[3] = add_75397 == 32'h0000_0003 ? 32'h0000_0000 : array_index_75395[3];
  assign array_update_75398[4] = add_75397 == 32'h0000_0004 ? 32'h0000_0000 : array_index_75395[4];
  assign array_update_75398[5] = add_75397 == 32'h0000_0005 ? 32'h0000_0000 : array_index_75395[5];
  assign array_update_75398[6] = add_75397 == 32'h0000_0006 ? 32'h0000_0000 : array_index_75395[6];
  assign array_update_75398[7] = add_75397 == 32'h0000_0007 ? 32'h0000_0000 : array_index_75395[7];
  assign array_update_75398[8] = add_75397 == 32'h0000_0008 ? 32'h0000_0000 : array_index_75395[8];
  assign array_update_75398[9] = add_75397 == 32'h0000_0009 ? 32'h0000_0000 : array_index_75395[9];
  assign literal_75399 = 32'h0000_0000;
  assign array_update_75400[0] = add_74719 == 32'h0000_0000 ? array_update_75398 : array_update_75393[0];
  assign array_update_75400[1] = add_74719 == 32'h0000_0001 ? array_update_75398 : array_update_75393[1];
  assign array_update_75400[2] = add_74719 == 32'h0000_0002 ? array_update_75398 : array_update_75393[2];
  assign array_update_75400[3] = add_74719 == 32'h0000_0003 ? array_update_75398 : array_update_75393[3];
  assign array_update_75400[4] = add_74719 == 32'h0000_0004 ? array_update_75398 : array_update_75393[4];
  assign array_update_75400[5] = add_74719 == 32'h0000_0005 ? array_update_75398 : array_update_75393[5];
  assign array_update_75400[6] = add_74719 == 32'h0000_0006 ? array_update_75398 : array_update_75393[6];
  assign array_update_75400[7] = add_74719 == 32'h0000_0007 ? array_update_75398 : array_update_75393[7];
  assign array_update_75400[8] = add_74719 == 32'h0000_0008 ? array_update_75398 : array_update_75393[8];
  assign array_update_75400[9] = add_74719 == 32'h0000_0009 ? array_update_75398 : array_update_75393[9];
  assign array_index_75402 = array_update_72021[literal_75399 > 32'h0000_0009 ? 4'h9 : literal_75399[3:0]];
  assign array_index_75403 = array_update_75400[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_75407 = smul32b_32b_x_32b(array_index_74726[literal_75399 > 32'h0000_0009 ? 4'h9 : literal_75399[3:0]], array_index_75402[add_75397 > 32'h0000_0009 ? 4'h9 : add_75397[3:0]]);
  assign add_75409 = array_index_75403[add_75397 > 32'h0000_0009 ? 4'h9 : add_75397[3:0]] + smul_75407;
  assign array_update_75411[0] = add_75397 == 32'h0000_0000 ? add_75409 : array_index_75403[0];
  assign array_update_75411[1] = add_75397 == 32'h0000_0001 ? add_75409 : array_index_75403[1];
  assign array_update_75411[2] = add_75397 == 32'h0000_0002 ? add_75409 : array_index_75403[2];
  assign array_update_75411[3] = add_75397 == 32'h0000_0003 ? add_75409 : array_index_75403[3];
  assign array_update_75411[4] = add_75397 == 32'h0000_0004 ? add_75409 : array_index_75403[4];
  assign array_update_75411[5] = add_75397 == 32'h0000_0005 ? add_75409 : array_index_75403[5];
  assign array_update_75411[6] = add_75397 == 32'h0000_0006 ? add_75409 : array_index_75403[6];
  assign array_update_75411[7] = add_75397 == 32'h0000_0007 ? add_75409 : array_index_75403[7];
  assign array_update_75411[8] = add_75397 == 32'h0000_0008 ? add_75409 : array_index_75403[8];
  assign array_update_75411[9] = add_75397 == 32'h0000_0009 ? add_75409 : array_index_75403[9];
  assign add_75412 = literal_75399 + 32'h0000_0001;
  assign array_update_75413[0] = add_74719 == 32'h0000_0000 ? array_update_75411 : array_update_75400[0];
  assign array_update_75413[1] = add_74719 == 32'h0000_0001 ? array_update_75411 : array_update_75400[1];
  assign array_update_75413[2] = add_74719 == 32'h0000_0002 ? array_update_75411 : array_update_75400[2];
  assign array_update_75413[3] = add_74719 == 32'h0000_0003 ? array_update_75411 : array_update_75400[3];
  assign array_update_75413[4] = add_74719 == 32'h0000_0004 ? array_update_75411 : array_update_75400[4];
  assign array_update_75413[5] = add_74719 == 32'h0000_0005 ? array_update_75411 : array_update_75400[5];
  assign array_update_75413[6] = add_74719 == 32'h0000_0006 ? array_update_75411 : array_update_75400[6];
  assign array_update_75413[7] = add_74719 == 32'h0000_0007 ? array_update_75411 : array_update_75400[7];
  assign array_update_75413[8] = add_74719 == 32'h0000_0008 ? array_update_75411 : array_update_75400[8];
  assign array_update_75413[9] = add_74719 == 32'h0000_0009 ? array_update_75411 : array_update_75400[9];
  assign array_index_75415 = array_update_72021[add_75412 > 32'h0000_0009 ? 4'h9 : add_75412[3:0]];
  assign array_index_75416 = array_update_75413[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_75420 = smul32b_32b_x_32b(array_index_74726[add_75412 > 32'h0000_0009 ? 4'h9 : add_75412[3:0]], array_index_75415[add_75397 > 32'h0000_0009 ? 4'h9 : add_75397[3:0]]);
  assign add_75422 = array_index_75416[add_75397 > 32'h0000_0009 ? 4'h9 : add_75397[3:0]] + smul_75420;
  assign array_update_75424[0] = add_75397 == 32'h0000_0000 ? add_75422 : array_index_75416[0];
  assign array_update_75424[1] = add_75397 == 32'h0000_0001 ? add_75422 : array_index_75416[1];
  assign array_update_75424[2] = add_75397 == 32'h0000_0002 ? add_75422 : array_index_75416[2];
  assign array_update_75424[3] = add_75397 == 32'h0000_0003 ? add_75422 : array_index_75416[3];
  assign array_update_75424[4] = add_75397 == 32'h0000_0004 ? add_75422 : array_index_75416[4];
  assign array_update_75424[5] = add_75397 == 32'h0000_0005 ? add_75422 : array_index_75416[5];
  assign array_update_75424[6] = add_75397 == 32'h0000_0006 ? add_75422 : array_index_75416[6];
  assign array_update_75424[7] = add_75397 == 32'h0000_0007 ? add_75422 : array_index_75416[7];
  assign array_update_75424[8] = add_75397 == 32'h0000_0008 ? add_75422 : array_index_75416[8];
  assign array_update_75424[9] = add_75397 == 32'h0000_0009 ? add_75422 : array_index_75416[9];
  assign add_75425 = add_75412 + 32'h0000_0001;
  assign array_update_75426[0] = add_74719 == 32'h0000_0000 ? array_update_75424 : array_update_75413[0];
  assign array_update_75426[1] = add_74719 == 32'h0000_0001 ? array_update_75424 : array_update_75413[1];
  assign array_update_75426[2] = add_74719 == 32'h0000_0002 ? array_update_75424 : array_update_75413[2];
  assign array_update_75426[3] = add_74719 == 32'h0000_0003 ? array_update_75424 : array_update_75413[3];
  assign array_update_75426[4] = add_74719 == 32'h0000_0004 ? array_update_75424 : array_update_75413[4];
  assign array_update_75426[5] = add_74719 == 32'h0000_0005 ? array_update_75424 : array_update_75413[5];
  assign array_update_75426[6] = add_74719 == 32'h0000_0006 ? array_update_75424 : array_update_75413[6];
  assign array_update_75426[7] = add_74719 == 32'h0000_0007 ? array_update_75424 : array_update_75413[7];
  assign array_update_75426[8] = add_74719 == 32'h0000_0008 ? array_update_75424 : array_update_75413[8];
  assign array_update_75426[9] = add_74719 == 32'h0000_0009 ? array_update_75424 : array_update_75413[9];
  assign array_index_75428 = array_update_72021[add_75425 > 32'h0000_0009 ? 4'h9 : add_75425[3:0]];
  assign array_index_75429 = array_update_75426[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_75433 = smul32b_32b_x_32b(array_index_74726[add_75425 > 32'h0000_0009 ? 4'h9 : add_75425[3:0]], array_index_75428[add_75397 > 32'h0000_0009 ? 4'h9 : add_75397[3:0]]);
  assign add_75435 = array_index_75429[add_75397 > 32'h0000_0009 ? 4'h9 : add_75397[3:0]] + smul_75433;
  assign array_update_75437[0] = add_75397 == 32'h0000_0000 ? add_75435 : array_index_75429[0];
  assign array_update_75437[1] = add_75397 == 32'h0000_0001 ? add_75435 : array_index_75429[1];
  assign array_update_75437[2] = add_75397 == 32'h0000_0002 ? add_75435 : array_index_75429[2];
  assign array_update_75437[3] = add_75397 == 32'h0000_0003 ? add_75435 : array_index_75429[3];
  assign array_update_75437[4] = add_75397 == 32'h0000_0004 ? add_75435 : array_index_75429[4];
  assign array_update_75437[5] = add_75397 == 32'h0000_0005 ? add_75435 : array_index_75429[5];
  assign array_update_75437[6] = add_75397 == 32'h0000_0006 ? add_75435 : array_index_75429[6];
  assign array_update_75437[7] = add_75397 == 32'h0000_0007 ? add_75435 : array_index_75429[7];
  assign array_update_75437[8] = add_75397 == 32'h0000_0008 ? add_75435 : array_index_75429[8];
  assign array_update_75437[9] = add_75397 == 32'h0000_0009 ? add_75435 : array_index_75429[9];
  assign add_75438 = add_75425 + 32'h0000_0001;
  assign array_update_75439[0] = add_74719 == 32'h0000_0000 ? array_update_75437 : array_update_75426[0];
  assign array_update_75439[1] = add_74719 == 32'h0000_0001 ? array_update_75437 : array_update_75426[1];
  assign array_update_75439[2] = add_74719 == 32'h0000_0002 ? array_update_75437 : array_update_75426[2];
  assign array_update_75439[3] = add_74719 == 32'h0000_0003 ? array_update_75437 : array_update_75426[3];
  assign array_update_75439[4] = add_74719 == 32'h0000_0004 ? array_update_75437 : array_update_75426[4];
  assign array_update_75439[5] = add_74719 == 32'h0000_0005 ? array_update_75437 : array_update_75426[5];
  assign array_update_75439[6] = add_74719 == 32'h0000_0006 ? array_update_75437 : array_update_75426[6];
  assign array_update_75439[7] = add_74719 == 32'h0000_0007 ? array_update_75437 : array_update_75426[7];
  assign array_update_75439[8] = add_74719 == 32'h0000_0008 ? array_update_75437 : array_update_75426[8];
  assign array_update_75439[9] = add_74719 == 32'h0000_0009 ? array_update_75437 : array_update_75426[9];
  assign array_index_75441 = array_update_72021[add_75438 > 32'h0000_0009 ? 4'h9 : add_75438[3:0]];
  assign array_index_75442 = array_update_75439[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_75446 = smul32b_32b_x_32b(array_index_74726[add_75438 > 32'h0000_0009 ? 4'h9 : add_75438[3:0]], array_index_75441[add_75397 > 32'h0000_0009 ? 4'h9 : add_75397[3:0]]);
  assign add_75448 = array_index_75442[add_75397 > 32'h0000_0009 ? 4'h9 : add_75397[3:0]] + smul_75446;
  assign array_update_75450[0] = add_75397 == 32'h0000_0000 ? add_75448 : array_index_75442[0];
  assign array_update_75450[1] = add_75397 == 32'h0000_0001 ? add_75448 : array_index_75442[1];
  assign array_update_75450[2] = add_75397 == 32'h0000_0002 ? add_75448 : array_index_75442[2];
  assign array_update_75450[3] = add_75397 == 32'h0000_0003 ? add_75448 : array_index_75442[3];
  assign array_update_75450[4] = add_75397 == 32'h0000_0004 ? add_75448 : array_index_75442[4];
  assign array_update_75450[5] = add_75397 == 32'h0000_0005 ? add_75448 : array_index_75442[5];
  assign array_update_75450[6] = add_75397 == 32'h0000_0006 ? add_75448 : array_index_75442[6];
  assign array_update_75450[7] = add_75397 == 32'h0000_0007 ? add_75448 : array_index_75442[7];
  assign array_update_75450[8] = add_75397 == 32'h0000_0008 ? add_75448 : array_index_75442[8];
  assign array_update_75450[9] = add_75397 == 32'h0000_0009 ? add_75448 : array_index_75442[9];
  assign add_75451 = add_75438 + 32'h0000_0001;
  assign array_update_75452[0] = add_74719 == 32'h0000_0000 ? array_update_75450 : array_update_75439[0];
  assign array_update_75452[1] = add_74719 == 32'h0000_0001 ? array_update_75450 : array_update_75439[1];
  assign array_update_75452[2] = add_74719 == 32'h0000_0002 ? array_update_75450 : array_update_75439[2];
  assign array_update_75452[3] = add_74719 == 32'h0000_0003 ? array_update_75450 : array_update_75439[3];
  assign array_update_75452[4] = add_74719 == 32'h0000_0004 ? array_update_75450 : array_update_75439[4];
  assign array_update_75452[5] = add_74719 == 32'h0000_0005 ? array_update_75450 : array_update_75439[5];
  assign array_update_75452[6] = add_74719 == 32'h0000_0006 ? array_update_75450 : array_update_75439[6];
  assign array_update_75452[7] = add_74719 == 32'h0000_0007 ? array_update_75450 : array_update_75439[7];
  assign array_update_75452[8] = add_74719 == 32'h0000_0008 ? array_update_75450 : array_update_75439[8];
  assign array_update_75452[9] = add_74719 == 32'h0000_0009 ? array_update_75450 : array_update_75439[9];
  assign array_index_75454 = array_update_72021[add_75451 > 32'h0000_0009 ? 4'h9 : add_75451[3:0]];
  assign array_index_75455 = array_update_75452[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_75459 = smul32b_32b_x_32b(array_index_74726[add_75451 > 32'h0000_0009 ? 4'h9 : add_75451[3:0]], array_index_75454[add_75397 > 32'h0000_0009 ? 4'h9 : add_75397[3:0]]);
  assign add_75461 = array_index_75455[add_75397 > 32'h0000_0009 ? 4'h9 : add_75397[3:0]] + smul_75459;
  assign array_update_75463[0] = add_75397 == 32'h0000_0000 ? add_75461 : array_index_75455[0];
  assign array_update_75463[1] = add_75397 == 32'h0000_0001 ? add_75461 : array_index_75455[1];
  assign array_update_75463[2] = add_75397 == 32'h0000_0002 ? add_75461 : array_index_75455[2];
  assign array_update_75463[3] = add_75397 == 32'h0000_0003 ? add_75461 : array_index_75455[3];
  assign array_update_75463[4] = add_75397 == 32'h0000_0004 ? add_75461 : array_index_75455[4];
  assign array_update_75463[5] = add_75397 == 32'h0000_0005 ? add_75461 : array_index_75455[5];
  assign array_update_75463[6] = add_75397 == 32'h0000_0006 ? add_75461 : array_index_75455[6];
  assign array_update_75463[7] = add_75397 == 32'h0000_0007 ? add_75461 : array_index_75455[7];
  assign array_update_75463[8] = add_75397 == 32'h0000_0008 ? add_75461 : array_index_75455[8];
  assign array_update_75463[9] = add_75397 == 32'h0000_0009 ? add_75461 : array_index_75455[9];
  assign add_75464 = add_75451 + 32'h0000_0001;
  assign array_update_75465[0] = add_74719 == 32'h0000_0000 ? array_update_75463 : array_update_75452[0];
  assign array_update_75465[1] = add_74719 == 32'h0000_0001 ? array_update_75463 : array_update_75452[1];
  assign array_update_75465[2] = add_74719 == 32'h0000_0002 ? array_update_75463 : array_update_75452[2];
  assign array_update_75465[3] = add_74719 == 32'h0000_0003 ? array_update_75463 : array_update_75452[3];
  assign array_update_75465[4] = add_74719 == 32'h0000_0004 ? array_update_75463 : array_update_75452[4];
  assign array_update_75465[5] = add_74719 == 32'h0000_0005 ? array_update_75463 : array_update_75452[5];
  assign array_update_75465[6] = add_74719 == 32'h0000_0006 ? array_update_75463 : array_update_75452[6];
  assign array_update_75465[7] = add_74719 == 32'h0000_0007 ? array_update_75463 : array_update_75452[7];
  assign array_update_75465[8] = add_74719 == 32'h0000_0008 ? array_update_75463 : array_update_75452[8];
  assign array_update_75465[9] = add_74719 == 32'h0000_0009 ? array_update_75463 : array_update_75452[9];
  assign array_index_75467 = array_update_72021[add_75464 > 32'h0000_0009 ? 4'h9 : add_75464[3:0]];
  assign array_index_75468 = array_update_75465[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_75472 = smul32b_32b_x_32b(array_index_74726[add_75464 > 32'h0000_0009 ? 4'h9 : add_75464[3:0]], array_index_75467[add_75397 > 32'h0000_0009 ? 4'h9 : add_75397[3:0]]);
  assign add_75474 = array_index_75468[add_75397 > 32'h0000_0009 ? 4'h9 : add_75397[3:0]] + smul_75472;
  assign array_update_75476[0] = add_75397 == 32'h0000_0000 ? add_75474 : array_index_75468[0];
  assign array_update_75476[1] = add_75397 == 32'h0000_0001 ? add_75474 : array_index_75468[1];
  assign array_update_75476[2] = add_75397 == 32'h0000_0002 ? add_75474 : array_index_75468[2];
  assign array_update_75476[3] = add_75397 == 32'h0000_0003 ? add_75474 : array_index_75468[3];
  assign array_update_75476[4] = add_75397 == 32'h0000_0004 ? add_75474 : array_index_75468[4];
  assign array_update_75476[5] = add_75397 == 32'h0000_0005 ? add_75474 : array_index_75468[5];
  assign array_update_75476[6] = add_75397 == 32'h0000_0006 ? add_75474 : array_index_75468[6];
  assign array_update_75476[7] = add_75397 == 32'h0000_0007 ? add_75474 : array_index_75468[7];
  assign array_update_75476[8] = add_75397 == 32'h0000_0008 ? add_75474 : array_index_75468[8];
  assign array_update_75476[9] = add_75397 == 32'h0000_0009 ? add_75474 : array_index_75468[9];
  assign add_75477 = add_75464 + 32'h0000_0001;
  assign array_update_75478[0] = add_74719 == 32'h0000_0000 ? array_update_75476 : array_update_75465[0];
  assign array_update_75478[1] = add_74719 == 32'h0000_0001 ? array_update_75476 : array_update_75465[1];
  assign array_update_75478[2] = add_74719 == 32'h0000_0002 ? array_update_75476 : array_update_75465[2];
  assign array_update_75478[3] = add_74719 == 32'h0000_0003 ? array_update_75476 : array_update_75465[3];
  assign array_update_75478[4] = add_74719 == 32'h0000_0004 ? array_update_75476 : array_update_75465[4];
  assign array_update_75478[5] = add_74719 == 32'h0000_0005 ? array_update_75476 : array_update_75465[5];
  assign array_update_75478[6] = add_74719 == 32'h0000_0006 ? array_update_75476 : array_update_75465[6];
  assign array_update_75478[7] = add_74719 == 32'h0000_0007 ? array_update_75476 : array_update_75465[7];
  assign array_update_75478[8] = add_74719 == 32'h0000_0008 ? array_update_75476 : array_update_75465[8];
  assign array_update_75478[9] = add_74719 == 32'h0000_0009 ? array_update_75476 : array_update_75465[9];
  assign array_index_75480 = array_update_72021[add_75477 > 32'h0000_0009 ? 4'h9 : add_75477[3:0]];
  assign array_index_75481 = array_update_75478[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_75485 = smul32b_32b_x_32b(array_index_74726[add_75477 > 32'h0000_0009 ? 4'h9 : add_75477[3:0]], array_index_75480[add_75397 > 32'h0000_0009 ? 4'h9 : add_75397[3:0]]);
  assign add_75487 = array_index_75481[add_75397 > 32'h0000_0009 ? 4'h9 : add_75397[3:0]] + smul_75485;
  assign array_update_75489[0] = add_75397 == 32'h0000_0000 ? add_75487 : array_index_75481[0];
  assign array_update_75489[1] = add_75397 == 32'h0000_0001 ? add_75487 : array_index_75481[1];
  assign array_update_75489[2] = add_75397 == 32'h0000_0002 ? add_75487 : array_index_75481[2];
  assign array_update_75489[3] = add_75397 == 32'h0000_0003 ? add_75487 : array_index_75481[3];
  assign array_update_75489[4] = add_75397 == 32'h0000_0004 ? add_75487 : array_index_75481[4];
  assign array_update_75489[5] = add_75397 == 32'h0000_0005 ? add_75487 : array_index_75481[5];
  assign array_update_75489[6] = add_75397 == 32'h0000_0006 ? add_75487 : array_index_75481[6];
  assign array_update_75489[7] = add_75397 == 32'h0000_0007 ? add_75487 : array_index_75481[7];
  assign array_update_75489[8] = add_75397 == 32'h0000_0008 ? add_75487 : array_index_75481[8];
  assign array_update_75489[9] = add_75397 == 32'h0000_0009 ? add_75487 : array_index_75481[9];
  assign add_75490 = add_75477 + 32'h0000_0001;
  assign array_update_75491[0] = add_74719 == 32'h0000_0000 ? array_update_75489 : array_update_75478[0];
  assign array_update_75491[1] = add_74719 == 32'h0000_0001 ? array_update_75489 : array_update_75478[1];
  assign array_update_75491[2] = add_74719 == 32'h0000_0002 ? array_update_75489 : array_update_75478[2];
  assign array_update_75491[3] = add_74719 == 32'h0000_0003 ? array_update_75489 : array_update_75478[3];
  assign array_update_75491[4] = add_74719 == 32'h0000_0004 ? array_update_75489 : array_update_75478[4];
  assign array_update_75491[5] = add_74719 == 32'h0000_0005 ? array_update_75489 : array_update_75478[5];
  assign array_update_75491[6] = add_74719 == 32'h0000_0006 ? array_update_75489 : array_update_75478[6];
  assign array_update_75491[7] = add_74719 == 32'h0000_0007 ? array_update_75489 : array_update_75478[7];
  assign array_update_75491[8] = add_74719 == 32'h0000_0008 ? array_update_75489 : array_update_75478[8];
  assign array_update_75491[9] = add_74719 == 32'h0000_0009 ? array_update_75489 : array_update_75478[9];
  assign array_index_75493 = array_update_72021[add_75490 > 32'h0000_0009 ? 4'h9 : add_75490[3:0]];
  assign array_index_75494 = array_update_75491[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_75498 = smul32b_32b_x_32b(array_index_74726[add_75490 > 32'h0000_0009 ? 4'h9 : add_75490[3:0]], array_index_75493[add_75397 > 32'h0000_0009 ? 4'h9 : add_75397[3:0]]);
  assign add_75500 = array_index_75494[add_75397 > 32'h0000_0009 ? 4'h9 : add_75397[3:0]] + smul_75498;
  assign array_update_75502[0] = add_75397 == 32'h0000_0000 ? add_75500 : array_index_75494[0];
  assign array_update_75502[1] = add_75397 == 32'h0000_0001 ? add_75500 : array_index_75494[1];
  assign array_update_75502[2] = add_75397 == 32'h0000_0002 ? add_75500 : array_index_75494[2];
  assign array_update_75502[3] = add_75397 == 32'h0000_0003 ? add_75500 : array_index_75494[3];
  assign array_update_75502[4] = add_75397 == 32'h0000_0004 ? add_75500 : array_index_75494[4];
  assign array_update_75502[5] = add_75397 == 32'h0000_0005 ? add_75500 : array_index_75494[5];
  assign array_update_75502[6] = add_75397 == 32'h0000_0006 ? add_75500 : array_index_75494[6];
  assign array_update_75502[7] = add_75397 == 32'h0000_0007 ? add_75500 : array_index_75494[7];
  assign array_update_75502[8] = add_75397 == 32'h0000_0008 ? add_75500 : array_index_75494[8];
  assign array_update_75502[9] = add_75397 == 32'h0000_0009 ? add_75500 : array_index_75494[9];
  assign add_75503 = add_75490 + 32'h0000_0001;
  assign array_update_75504[0] = add_74719 == 32'h0000_0000 ? array_update_75502 : array_update_75491[0];
  assign array_update_75504[1] = add_74719 == 32'h0000_0001 ? array_update_75502 : array_update_75491[1];
  assign array_update_75504[2] = add_74719 == 32'h0000_0002 ? array_update_75502 : array_update_75491[2];
  assign array_update_75504[3] = add_74719 == 32'h0000_0003 ? array_update_75502 : array_update_75491[3];
  assign array_update_75504[4] = add_74719 == 32'h0000_0004 ? array_update_75502 : array_update_75491[4];
  assign array_update_75504[5] = add_74719 == 32'h0000_0005 ? array_update_75502 : array_update_75491[5];
  assign array_update_75504[6] = add_74719 == 32'h0000_0006 ? array_update_75502 : array_update_75491[6];
  assign array_update_75504[7] = add_74719 == 32'h0000_0007 ? array_update_75502 : array_update_75491[7];
  assign array_update_75504[8] = add_74719 == 32'h0000_0008 ? array_update_75502 : array_update_75491[8];
  assign array_update_75504[9] = add_74719 == 32'h0000_0009 ? array_update_75502 : array_update_75491[9];
  assign array_index_75506 = array_update_72021[add_75503 > 32'h0000_0009 ? 4'h9 : add_75503[3:0]];
  assign array_index_75507 = array_update_75504[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_75511 = smul32b_32b_x_32b(array_index_74726[add_75503 > 32'h0000_0009 ? 4'h9 : add_75503[3:0]], array_index_75506[add_75397 > 32'h0000_0009 ? 4'h9 : add_75397[3:0]]);
  assign add_75513 = array_index_75507[add_75397 > 32'h0000_0009 ? 4'h9 : add_75397[3:0]] + smul_75511;
  assign array_update_75515[0] = add_75397 == 32'h0000_0000 ? add_75513 : array_index_75507[0];
  assign array_update_75515[1] = add_75397 == 32'h0000_0001 ? add_75513 : array_index_75507[1];
  assign array_update_75515[2] = add_75397 == 32'h0000_0002 ? add_75513 : array_index_75507[2];
  assign array_update_75515[3] = add_75397 == 32'h0000_0003 ? add_75513 : array_index_75507[3];
  assign array_update_75515[4] = add_75397 == 32'h0000_0004 ? add_75513 : array_index_75507[4];
  assign array_update_75515[5] = add_75397 == 32'h0000_0005 ? add_75513 : array_index_75507[5];
  assign array_update_75515[6] = add_75397 == 32'h0000_0006 ? add_75513 : array_index_75507[6];
  assign array_update_75515[7] = add_75397 == 32'h0000_0007 ? add_75513 : array_index_75507[7];
  assign array_update_75515[8] = add_75397 == 32'h0000_0008 ? add_75513 : array_index_75507[8];
  assign array_update_75515[9] = add_75397 == 32'h0000_0009 ? add_75513 : array_index_75507[9];
  assign add_75516 = add_75503 + 32'h0000_0001;
  assign array_update_75517[0] = add_74719 == 32'h0000_0000 ? array_update_75515 : array_update_75504[0];
  assign array_update_75517[1] = add_74719 == 32'h0000_0001 ? array_update_75515 : array_update_75504[1];
  assign array_update_75517[2] = add_74719 == 32'h0000_0002 ? array_update_75515 : array_update_75504[2];
  assign array_update_75517[3] = add_74719 == 32'h0000_0003 ? array_update_75515 : array_update_75504[3];
  assign array_update_75517[4] = add_74719 == 32'h0000_0004 ? array_update_75515 : array_update_75504[4];
  assign array_update_75517[5] = add_74719 == 32'h0000_0005 ? array_update_75515 : array_update_75504[5];
  assign array_update_75517[6] = add_74719 == 32'h0000_0006 ? array_update_75515 : array_update_75504[6];
  assign array_update_75517[7] = add_74719 == 32'h0000_0007 ? array_update_75515 : array_update_75504[7];
  assign array_update_75517[8] = add_74719 == 32'h0000_0008 ? array_update_75515 : array_update_75504[8];
  assign array_update_75517[9] = add_74719 == 32'h0000_0009 ? array_update_75515 : array_update_75504[9];
  assign array_index_75519 = array_update_72021[add_75516 > 32'h0000_0009 ? 4'h9 : add_75516[3:0]];
  assign array_index_75520 = array_update_75517[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_75524 = smul32b_32b_x_32b(array_index_74726[add_75516 > 32'h0000_0009 ? 4'h9 : add_75516[3:0]], array_index_75519[add_75397 > 32'h0000_0009 ? 4'h9 : add_75397[3:0]]);
  assign add_75526 = array_index_75520[add_75397 > 32'h0000_0009 ? 4'h9 : add_75397[3:0]] + smul_75524;
  assign array_update_75527[0] = add_75397 == 32'h0000_0000 ? add_75526 : array_index_75520[0];
  assign array_update_75527[1] = add_75397 == 32'h0000_0001 ? add_75526 : array_index_75520[1];
  assign array_update_75527[2] = add_75397 == 32'h0000_0002 ? add_75526 : array_index_75520[2];
  assign array_update_75527[3] = add_75397 == 32'h0000_0003 ? add_75526 : array_index_75520[3];
  assign array_update_75527[4] = add_75397 == 32'h0000_0004 ? add_75526 : array_index_75520[4];
  assign array_update_75527[5] = add_75397 == 32'h0000_0005 ? add_75526 : array_index_75520[5];
  assign array_update_75527[6] = add_75397 == 32'h0000_0006 ? add_75526 : array_index_75520[6];
  assign array_update_75527[7] = add_75397 == 32'h0000_0007 ? add_75526 : array_index_75520[7];
  assign array_update_75527[8] = add_75397 == 32'h0000_0008 ? add_75526 : array_index_75520[8];
  assign array_update_75527[9] = add_75397 == 32'h0000_0009 ? add_75526 : array_index_75520[9];
  assign array_update_75528[0] = add_74719 == 32'h0000_0000 ? array_update_75527 : array_update_75517[0];
  assign array_update_75528[1] = add_74719 == 32'h0000_0001 ? array_update_75527 : array_update_75517[1];
  assign array_update_75528[2] = add_74719 == 32'h0000_0002 ? array_update_75527 : array_update_75517[2];
  assign array_update_75528[3] = add_74719 == 32'h0000_0003 ? array_update_75527 : array_update_75517[3];
  assign array_update_75528[4] = add_74719 == 32'h0000_0004 ? array_update_75527 : array_update_75517[4];
  assign array_update_75528[5] = add_74719 == 32'h0000_0005 ? array_update_75527 : array_update_75517[5];
  assign array_update_75528[6] = add_74719 == 32'h0000_0006 ? array_update_75527 : array_update_75517[6];
  assign array_update_75528[7] = add_74719 == 32'h0000_0007 ? array_update_75527 : array_update_75517[7];
  assign array_update_75528[8] = add_74719 == 32'h0000_0008 ? array_update_75527 : array_update_75517[8];
  assign array_update_75528[9] = add_74719 == 32'h0000_0009 ? array_update_75527 : array_update_75517[9];
  assign array_index_75530 = array_update_75528[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign add_75532 = add_75397 + 32'h0000_0001;
  assign array_update_75533[0] = add_75532 == 32'h0000_0000 ? 32'h0000_0000 : array_index_75530[0];
  assign array_update_75533[1] = add_75532 == 32'h0000_0001 ? 32'h0000_0000 : array_index_75530[1];
  assign array_update_75533[2] = add_75532 == 32'h0000_0002 ? 32'h0000_0000 : array_index_75530[2];
  assign array_update_75533[3] = add_75532 == 32'h0000_0003 ? 32'h0000_0000 : array_index_75530[3];
  assign array_update_75533[4] = add_75532 == 32'h0000_0004 ? 32'h0000_0000 : array_index_75530[4];
  assign array_update_75533[5] = add_75532 == 32'h0000_0005 ? 32'h0000_0000 : array_index_75530[5];
  assign array_update_75533[6] = add_75532 == 32'h0000_0006 ? 32'h0000_0000 : array_index_75530[6];
  assign array_update_75533[7] = add_75532 == 32'h0000_0007 ? 32'h0000_0000 : array_index_75530[7];
  assign array_update_75533[8] = add_75532 == 32'h0000_0008 ? 32'h0000_0000 : array_index_75530[8];
  assign array_update_75533[9] = add_75532 == 32'h0000_0009 ? 32'h0000_0000 : array_index_75530[9];
  assign literal_75534 = 32'h0000_0000;
  assign array_update_75535[0] = add_74719 == 32'h0000_0000 ? array_update_75533 : array_update_75528[0];
  assign array_update_75535[1] = add_74719 == 32'h0000_0001 ? array_update_75533 : array_update_75528[1];
  assign array_update_75535[2] = add_74719 == 32'h0000_0002 ? array_update_75533 : array_update_75528[2];
  assign array_update_75535[3] = add_74719 == 32'h0000_0003 ? array_update_75533 : array_update_75528[3];
  assign array_update_75535[4] = add_74719 == 32'h0000_0004 ? array_update_75533 : array_update_75528[4];
  assign array_update_75535[5] = add_74719 == 32'h0000_0005 ? array_update_75533 : array_update_75528[5];
  assign array_update_75535[6] = add_74719 == 32'h0000_0006 ? array_update_75533 : array_update_75528[6];
  assign array_update_75535[7] = add_74719 == 32'h0000_0007 ? array_update_75533 : array_update_75528[7];
  assign array_update_75535[8] = add_74719 == 32'h0000_0008 ? array_update_75533 : array_update_75528[8];
  assign array_update_75535[9] = add_74719 == 32'h0000_0009 ? array_update_75533 : array_update_75528[9];
  assign array_index_75537 = array_update_72021[literal_75534 > 32'h0000_0009 ? 4'h9 : literal_75534[3:0]];
  assign array_index_75538 = array_update_75535[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_75542 = smul32b_32b_x_32b(array_index_74726[literal_75534 > 32'h0000_0009 ? 4'h9 : literal_75534[3:0]], array_index_75537[add_75532 > 32'h0000_0009 ? 4'h9 : add_75532[3:0]]);
  assign add_75544 = array_index_75538[add_75532 > 32'h0000_0009 ? 4'h9 : add_75532[3:0]] + smul_75542;
  assign array_update_75546[0] = add_75532 == 32'h0000_0000 ? add_75544 : array_index_75538[0];
  assign array_update_75546[1] = add_75532 == 32'h0000_0001 ? add_75544 : array_index_75538[1];
  assign array_update_75546[2] = add_75532 == 32'h0000_0002 ? add_75544 : array_index_75538[2];
  assign array_update_75546[3] = add_75532 == 32'h0000_0003 ? add_75544 : array_index_75538[3];
  assign array_update_75546[4] = add_75532 == 32'h0000_0004 ? add_75544 : array_index_75538[4];
  assign array_update_75546[5] = add_75532 == 32'h0000_0005 ? add_75544 : array_index_75538[5];
  assign array_update_75546[6] = add_75532 == 32'h0000_0006 ? add_75544 : array_index_75538[6];
  assign array_update_75546[7] = add_75532 == 32'h0000_0007 ? add_75544 : array_index_75538[7];
  assign array_update_75546[8] = add_75532 == 32'h0000_0008 ? add_75544 : array_index_75538[8];
  assign array_update_75546[9] = add_75532 == 32'h0000_0009 ? add_75544 : array_index_75538[9];
  assign add_75547 = literal_75534 + 32'h0000_0001;
  assign array_update_75548[0] = add_74719 == 32'h0000_0000 ? array_update_75546 : array_update_75535[0];
  assign array_update_75548[1] = add_74719 == 32'h0000_0001 ? array_update_75546 : array_update_75535[1];
  assign array_update_75548[2] = add_74719 == 32'h0000_0002 ? array_update_75546 : array_update_75535[2];
  assign array_update_75548[3] = add_74719 == 32'h0000_0003 ? array_update_75546 : array_update_75535[3];
  assign array_update_75548[4] = add_74719 == 32'h0000_0004 ? array_update_75546 : array_update_75535[4];
  assign array_update_75548[5] = add_74719 == 32'h0000_0005 ? array_update_75546 : array_update_75535[5];
  assign array_update_75548[6] = add_74719 == 32'h0000_0006 ? array_update_75546 : array_update_75535[6];
  assign array_update_75548[7] = add_74719 == 32'h0000_0007 ? array_update_75546 : array_update_75535[7];
  assign array_update_75548[8] = add_74719 == 32'h0000_0008 ? array_update_75546 : array_update_75535[8];
  assign array_update_75548[9] = add_74719 == 32'h0000_0009 ? array_update_75546 : array_update_75535[9];
  assign array_index_75550 = array_update_72021[add_75547 > 32'h0000_0009 ? 4'h9 : add_75547[3:0]];
  assign array_index_75551 = array_update_75548[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_75555 = smul32b_32b_x_32b(array_index_74726[add_75547 > 32'h0000_0009 ? 4'h9 : add_75547[3:0]], array_index_75550[add_75532 > 32'h0000_0009 ? 4'h9 : add_75532[3:0]]);
  assign add_75557 = array_index_75551[add_75532 > 32'h0000_0009 ? 4'h9 : add_75532[3:0]] + smul_75555;
  assign array_update_75559[0] = add_75532 == 32'h0000_0000 ? add_75557 : array_index_75551[0];
  assign array_update_75559[1] = add_75532 == 32'h0000_0001 ? add_75557 : array_index_75551[1];
  assign array_update_75559[2] = add_75532 == 32'h0000_0002 ? add_75557 : array_index_75551[2];
  assign array_update_75559[3] = add_75532 == 32'h0000_0003 ? add_75557 : array_index_75551[3];
  assign array_update_75559[4] = add_75532 == 32'h0000_0004 ? add_75557 : array_index_75551[4];
  assign array_update_75559[5] = add_75532 == 32'h0000_0005 ? add_75557 : array_index_75551[5];
  assign array_update_75559[6] = add_75532 == 32'h0000_0006 ? add_75557 : array_index_75551[6];
  assign array_update_75559[7] = add_75532 == 32'h0000_0007 ? add_75557 : array_index_75551[7];
  assign array_update_75559[8] = add_75532 == 32'h0000_0008 ? add_75557 : array_index_75551[8];
  assign array_update_75559[9] = add_75532 == 32'h0000_0009 ? add_75557 : array_index_75551[9];
  assign add_75560 = add_75547 + 32'h0000_0001;
  assign array_update_75561[0] = add_74719 == 32'h0000_0000 ? array_update_75559 : array_update_75548[0];
  assign array_update_75561[1] = add_74719 == 32'h0000_0001 ? array_update_75559 : array_update_75548[1];
  assign array_update_75561[2] = add_74719 == 32'h0000_0002 ? array_update_75559 : array_update_75548[2];
  assign array_update_75561[3] = add_74719 == 32'h0000_0003 ? array_update_75559 : array_update_75548[3];
  assign array_update_75561[4] = add_74719 == 32'h0000_0004 ? array_update_75559 : array_update_75548[4];
  assign array_update_75561[5] = add_74719 == 32'h0000_0005 ? array_update_75559 : array_update_75548[5];
  assign array_update_75561[6] = add_74719 == 32'h0000_0006 ? array_update_75559 : array_update_75548[6];
  assign array_update_75561[7] = add_74719 == 32'h0000_0007 ? array_update_75559 : array_update_75548[7];
  assign array_update_75561[8] = add_74719 == 32'h0000_0008 ? array_update_75559 : array_update_75548[8];
  assign array_update_75561[9] = add_74719 == 32'h0000_0009 ? array_update_75559 : array_update_75548[9];
  assign array_index_75563 = array_update_72021[add_75560 > 32'h0000_0009 ? 4'h9 : add_75560[3:0]];
  assign array_index_75564 = array_update_75561[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_75568 = smul32b_32b_x_32b(array_index_74726[add_75560 > 32'h0000_0009 ? 4'h9 : add_75560[3:0]], array_index_75563[add_75532 > 32'h0000_0009 ? 4'h9 : add_75532[3:0]]);
  assign add_75570 = array_index_75564[add_75532 > 32'h0000_0009 ? 4'h9 : add_75532[3:0]] + smul_75568;
  assign array_update_75572[0] = add_75532 == 32'h0000_0000 ? add_75570 : array_index_75564[0];
  assign array_update_75572[1] = add_75532 == 32'h0000_0001 ? add_75570 : array_index_75564[1];
  assign array_update_75572[2] = add_75532 == 32'h0000_0002 ? add_75570 : array_index_75564[2];
  assign array_update_75572[3] = add_75532 == 32'h0000_0003 ? add_75570 : array_index_75564[3];
  assign array_update_75572[4] = add_75532 == 32'h0000_0004 ? add_75570 : array_index_75564[4];
  assign array_update_75572[5] = add_75532 == 32'h0000_0005 ? add_75570 : array_index_75564[5];
  assign array_update_75572[6] = add_75532 == 32'h0000_0006 ? add_75570 : array_index_75564[6];
  assign array_update_75572[7] = add_75532 == 32'h0000_0007 ? add_75570 : array_index_75564[7];
  assign array_update_75572[8] = add_75532 == 32'h0000_0008 ? add_75570 : array_index_75564[8];
  assign array_update_75572[9] = add_75532 == 32'h0000_0009 ? add_75570 : array_index_75564[9];
  assign add_75573 = add_75560 + 32'h0000_0001;
  assign array_update_75574[0] = add_74719 == 32'h0000_0000 ? array_update_75572 : array_update_75561[0];
  assign array_update_75574[1] = add_74719 == 32'h0000_0001 ? array_update_75572 : array_update_75561[1];
  assign array_update_75574[2] = add_74719 == 32'h0000_0002 ? array_update_75572 : array_update_75561[2];
  assign array_update_75574[3] = add_74719 == 32'h0000_0003 ? array_update_75572 : array_update_75561[3];
  assign array_update_75574[4] = add_74719 == 32'h0000_0004 ? array_update_75572 : array_update_75561[4];
  assign array_update_75574[5] = add_74719 == 32'h0000_0005 ? array_update_75572 : array_update_75561[5];
  assign array_update_75574[6] = add_74719 == 32'h0000_0006 ? array_update_75572 : array_update_75561[6];
  assign array_update_75574[7] = add_74719 == 32'h0000_0007 ? array_update_75572 : array_update_75561[7];
  assign array_update_75574[8] = add_74719 == 32'h0000_0008 ? array_update_75572 : array_update_75561[8];
  assign array_update_75574[9] = add_74719 == 32'h0000_0009 ? array_update_75572 : array_update_75561[9];
  assign array_index_75576 = array_update_72021[add_75573 > 32'h0000_0009 ? 4'h9 : add_75573[3:0]];
  assign array_index_75577 = array_update_75574[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_75581 = smul32b_32b_x_32b(array_index_74726[add_75573 > 32'h0000_0009 ? 4'h9 : add_75573[3:0]], array_index_75576[add_75532 > 32'h0000_0009 ? 4'h9 : add_75532[3:0]]);
  assign add_75583 = array_index_75577[add_75532 > 32'h0000_0009 ? 4'h9 : add_75532[3:0]] + smul_75581;
  assign array_update_75585[0] = add_75532 == 32'h0000_0000 ? add_75583 : array_index_75577[0];
  assign array_update_75585[1] = add_75532 == 32'h0000_0001 ? add_75583 : array_index_75577[1];
  assign array_update_75585[2] = add_75532 == 32'h0000_0002 ? add_75583 : array_index_75577[2];
  assign array_update_75585[3] = add_75532 == 32'h0000_0003 ? add_75583 : array_index_75577[3];
  assign array_update_75585[4] = add_75532 == 32'h0000_0004 ? add_75583 : array_index_75577[4];
  assign array_update_75585[5] = add_75532 == 32'h0000_0005 ? add_75583 : array_index_75577[5];
  assign array_update_75585[6] = add_75532 == 32'h0000_0006 ? add_75583 : array_index_75577[6];
  assign array_update_75585[7] = add_75532 == 32'h0000_0007 ? add_75583 : array_index_75577[7];
  assign array_update_75585[8] = add_75532 == 32'h0000_0008 ? add_75583 : array_index_75577[8];
  assign array_update_75585[9] = add_75532 == 32'h0000_0009 ? add_75583 : array_index_75577[9];
  assign add_75586 = add_75573 + 32'h0000_0001;
  assign array_update_75587[0] = add_74719 == 32'h0000_0000 ? array_update_75585 : array_update_75574[0];
  assign array_update_75587[1] = add_74719 == 32'h0000_0001 ? array_update_75585 : array_update_75574[1];
  assign array_update_75587[2] = add_74719 == 32'h0000_0002 ? array_update_75585 : array_update_75574[2];
  assign array_update_75587[3] = add_74719 == 32'h0000_0003 ? array_update_75585 : array_update_75574[3];
  assign array_update_75587[4] = add_74719 == 32'h0000_0004 ? array_update_75585 : array_update_75574[4];
  assign array_update_75587[5] = add_74719 == 32'h0000_0005 ? array_update_75585 : array_update_75574[5];
  assign array_update_75587[6] = add_74719 == 32'h0000_0006 ? array_update_75585 : array_update_75574[6];
  assign array_update_75587[7] = add_74719 == 32'h0000_0007 ? array_update_75585 : array_update_75574[7];
  assign array_update_75587[8] = add_74719 == 32'h0000_0008 ? array_update_75585 : array_update_75574[8];
  assign array_update_75587[9] = add_74719 == 32'h0000_0009 ? array_update_75585 : array_update_75574[9];
  assign array_index_75589 = array_update_72021[add_75586 > 32'h0000_0009 ? 4'h9 : add_75586[3:0]];
  assign array_index_75590 = array_update_75587[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_75594 = smul32b_32b_x_32b(array_index_74726[add_75586 > 32'h0000_0009 ? 4'h9 : add_75586[3:0]], array_index_75589[add_75532 > 32'h0000_0009 ? 4'h9 : add_75532[3:0]]);
  assign add_75596 = array_index_75590[add_75532 > 32'h0000_0009 ? 4'h9 : add_75532[3:0]] + smul_75594;
  assign array_update_75598[0] = add_75532 == 32'h0000_0000 ? add_75596 : array_index_75590[0];
  assign array_update_75598[1] = add_75532 == 32'h0000_0001 ? add_75596 : array_index_75590[1];
  assign array_update_75598[2] = add_75532 == 32'h0000_0002 ? add_75596 : array_index_75590[2];
  assign array_update_75598[3] = add_75532 == 32'h0000_0003 ? add_75596 : array_index_75590[3];
  assign array_update_75598[4] = add_75532 == 32'h0000_0004 ? add_75596 : array_index_75590[4];
  assign array_update_75598[5] = add_75532 == 32'h0000_0005 ? add_75596 : array_index_75590[5];
  assign array_update_75598[6] = add_75532 == 32'h0000_0006 ? add_75596 : array_index_75590[6];
  assign array_update_75598[7] = add_75532 == 32'h0000_0007 ? add_75596 : array_index_75590[7];
  assign array_update_75598[8] = add_75532 == 32'h0000_0008 ? add_75596 : array_index_75590[8];
  assign array_update_75598[9] = add_75532 == 32'h0000_0009 ? add_75596 : array_index_75590[9];
  assign add_75599 = add_75586 + 32'h0000_0001;
  assign array_update_75600[0] = add_74719 == 32'h0000_0000 ? array_update_75598 : array_update_75587[0];
  assign array_update_75600[1] = add_74719 == 32'h0000_0001 ? array_update_75598 : array_update_75587[1];
  assign array_update_75600[2] = add_74719 == 32'h0000_0002 ? array_update_75598 : array_update_75587[2];
  assign array_update_75600[3] = add_74719 == 32'h0000_0003 ? array_update_75598 : array_update_75587[3];
  assign array_update_75600[4] = add_74719 == 32'h0000_0004 ? array_update_75598 : array_update_75587[4];
  assign array_update_75600[5] = add_74719 == 32'h0000_0005 ? array_update_75598 : array_update_75587[5];
  assign array_update_75600[6] = add_74719 == 32'h0000_0006 ? array_update_75598 : array_update_75587[6];
  assign array_update_75600[7] = add_74719 == 32'h0000_0007 ? array_update_75598 : array_update_75587[7];
  assign array_update_75600[8] = add_74719 == 32'h0000_0008 ? array_update_75598 : array_update_75587[8];
  assign array_update_75600[9] = add_74719 == 32'h0000_0009 ? array_update_75598 : array_update_75587[9];
  assign array_index_75602 = array_update_72021[add_75599 > 32'h0000_0009 ? 4'h9 : add_75599[3:0]];
  assign array_index_75603 = array_update_75600[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_75607 = smul32b_32b_x_32b(array_index_74726[add_75599 > 32'h0000_0009 ? 4'h9 : add_75599[3:0]], array_index_75602[add_75532 > 32'h0000_0009 ? 4'h9 : add_75532[3:0]]);
  assign add_75609 = array_index_75603[add_75532 > 32'h0000_0009 ? 4'h9 : add_75532[3:0]] + smul_75607;
  assign array_update_75611[0] = add_75532 == 32'h0000_0000 ? add_75609 : array_index_75603[0];
  assign array_update_75611[1] = add_75532 == 32'h0000_0001 ? add_75609 : array_index_75603[1];
  assign array_update_75611[2] = add_75532 == 32'h0000_0002 ? add_75609 : array_index_75603[2];
  assign array_update_75611[3] = add_75532 == 32'h0000_0003 ? add_75609 : array_index_75603[3];
  assign array_update_75611[4] = add_75532 == 32'h0000_0004 ? add_75609 : array_index_75603[4];
  assign array_update_75611[5] = add_75532 == 32'h0000_0005 ? add_75609 : array_index_75603[5];
  assign array_update_75611[6] = add_75532 == 32'h0000_0006 ? add_75609 : array_index_75603[6];
  assign array_update_75611[7] = add_75532 == 32'h0000_0007 ? add_75609 : array_index_75603[7];
  assign array_update_75611[8] = add_75532 == 32'h0000_0008 ? add_75609 : array_index_75603[8];
  assign array_update_75611[9] = add_75532 == 32'h0000_0009 ? add_75609 : array_index_75603[9];
  assign add_75612 = add_75599 + 32'h0000_0001;
  assign array_update_75613[0] = add_74719 == 32'h0000_0000 ? array_update_75611 : array_update_75600[0];
  assign array_update_75613[1] = add_74719 == 32'h0000_0001 ? array_update_75611 : array_update_75600[1];
  assign array_update_75613[2] = add_74719 == 32'h0000_0002 ? array_update_75611 : array_update_75600[2];
  assign array_update_75613[3] = add_74719 == 32'h0000_0003 ? array_update_75611 : array_update_75600[3];
  assign array_update_75613[4] = add_74719 == 32'h0000_0004 ? array_update_75611 : array_update_75600[4];
  assign array_update_75613[5] = add_74719 == 32'h0000_0005 ? array_update_75611 : array_update_75600[5];
  assign array_update_75613[6] = add_74719 == 32'h0000_0006 ? array_update_75611 : array_update_75600[6];
  assign array_update_75613[7] = add_74719 == 32'h0000_0007 ? array_update_75611 : array_update_75600[7];
  assign array_update_75613[8] = add_74719 == 32'h0000_0008 ? array_update_75611 : array_update_75600[8];
  assign array_update_75613[9] = add_74719 == 32'h0000_0009 ? array_update_75611 : array_update_75600[9];
  assign array_index_75615 = array_update_72021[add_75612 > 32'h0000_0009 ? 4'h9 : add_75612[3:0]];
  assign array_index_75616 = array_update_75613[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_75620 = smul32b_32b_x_32b(array_index_74726[add_75612 > 32'h0000_0009 ? 4'h9 : add_75612[3:0]], array_index_75615[add_75532 > 32'h0000_0009 ? 4'h9 : add_75532[3:0]]);
  assign add_75622 = array_index_75616[add_75532 > 32'h0000_0009 ? 4'h9 : add_75532[3:0]] + smul_75620;
  assign array_update_75624[0] = add_75532 == 32'h0000_0000 ? add_75622 : array_index_75616[0];
  assign array_update_75624[1] = add_75532 == 32'h0000_0001 ? add_75622 : array_index_75616[1];
  assign array_update_75624[2] = add_75532 == 32'h0000_0002 ? add_75622 : array_index_75616[2];
  assign array_update_75624[3] = add_75532 == 32'h0000_0003 ? add_75622 : array_index_75616[3];
  assign array_update_75624[4] = add_75532 == 32'h0000_0004 ? add_75622 : array_index_75616[4];
  assign array_update_75624[5] = add_75532 == 32'h0000_0005 ? add_75622 : array_index_75616[5];
  assign array_update_75624[6] = add_75532 == 32'h0000_0006 ? add_75622 : array_index_75616[6];
  assign array_update_75624[7] = add_75532 == 32'h0000_0007 ? add_75622 : array_index_75616[7];
  assign array_update_75624[8] = add_75532 == 32'h0000_0008 ? add_75622 : array_index_75616[8];
  assign array_update_75624[9] = add_75532 == 32'h0000_0009 ? add_75622 : array_index_75616[9];
  assign add_75625 = add_75612 + 32'h0000_0001;
  assign array_update_75626[0] = add_74719 == 32'h0000_0000 ? array_update_75624 : array_update_75613[0];
  assign array_update_75626[1] = add_74719 == 32'h0000_0001 ? array_update_75624 : array_update_75613[1];
  assign array_update_75626[2] = add_74719 == 32'h0000_0002 ? array_update_75624 : array_update_75613[2];
  assign array_update_75626[3] = add_74719 == 32'h0000_0003 ? array_update_75624 : array_update_75613[3];
  assign array_update_75626[4] = add_74719 == 32'h0000_0004 ? array_update_75624 : array_update_75613[4];
  assign array_update_75626[5] = add_74719 == 32'h0000_0005 ? array_update_75624 : array_update_75613[5];
  assign array_update_75626[6] = add_74719 == 32'h0000_0006 ? array_update_75624 : array_update_75613[6];
  assign array_update_75626[7] = add_74719 == 32'h0000_0007 ? array_update_75624 : array_update_75613[7];
  assign array_update_75626[8] = add_74719 == 32'h0000_0008 ? array_update_75624 : array_update_75613[8];
  assign array_update_75626[9] = add_74719 == 32'h0000_0009 ? array_update_75624 : array_update_75613[9];
  assign array_index_75628 = array_update_72021[add_75625 > 32'h0000_0009 ? 4'h9 : add_75625[3:0]];
  assign array_index_75629 = array_update_75626[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_75633 = smul32b_32b_x_32b(array_index_74726[add_75625 > 32'h0000_0009 ? 4'h9 : add_75625[3:0]], array_index_75628[add_75532 > 32'h0000_0009 ? 4'h9 : add_75532[3:0]]);
  assign add_75635 = array_index_75629[add_75532 > 32'h0000_0009 ? 4'h9 : add_75532[3:0]] + smul_75633;
  assign array_update_75637[0] = add_75532 == 32'h0000_0000 ? add_75635 : array_index_75629[0];
  assign array_update_75637[1] = add_75532 == 32'h0000_0001 ? add_75635 : array_index_75629[1];
  assign array_update_75637[2] = add_75532 == 32'h0000_0002 ? add_75635 : array_index_75629[2];
  assign array_update_75637[3] = add_75532 == 32'h0000_0003 ? add_75635 : array_index_75629[3];
  assign array_update_75637[4] = add_75532 == 32'h0000_0004 ? add_75635 : array_index_75629[4];
  assign array_update_75637[5] = add_75532 == 32'h0000_0005 ? add_75635 : array_index_75629[5];
  assign array_update_75637[6] = add_75532 == 32'h0000_0006 ? add_75635 : array_index_75629[6];
  assign array_update_75637[7] = add_75532 == 32'h0000_0007 ? add_75635 : array_index_75629[7];
  assign array_update_75637[8] = add_75532 == 32'h0000_0008 ? add_75635 : array_index_75629[8];
  assign array_update_75637[9] = add_75532 == 32'h0000_0009 ? add_75635 : array_index_75629[9];
  assign add_75638 = add_75625 + 32'h0000_0001;
  assign array_update_75639[0] = add_74719 == 32'h0000_0000 ? array_update_75637 : array_update_75626[0];
  assign array_update_75639[1] = add_74719 == 32'h0000_0001 ? array_update_75637 : array_update_75626[1];
  assign array_update_75639[2] = add_74719 == 32'h0000_0002 ? array_update_75637 : array_update_75626[2];
  assign array_update_75639[3] = add_74719 == 32'h0000_0003 ? array_update_75637 : array_update_75626[3];
  assign array_update_75639[4] = add_74719 == 32'h0000_0004 ? array_update_75637 : array_update_75626[4];
  assign array_update_75639[5] = add_74719 == 32'h0000_0005 ? array_update_75637 : array_update_75626[5];
  assign array_update_75639[6] = add_74719 == 32'h0000_0006 ? array_update_75637 : array_update_75626[6];
  assign array_update_75639[7] = add_74719 == 32'h0000_0007 ? array_update_75637 : array_update_75626[7];
  assign array_update_75639[8] = add_74719 == 32'h0000_0008 ? array_update_75637 : array_update_75626[8];
  assign array_update_75639[9] = add_74719 == 32'h0000_0009 ? array_update_75637 : array_update_75626[9];
  assign array_index_75641 = array_update_72021[add_75638 > 32'h0000_0009 ? 4'h9 : add_75638[3:0]];
  assign array_index_75642 = array_update_75639[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_75646 = smul32b_32b_x_32b(array_index_74726[add_75638 > 32'h0000_0009 ? 4'h9 : add_75638[3:0]], array_index_75641[add_75532 > 32'h0000_0009 ? 4'h9 : add_75532[3:0]]);
  assign add_75648 = array_index_75642[add_75532 > 32'h0000_0009 ? 4'h9 : add_75532[3:0]] + smul_75646;
  assign array_update_75650[0] = add_75532 == 32'h0000_0000 ? add_75648 : array_index_75642[0];
  assign array_update_75650[1] = add_75532 == 32'h0000_0001 ? add_75648 : array_index_75642[1];
  assign array_update_75650[2] = add_75532 == 32'h0000_0002 ? add_75648 : array_index_75642[2];
  assign array_update_75650[3] = add_75532 == 32'h0000_0003 ? add_75648 : array_index_75642[3];
  assign array_update_75650[4] = add_75532 == 32'h0000_0004 ? add_75648 : array_index_75642[4];
  assign array_update_75650[5] = add_75532 == 32'h0000_0005 ? add_75648 : array_index_75642[5];
  assign array_update_75650[6] = add_75532 == 32'h0000_0006 ? add_75648 : array_index_75642[6];
  assign array_update_75650[7] = add_75532 == 32'h0000_0007 ? add_75648 : array_index_75642[7];
  assign array_update_75650[8] = add_75532 == 32'h0000_0008 ? add_75648 : array_index_75642[8];
  assign array_update_75650[9] = add_75532 == 32'h0000_0009 ? add_75648 : array_index_75642[9];
  assign add_75651 = add_75638 + 32'h0000_0001;
  assign array_update_75652[0] = add_74719 == 32'h0000_0000 ? array_update_75650 : array_update_75639[0];
  assign array_update_75652[1] = add_74719 == 32'h0000_0001 ? array_update_75650 : array_update_75639[1];
  assign array_update_75652[2] = add_74719 == 32'h0000_0002 ? array_update_75650 : array_update_75639[2];
  assign array_update_75652[3] = add_74719 == 32'h0000_0003 ? array_update_75650 : array_update_75639[3];
  assign array_update_75652[4] = add_74719 == 32'h0000_0004 ? array_update_75650 : array_update_75639[4];
  assign array_update_75652[5] = add_74719 == 32'h0000_0005 ? array_update_75650 : array_update_75639[5];
  assign array_update_75652[6] = add_74719 == 32'h0000_0006 ? array_update_75650 : array_update_75639[6];
  assign array_update_75652[7] = add_74719 == 32'h0000_0007 ? array_update_75650 : array_update_75639[7];
  assign array_update_75652[8] = add_74719 == 32'h0000_0008 ? array_update_75650 : array_update_75639[8];
  assign array_update_75652[9] = add_74719 == 32'h0000_0009 ? array_update_75650 : array_update_75639[9];
  assign array_index_75654 = array_update_72021[add_75651 > 32'h0000_0009 ? 4'h9 : add_75651[3:0]];
  assign array_index_75655 = array_update_75652[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_75659 = smul32b_32b_x_32b(array_index_74726[add_75651 > 32'h0000_0009 ? 4'h9 : add_75651[3:0]], array_index_75654[add_75532 > 32'h0000_0009 ? 4'h9 : add_75532[3:0]]);
  assign add_75661 = array_index_75655[add_75532 > 32'h0000_0009 ? 4'h9 : add_75532[3:0]] + smul_75659;
  assign array_update_75662[0] = add_75532 == 32'h0000_0000 ? add_75661 : array_index_75655[0];
  assign array_update_75662[1] = add_75532 == 32'h0000_0001 ? add_75661 : array_index_75655[1];
  assign array_update_75662[2] = add_75532 == 32'h0000_0002 ? add_75661 : array_index_75655[2];
  assign array_update_75662[3] = add_75532 == 32'h0000_0003 ? add_75661 : array_index_75655[3];
  assign array_update_75662[4] = add_75532 == 32'h0000_0004 ? add_75661 : array_index_75655[4];
  assign array_update_75662[5] = add_75532 == 32'h0000_0005 ? add_75661 : array_index_75655[5];
  assign array_update_75662[6] = add_75532 == 32'h0000_0006 ? add_75661 : array_index_75655[6];
  assign array_update_75662[7] = add_75532 == 32'h0000_0007 ? add_75661 : array_index_75655[7];
  assign array_update_75662[8] = add_75532 == 32'h0000_0008 ? add_75661 : array_index_75655[8];
  assign array_update_75662[9] = add_75532 == 32'h0000_0009 ? add_75661 : array_index_75655[9];
  assign array_update_75663[0] = add_74719 == 32'h0000_0000 ? array_update_75662 : array_update_75652[0];
  assign array_update_75663[1] = add_74719 == 32'h0000_0001 ? array_update_75662 : array_update_75652[1];
  assign array_update_75663[2] = add_74719 == 32'h0000_0002 ? array_update_75662 : array_update_75652[2];
  assign array_update_75663[3] = add_74719 == 32'h0000_0003 ? array_update_75662 : array_update_75652[3];
  assign array_update_75663[4] = add_74719 == 32'h0000_0004 ? array_update_75662 : array_update_75652[4];
  assign array_update_75663[5] = add_74719 == 32'h0000_0005 ? array_update_75662 : array_update_75652[5];
  assign array_update_75663[6] = add_74719 == 32'h0000_0006 ? array_update_75662 : array_update_75652[6];
  assign array_update_75663[7] = add_74719 == 32'h0000_0007 ? array_update_75662 : array_update_75652[7];
  assign array_update_75663[8] = add_74719 == 32'h0000_0008 ? array_update_75662 : array_update_75652[8];
  assign array_update_75663[9] = add_74719 == 32'h0000_0009 ? array_update_75662 : array_update_75652[9];
  assign array_index_75665 = array_update_75663[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign add_75667 = add_75532 + 32'h0000_0001;
  assign array_update_75668[0] = add_75667 == 32'h0000_0000 ? 32'h0000_0000 : array_index_75665[0];
  assign array_update_75668[1] = add_75667 == 32'h0000_0001 ? 32'h0000_0000 : array_index_75665[1];
  assign array_update_75668[2] = add_75667 == 32'h0000_0002 ? 32'h0000_0000 : array_index_75665[2];
  assign array_update_75668[3] = add_75667 == 32'h0000_0003 ? 32'h0000_0000 : array_index_75665[3];
  assign array_update_75668[4] = add_75667 == 32'h0000_0004 ? 32'h0000_0000 : array_index_75665[4];
  assign array_update_75668[5] = add_75667 == 32'h0000_0005 ? 32'h0000_0000 : array_index_75665[5];
  assign array_update_75668[6] = add_75667 == 32'h0000_0006 ? 32'h0000_0000 : array_index_75665[6];
  assign array_update_75668[7] = add_75667 == 32'h0000_0007 ? 32'h0000_0000 : array_index_75665[7];
  assign array_update_75668[8] = add_75667 == 32'h0000_0008 ? 32'h0000_0000 : array_index_75665[8];
  assign array_update_75668[9] = add_75667 == 32'h0000_0009 ? 32'h0000_0000 : array_index_75665[9];
  assign literal_75669 = 32'h0000_0000;
  assign array_update_75670[0] = add_74719 == 32'h0000_0000 ? array_update_75668 : array_update_75663[0];
  assign array_update_75670[1] = add_74719 == 32'h0000_0001 ? array_update_75668 : array_update_75663[1];
  assign array_update_75670[2] = add_74719 == 32'h0000_0002 ? array_update_75668 : array_update_75663[2];
  assign array_update_75670[3] = add_74719 == 32'h0000_0003 ? array_update_75668 : array_update_75663[3];
  assign array_update_75670[4] = add_74719 == 32'h0000_0004 ? array_update_75668 : array_update_75663[4];
  assign array_update_75670[5] = add_74719 == 32'h0000_0005 ? array_update_75668 : array_update_75663[5];
  assign array_update_75670[6] = add_74719 == 32'h0000_0006 ? array_update_75668 : array_update_75663[6];
  assign array_update_75670[7] = add_74719 == 32'h0000_0007 ? array_update_75668 : array_update_75663[7];
  assign array_update_75670[8] = add_74719 == 32'h0000_0008 ? array_update_75668 : array_update_75663[8];
  assign array_update_75670[9] = add_74719 == 32'h0000_0009 ? array_update_75668 : array_update_75663[9];
  assign array_index_75672 = array_update_72021[literal_75669 > 32'h0000_0009 ? 4'h9 : literal_75669[3:0]];
  assign array_index_75673 = array_update_75670[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_75677 = smul32b_32b_x_32b(array_index_74726[literal_75669 > 32'h0000_0009 ? 4'h9 : literal_75669[3:0]], array_index_75672[add_75667 > 32'h0000_0009 ? 4'h9 : add_75667[3:0]]);
  assign add_75679 = array_index_75673[add_75667 > 32'h0000_0009 ? 4'h9 : add_75667[3:0]] + smul_75677;
  assign array_update_75681[0] = add_75667 == 32'h0000_0000 ? add_75679 : array_index_75673[0];
  assign array_update_75681[1] = add_75667 == 32'h0000_0001 ? add_75679 : array_index_75673[1];
  assign array_update_75681[2] = add_75667 == 32'h0000_0002 ? add_75679 : array_index_75673[2];
  assign array_update_75681[3] = add_75667 == 32'h0000_0003 ? add_75679 : array_index_75673[3];
  assign array_update_75681[4] = add_75667 == 32'h0000_0004 ? add_75679 : array_index_75673[4];
  assign array_update_75681[5] = add_75667 == 32'h0000_0005 ? add_75679 : array_index_75673[5];
  assign array_update_75681[6] = add_75667 == 32'h0000_0006 ? add_75679 : array_index_75673[6];
  assign array_update_75681[7] = add_75667 == 32'h0000_0007 ? add_75679 : array_index_75673[7];
  assign array_update_75681[8] = add_75667 == 32'h0000_0008 ? add_75679 : array_index_75673[8];
  assign array_update_75681[9] = add_75667 == 32'h0000_0009 ? add_75679 : array_index_75673[9];
  assign add_75682 = literal_75669 + 32'h0000_0001;
  assign array_update_75683[0] = add_74719 == 32'h0000_0000 ? array_update_75681 : array_update_75670[0];
  assign array_update_75683[1] = add_74719 == 32'h0000_0001 ? array_update_75681 : array_update_75670[1];
  assign array_update_75683[2] = add_74719 == 32'h0000_0002 ? array_update_75681 : array_update_75670[2];
  assign array_update_75683[3] = add_74719 == 32'h0000_0003 ? array_update_75681 : array_update_75670[3];
  assign array_update_75683[4] = add_74719 == 32'h0000_0004 ? array_update_75681 : array_update_75670[4];
  assign array_update_75683[5] = add_74719 == 32'h0000_0005 ? array_update_75681 : array_update_75670[5];
  assign array_update_75683[6] = add_74719 == 32'h0000_0006 ? array_update_75681 : array_update_75670[6];
  assign array_update_75683[7] = add_74719 == 32'h0000_0007 ? array_update_75681 : array_update_75670[7];
  assign array_update_75683[8] = add_74719 == 32'h0000_0008 ? array_update_75681 : array_update_75670[8];
  assign array_update_75683[9] = add_74719 == 32'h0000_0009 ? array_update_75681 : array_update_75670[9];
  assign array_index_75685 = array_update_72021[add_75682 > 32'h0000_0009 ? 4'h9 : add_75682[3:0]];
  assign array_index_75686 = array_update_75683[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_75690 = smul32b_32b_x_32b(array_index_74726[add_75682 > 32'h0000_0009 ? 4'h9 : add_75682[3:0]], array_index_75685[add_75667 > 32'h0000_0009 ? 4'h9 : add_75667[3:0]]);
  assign add_75692 = array_index_75686[add_75667 > 32'h0000_0009 ? 4'h9 : add_75667[3:0]] + smul_75690;
  assign array_update_75694[0] = add_75667 == 32'h0000_0000 ? add_75692 : array_index_75686[0];
  assign array_update_75694[1] = add_75667 == 32'h0000_0001 ? add_75692 : array_index_75686[1];
  assign array_update_75694[2] = add_75667 == 32'h0000_0002 ? add_75692 : array_index_75686[2];
  assign array_update_75694[3] = add_75667 == 32'h0000_0003 ? add_75692 : array_index_75686[3];
  assign array_update_75694[4] = add_75667 == 32'h0000_0004 ? add_75692 : array_index_75686[4];
  assign array_update_75694[5] = add_75667 == 32'h0000_0005 ? add_75692 : array_index_75686[5];
  assign array_update_75694[6] = add_75667 == 32'h0000_0006 ? add_75692 : array_index_75686[6];
  assign array_update_75694[7] = add_75667 == 32'h0000_0007 ? add_75692 : array_index_75686[7];
  assign array_update_75694[8] = add_75667 == 32'h0000_0008 ? add_75692 : array_index_75686[8];
  assign array_update_75694[9] = add_75667 == 32'h0000_0009 ? add_75692 : array_index_75686[9];
  assign add_75695 = add_75682 + 32'h0000_0001;
  assign array_update_75696[0] = add_74719 == 32'h0000_0000 ? array_update_75694 : array_update_75683[0];
  assign array_update_75696[1] = add_74719 == 32'h0000_0001 ? array_update_75694 : array_update_75683[1];
  assign array_update_75696[2] = add_74719 == 32'h0000_0002 ? array_update_75694 : array_update_75683[2];
  assign array_update_75696[3] = add_74719 == 32'h0000_0003 ? array_update_75694 : array_update_75683[3];
  assign array_update_75696[4] = add_74719 == 32'h0000_0004 ? array_update_75694 : array_update_75683[4];
  assign array_update_75696[5] = add_74719 == 32'h0000_0005 ? array_update_75694 : array_update_75683[5];
  assign array_update_75696[6] = add_74719 == 32'h0000_0006 ? array_update_75694 : array_update_75683[6];
  assign array_update_75696[7] = add_74719 == 32'h0000_0007 ? array_update_75694 : array_update_75683[7];
  assign array_update_75696[8] = add_74719 == 32'h0000_0008 ? array_update_75694 : array_update_75683[8];
  assign array_update_75696[9] = add_74719 == 32'h0000_0009 ? array_update_75694 : array_update_75683[9];
  assign array_index_75698 = array_update_72021[add_75695 > 32'h0000_0009 ? 4'h9 : add_75695[3:0]];
  assign array_index_75699 = array_update_75696[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_75703 = smul32b_32b_x_32b(array_index_74726[add_75695 > 32'h0000_0009 ? 4'h9 : add_75695[3:0]], array_index_75698[add_75667 > 32'h0000_0009 ? 4'h9 : add_75667[3:0]]);
  assign add_75705 = array_index_75699[add_75667 > 32'h0000_0009 ? 4'h9 : add_75667[3:0]] + smul_75703;
  assign array_update_75707[0] = add_75667 == 32'h0000_0000 ? add_75705 : array_index_75699[0];
  assign array_update_75707[1] = add_75667 == 32'h0000_0001 ? add_75705 : array_index_75699[1];
  assign array_update_75707[2] = add_75667 == 32'h0000_0002 ? add_75705 : array_index_75699[2];
  assign array_update_75707[3] = add_75667 == 32'h0000_0003 ? add_75705 : array_index_75699[3];
  assign array_update_75707[4] = add_75667 == 32'h0000_0004 ? add_75705 : array_index_75699[4];
  assign array_update_75707[5] = add_75667 == 32'h0000_0005 ? add_75705 : array_index_75699[5];
  assign array_update_75707[6] = add_75667 == 32'h0000_0006 ? add_75705 : array_index_75699[6];
  assign array_update_75707[7] = add_75667 == 32'h0000_0007 ? add_75705 : array_index_75699[7];
  assign array_update_75707[8] = add_75667 == 32'h0000_0008 ? add_75705 : array_index_75699[8];
  assign array_update_75707[9] = add_75667 == 32'h0000_0009 ? add_75705 : array_index_75699[9];
  assign add_75708 = add_75695 + 32'h0000_0001;
  assign array_update_75709[0] = add_74719 == 32'h0000_0000 ? array_update_75707 : array_update_75696[0];
  assign array_update_75709[1] = add_74719 == 32'h0000_0001 ? array_update_75707 : array_update_75696[1];
  assign array_update_75709[2] = add_74719 == 32'h0000_0002 ? array_update_75707 : array_update_75696[2];
  assign array_update_75709[3] = add_74719 == 32'h0000_0003 ? array_update_75707 : array_update_75696[3];
  assign array_update_75709[4] = add_74719 == 32'h0000_0004 ? array_update_75707 : array_update_75696[4];
  assign array_update_75709[5] = add_74719 == 32'h0000_0005 ? array_update_75707 : array_update_75696[5];
  assign array_update_75709[6] = add_74719 == 32'h0000_0006 ? array_update_75707 : array_update_75696[6];
  assign array_update_75709[7] = add_74719 == 32'h0000_0007 ? array_update_75707 : array_update_75696[7];
  assign array_update_75709[8] = add_74719 == 32'h0000_0008 ? array_update_75707 : array_update_75696[8];
  assign array_update_75709[9] = add_74719 == 32'h0000_0009 ? array_update_75707 : array_update_75696[9];
  assign array_index_75711 = array_update_72021[add_75708 > 32'h0000_0009 ? 4'h9 : add_75708[3:0]];
  assign array_index_75712 = array_update_75709[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_75716 = smul32b_32b_x_32b(array_index_74726[add_75708 > 32'h0000_0009 ? 4'h9 : add_75708[3:0]], array_index_75711[add_75667 > 32'h0000_0009 ? 4'h9 : add_75667[3:0]]);
  assign add_75718 = array_index_75712[add_75667 > 32'h0000_0009 ? 4'h9 : add_75667[3:0]] + smul_75716;
  assign array_update_75720[0] = add_75667 == 32'h0000_0000 ? add_75718 : array_index_75712[0];
  assign array_update_75720[1] = add_75667 == 32'h0000_0001 ? add_75718 : array_index_75712[1];
  assign array_update_75720[2] = add_75667 == 32'h0000_0002 ? add_75718 : array_index_75712[2];
  assign array_update_75720[3] = add_75667 == 32'h0000_0003 ? add_75718 : array_index_75712[3];
  assign array_update_75720[4] = add_75667 == 32'h0000_0004 ? add_75718 : array_index_75712[4];
  assign array_update_75720[5] = add_75667 == 32'h0000_0005 ? add_75718 : array_index_75712[5];
  assign array_update_75720[6] = add_75667 == 32'h0000_0006 ? add_75718 : array_index_75712[6];
  assign array_update_75720[7] = add_75667 == 32'h0000_0007 ? add_75718 : array_index_75712[7];
  assign array_update_75720[8] = add_75667 == 32'h0000_0008 ? add_75718 : array_index_75712[8];
  assign array_update_75720[9] = add_75667 == 32'h0000_0009 ? add_75718 : array_index_75712[9];
  assign add_75721 = add_75708 + 32'h0000_0001;
  assign array_update_75722[0] = add_74719 == 32'h0000_0000 ? array_update_75720 : array_update_75709[0];
  assign array_update_75722[1] = add_74719 == 32'h0000_0001 ? array_update_75720 : array_update_75709[1];
  assign array_update_75722[2] = add_74719 == 32'h0000_0002 ? array_update_75720 : array_update_75709[2];
  assign array_update_75722[3] = add_74719 == 32'h0000_0003 ? array_update_75720 : array_update_75709[3];
  assign array_update_75722[4] = add_74719 == 32'h0000_0004 ? array_update_75720 : array_update_75709[4];
  assign array_update_75722[5] = add_74719 == 32'h0000_0005 ? array_update_75720 : array_update_75709[5];
  assign array_update_75722[6] = add_74719 == 32'h0000_0006 ? array_update_75720 : array_update_75709[6];
  assign array_update_75722[7] = add_74719 == 32'h0000_0007 ? array_update_75720 : array_update_75709[7];
  assign array_update_75722[8] = add_74719 == 32'h0000_0008 ? array_update_75720 : array_update_75709[8];
  assign array_update_75722[9] = add_74719 == 32'h0000_0009 ? array_update_75720 : array_update_75709[9];
  assign array_index_75724 = array_update_72021[add_75721 > 32'h0000_0009 ? 4'h9 : add_75721[3:0]];
  assign array_index_75725 = array_update_75722[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_75729 = smul32b_32b_x_32b(array_index_74726[add_75721 > 32'h0000_0009 ? 4'h9 : add_75721[3:0]], array_index_75724[add_75667 > 32'h0000_0009 ? 4'h9 : add_75667[3:0]]);
  assign add_75731 = array_index_75725[add_75667 > 32'h0000_0009 ? 4'h9 : add_75667[3:0]] + smul_75729;
  assign array_update_75733[0] = add_75667 == 32'h0000_0000 ? add_75731 : array_index_75725[0];
  assign array_update_75733[1] = add_75667 == 32'h0000_0001 ? add_75731 : array_index_75725[1];
  assign array_update_75733[2] = add_75667 == 32'h0000_0002 ? add_75731 : array_index_75725[2];
  assign array_update_75733[3] = add_75667 == 32'h0000_0003 ? add_75731 : array_index_75725[3];
  assign array_update_75733[4] = add_75667 == 32'h0000_0004 ? add_75731 : array_index_75725[4];
  assign array_update_75733[5] = add_75667 == 32'h0000_0005 ? add_75731 : array_index_75725[5];
  assign array_update_75733[6] = add_75667 == 32'h0000_0006 ? add_75731 : array_index_75725[6];
  assign array_update_75733[7] = add_75667 == 32'h0000_0007 ? add_75731 : array_index_75725[7];
  assign array_update_75733[8] = add_75667 == 32'h0000_0008 ? add_75731 : array_index_75725[8];
  assign array_update_75733[9] = add_75667 == 32'h0000_0009 ? add_75731 : array_index_75725[9];
  assign add_75734 = add_75721 + 32'h0000_0001;
  assign array_update_75735[0] = add_74719 == 32'h0000_0000 ? array_update_75733 : array_update_75722[0];
  assign array_update_75735[1] = add_74719 == 32'h0000_0001 ? array_update_75733 : array_update_75722[1];
  assign array_update_75735[2] = add_74719 == 32'h0000_0002 ? array_update_75733 : array_update_75722[2];
  assign array_update_75735[3] = add_74719 == 32'h0000_0003 ? array_update_75733 : array_update_75722[3];
  assign array_update_75735[4] = add_74719 == 32'h0000_0004 ? array_update_75733 : array_update_75722[4];
  assign array_update_75735[5] = add_74719 == 32'h0000_0005 ? array_update_75733 : array_update_75722[5];
  assign array_update_75735[6] = add_74719 == 32'h0000_0006 ? array_update_75733 : array_update_75722[6];
  assign array_update_75735[7] = add_74719 == 32'h0000_0007 ? array_update_75733 : array_update_75722[7];
  assign array_update_75735[8] = add_74719 == 32'h0000_0008 ? array_update_75733 : array_update_75722[8];
  assign array_update_75735[9] = add_74719 == 32'h0000_0009 ? array_update_75733 : array_update_75722[9];
  assign array_index_75737 = array_update_72021[add_75734 > 32'h0000_0009 ? 4'h9 : add_75734[3:0]];
  assign array_index_75738 = array_update_75735[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_75742 = smul32b_32b_x_32b(array_index_74726[add_75734 > 32'h0000_0009 ? 4'h9 : add_75734[3:0]], array_index_75737[add_75667 > 32'h0000_0009 ? 4'h9 : add_75667[3:0]]);
  assign add_75744 = array_index_75738[add_75667 > 32'h0000_0009 ? 4'h9 : add_75667[3:0]] + smul_75742;
  assign array_update_75746[0] = add_75667 == 32'h0000_0000 ? add_75744 : array_index_75738[0];
  assign array_update_75746[1] = add_75667 == 32'h0000_0001 ? add_75744 : array_index_75738[1];
  assign array_update_75746[2] = add_75667 == 32'h0000_0002 ? add_75744 : array_index_75738[2];
  assign array_update_75746[3] = add_75667 == 32'h0000_0003 ? add_75744 : array_index_75738[3];
  assign array_update_75746[4] = add_75667 == 32'h0000_0004 ? add_75744 : array_index_75738[4];
  assign array_update_75746[5] = add_75667 == 32'h0000_0005 ? add_75744 : array_index_75738[5];
  assign array_update_75746[6] = add_75667 == 32'h0000_0006 ? add_75744 : array_index_75738[6];
  assign array_update_75746[7] = add_75667 == 32'h0000_0007 ? add_75744 : array_index_75738[7];
  assign array_update_75746[8] = add_75667 == 32'h0000_0008 ? add_75744 : array_index_75738[8];
  assign array_update_75746[9] = add_75667 == 32'h0000_0009 ? add_75744 : array_index_75738[9];
  assign add_75747 = add_75734 + 32'h0000_0001;
  assign array_update_75748[0] = add_74719 == 32'h0000_0000 ? array_update_75746 : array_update_75735[0];
  assign array_update_75748[1] = add_74719 == 32'h0000_0001 ? array_update_75746 : array_update_75735[1];
  assign array_update_75748[2] = add_74719 == 32'h0000_0002 ? array_update_75746 : array_update_75735[2];
  assign array_update_75748[3] = add_74719 == 32'h0000_0003 ? array_update_75746 : array_update_75735[3];
  assign array_update_75748[4] = add_74719 == 32'h0000_0004 ? array_update_75746 : array_update_75735[4];
  assign array_update_75748[5] = add_74719 == 32'h0000_0005 ? array_update_75746 : array_update_75735[5];
  assign array_update_75748[6] = add_74719 == 32'h0000_0006 ? array_update_75746 : array_update_75735[6];
  assign array_update_75748[7] = add_74719 == 32'h0000_0007 ? array_update_75746 : array_update_75735[7];
  assign array_update_75748[8] = add_74719 == 32'h0000_0008 ? array_update_75746 : array_update_75735[8];
  assign array_update_75748[9] = add_74719 == 32'h0000_0009 ? array_update_75746 : array_update_75735[9];
  assign array_index_75750 = array_update_72021[add_75747 > 32'h0000_0009 ? 4'h9 : add_75747[3:0]];
  assign array_index_75751 = array_update_75748[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_75755 = smul32b_32b_x_32b(array_index_74726[add_75747 > 32'h0000_0009 ? 4'h9 : add_75747[3:0]], array_index_75750[add_75667 > 32'h0000_0009 ? 4'h9 : add_75667[3:0]]);
  assign add_75757 = array_index_75751[add_75667 > 32'h0000_0009 ? 4'h9 : add_75667[3:0]] + smul_75755;
  assign array_update_75759[0] = add_75667 == 32'h0000_0000 ? add_75757 : array_index_75751[0];
  assign array_update_75759[1] = add_75667 == 32'h0000_0001 ? add_75757 : array_index_75751[1];
  assign array_update_75759[2] = add_75667 == 32'h0000_0002 ? add_75757 : array_index_75751[2];
  assign array_update_75759[3] = add_75667 == 32'h0000_0003 ? add_75757 : array_index_75751[3];
  assign array_update_75759[4] = add_75667 == 32'h0000_0004 ? add_75757 : array_index_75751[4];
  assign array_update_75759[5] = add_75667 == 32'h0000_0005 ? add_75757 : array_index_75751[5];
  assign array_update_75759[6] = add_75667 == 32'h0000_0006 ? add_75757 : array_index_75751[6];
  assign array_update_75759[7] = add_75667 == 32'h0000_0007 ? add_75757 : array_index_75751[7];
  assign array_update_75759[8] = add_75667 == 32'h0000_0008 ? add_75757 : array_index_75751[8];
  assign array_update_75759[9] = add_75667 == 32'h0000_0009 ? add_75757 : array_index_75751[9];
  assign add_75760 = add_75747 + 32'h0000_0001;
  assign array_update_75761[0] = add_74719 == 32'h0000_0000 ? array_update_75759 : array_update_75748[0];
  assign array_update_75761[1] = add_74719 == 32'h0000_0001 ? array_update_75759 : array_update_75748[1];
  assign array_update_75761[2] = add_74719 == 32'h0000_0002 ? array_update_75759 : array_update_75748[2];
  assign array_update_75761[3] = add_74719 == 32'h0000_0003 ? array_update_75759 : array_update_75748[3];
  assign array_update_75761[4] = add_74719 == 32'h0000_0004 ? array_update_75759 : array_update_75748[4];
  assign array_update_75761[5] = add_74719 == 32'h0000_0005 ? array_update_75759 : array_update_75748[5];
  assign array_update_75761[6] = add_74719 == 32'h0000_0006 ? array_update_75759 : array_update_75748[6];
  assign array_update_75761[7] = add_74719 == 32'h0000_0007 ? array_update_75759 : array_update_75748[7];
  assign array_update_75761[8] = add_74719 == 32'h0000_0008 ? array_update_75759 : array_update_75748[8];
  assign array_update_75761[9] = add_74719 == 32'h0000_0009 ? array_update_75759 : array_update_75748[9];
  assign array_index_75763 = array_update_72021[add_75760 > 32'h0000_0009 ? 4'h9 : add_75760[3:0]];
  assign array_index_75764 = array_update_75761[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_75768 = smul32b_32b_x_32b(array_index_74726[add_75760 > 32'h0000_0009 ? 4'h9 : add_75760[3:0]], array_index_75763[add_75667 > 32'h0000_0009 ? 4'h9 : add_75667[3:0]]);
  assign add_75770 = array_index_75764[add_75667 > 32'h0000_0009 ? 4'h9 : add_75667[3:0]] + smul_75768;
  assign array_update_75772[0] = add_75667 == 32'h0000_0000 ? add_75770 : array_index_75764[0];
  assign array_update_75772[1] = add_75667 == 32'h0000_0001 ? add_75770 : array_index_75764[1];
  assign array_update_75772[2] = add_75667 == 32'h0000_0002 ? add_75770 : array_index_75764[2];
  assign array_update_75772[3] = add_75667 == 32'h0000_0003 ? add_75770 : array_index_75764[3];
  assign array_update_75772[4] = add_75667 == 32'h0000_0004 ? add_75770 : array_index_75764[4];
  assign array_update_75772[5] = add_75667 == 32'h0000_0005 ? add_75770 : array_index_75764[5];
  assign array_update_75772[6] = add_75667 == 32'h0000_0006 ? add_75770 : array_index_75764[6];
  assign array_update_75772[7] = add_75667 == 32'h0000_0007 ? add_75770 : array_index_75764[7];
  assign array_update_75772[8] = add_75667 == 32'h0000_0008 ? add_75770 : array_index_75764[8];
  assign array_update_75772[9] = add_75667 == 32'h0000_0009 ? add_75770 : array_index_75764[9];
  assign add_75773 = add_75760 + 32'h0000_0001;
  assign array_update_75774[0] = add_74719 == 32'h0000_0000 ? array_update_75772 : array_update_75761[0];
  assign array_update_75774[1] = add_74719 == 32'h0000_0001 ? array_update_75772 : array_update_75761[1];
  assign array_update_75774[2] = add_74719 == 32'h0000_0002 ? array_update_75772 : array_update_75761[2];
  assign array_update_75774[3] = add_74719 == 32'h0000_0003 ? array_update_75772 : array_update_75761[3];
  assign array_update_75774[4] = add_74719 == 32'h0000_0004 ? array_update_75772 : array_update_75761[4];
  assign array_update_75774[5] = add_74719 == 32'h0000_0005 ? array_update_75772 : array_update_75761[5];
  assign array_update_75774[6] = add_74719 == 32'h0000_0006 ? array_update_75772 : array_update_75761[6];
  assign array_update_75774[7] = add_74719 == 32'h0000_0007 ? array_update_75772 : array_update_75761[7];
  assign array_update_75774[8] = add_74719 == 32'h0000_0008 ? array_update_75772 : array_update_75761[8];
  assign array_update_75774[9] = add_74719 == 32'h0000_0009 ? array_update_75772 : array_update_75761[9];
  assign array_index_75776 = array_update_72021[add_75773 > 32'h0000_0009 ? 4'h9 : add_75773[3:0]];
  assign array_index_75777 = array_update_75774[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_75781 = smul32b_32b_x_32b(array_index_74726[add_75773 > 32'h0000_0009 ? 4'h9 : add_75773[3:0]], array_index_75776[add_75667 > 32'h0000_0009 ? 4'h9 : add_75667[3:0]]);
  assign add_75783 = array_index_75777[add_75667 > 32'h0000_0009 ? 4'h9 : add_75667[3:0]] + smul_75781;
  assign array_update_75785[0] = add_75667 == 32'h0000_0000 ? add_75783 : array_index_75777[0];
  assign array_update_75785[1] = add_75667 == 32'h0000_0001 ? add_75783 : array_index_75777[1];
  assign array_update_75785[2] = add_75667 == 32'h0000_0002 ? add_75783 : array_index_75777[2];
  assign array_update_75785[3] = add_75667 == 32'h0000_0003 ? add_75783 : array_index_75777[3];
  assign array_update_75785[4] = add_75667 == 32'h0000_0004 ? add_75783 : array_index_75777[4];
  assign array_update_75785[5] = add_75667 == 32'h0000_0005 ? add_75783 : array_index_75777[5];
  assign array_update_75785[6] = add_75667 == 32'h0000_0006 ? add_75783 : array_index_75777[6];
  assign array_update_75785[7] = add_75667 == 32'h0000_0007 ? add_75783 : array_index_75777[7];
  assign array_update_75785[8] = add_75667 == 32'h0000_0008 ? add_75783 : array_index_75777[8];
  assign array_update_75785[9] = add_75667 == 32'h0000_0009 ? add_75783 : array_index_75777[9];
  assign add_75786 = add_75773 + 32'h0000_0001;
  assign array_update_75787[0] = add_74719 == 32'h0000_0000 ? array_update_75785 : array_update_75774[0];
  assign array_update_75787[1] = add_74719 == 32'h0000_0001 ? array_update_75785 : array_update_75774[1];
  assign array_update_75787[2] = add_74719 == 32'h0000_0002 ? array_update_75785 : array_update_75774[2];
  assign array_update_75787[3] = add_74719 == 32'h0000_0003 ? array_update_75785 : array_update_75774[3];
  assign array_update_75787[4] = add_74719 == 32'h0000_0004 ? array_update_75785 : array_update_75774[4];
  assign array_update_75787[5] = add_74719 == 32'h0000_0005 ? array_update_75785 : array_update_75774[5];
  assign array_update_75787[6] = add_74719 == 32'h0000_0006 ? array_update_75785 : array_update_75774[6];
  assign array_update_75787[7] = add_74719 == 32'h0000_0007 ? array_update_75785 : array_update_75774[7];
  assign array_update_75787[8] = add_74719 == 32'h0000_0008 ? array_update_75785 : array_update_75774[8];
  assign array_update_75787[9] = add_74719 == 32'h0000_0009 ? array_update_75785 : array_update_75774[9];
  assign array_index_75789 = array_update_72021[add_75786 > 32'h0000_0009 ? 4'h9 : add_75786[3:0]];
  assign array_index_75790 = array_update_75787[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_75794 = smul32b_32b_x_32b(array_index_74726[add_75786 > 32'h0000_0009 ? 4'h9 : add_75786[3:0]], array_index_75789[add_75667 > 32'h0000_0009 ? 4'h9 : add_75667[3:0]]);
  assign add_75796 = array_index_75790[add_75667 > 32'h0000_0009 ? 4'h9 : add_75667[3:0]] + smul_75794;
  assign array_update_75797[0] = add_75667 == 32'h0000_0000 ? add_75796 : array_index_75790[0];
  assign array_update_75797[1] = add_75667 == 32'h0000_0001 ? add_75796 : array_index_75790[1];
  assign array_update_75797[2] = add_75667 == 32'h0000_0002 ? add_75796 : array_index_75790[2];
  assign array_update_75797[3] = add_75667 == 32'h0000_0003 ? add_75796 : array_index_75790[3];
  assign array_update_75797[4] = add_75667 == 32'h0000_0004 ? add_75796 : array_index_75790[4];
  assign array_update_75797[5] = add_75667 == 32'h0000_0005 ? add_75796 : array_index_75790[5];
  assign array_update_75797[6] = add_75667 == 32'h0000_0006 ? add_75796 : array_index_75790[6];
  assign array_update_75797[7] = add_75667 == 32'h0000_0007 ? add_75796 : array_index_75790[7];
  assign array_update_75797[8] = add_75667 == 32'h0000_0008 ? add_75796 : array_index_75790[8];
  assign array_update_75797[9] = add_75667 == 32'h0000_0009 ? add_75796 : array_index_75790[9];
  assign array_update_75798[0] = add_74719 == 32'h0000_0000 ? array_update_75797 : array_update_75787[0];
  assign array_update_75798[1] = add_74719 == 32'h0000_0001 ? array_update_75797 : array_update_75787[1];
  assign array_update_75798[2] = add_74719 == 32'h0000_0002 ? array_update_75797 : array_update_75787[2];
  assign array_update_75798[3] = add_74719 == 32'h0000_0003 ? array_update_75797 : array_update_75787[3];
  assign array_update_75798[4] = add_74719 == 32'h0000_0004 ? array_update_75797 : array_update_75787[4];
  assign array_update_75798[5] = add_74719 == 32'h0000_0005 ? array_update_75797 : array_update_75787[5];
  assign array_update_75798[6] = add_74719 == 32'h0000_0006 ? array_update_75797 : array_update_75787[6];
  assign array_update_75798[7] = add_74719 == 32'h0000_0007 ? array_update_75797 : array_update_75787[7];
  assign array_update_75798[8] = add_74719 == 32'h0000_0008 ? array_update_75797 : array_update_75787[8];
  assign array_update_75798[9] = add_74719 == 32'h0000_0009 ? array_update_75797 : array_update_75787[9];
  assign array_index_75800 = array_update_75798[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign add_75802 = add_75667 + 32'h0000_0001;
  assign array_update_75803[0] = add_75802 == 32'h0000_0000 ? 32'h0000_0000 : array_index_75800[0];
  assign array_update_75803[1] = add_75802 == 32'h0000_0001 ? 32'h0000_0000 : array_index_75800[1];
  assign array_update_75803[2] = add_75802 == 32'h0000_0002 ? 32'h0000_0000 : array_index_75800[2];
  assign array_update_75803[3] = add_75802 == 32'h0000_0003 ? 32'h0000_0000 : array_index_75800[3];
  assign array_update_75803[4] = add_75802 == 32'h0000_0004 ? 32'h0000_0000 : array_index_75800[4];
  assign array_update_75803[5] = add_75802 == 32'h0000_0005 ? 32'h0000_0000 : array_index_75800[5];
  assign array_update_75803[6] = add_75802 == 32'h0000_0006 ? 32'h0000_0000 : array_index_75800[6];
  assign array_update_75803[7] = add_75802 == 32'h0000_0007 ? 32'h0000_0000 : array_index_75800[7];
  assign array_update_75803[8] = add_75802 == 32'h0000_0008 ? 32'h0000_0000 : array_index_75800[8];
  assign array_update_75803[9] = add_75802 == 32'h0000_0009 ? 32'h0000_0000 : array_index_75800[9];
  assign literal_75804 = 32'h0000_0000;
  assign array_update_75805[0] = add_74719 == 32'h0000_0000 ? array_update_75803 : array_update_75798[0];
  assign array_update_75805[1] = add_74719 == 32'h0000_0001 ? array_update_75803 : array_update_75798[1];
  assign array_update_75805[2] = add_74719 == 32'h0000_0002 ? array_update_75803 : array_update_75798[2];
  assign array_update_75805[3] = add_74719 == 32'h0000_0003 ? array_update_75803 : array_update_75798[3];
  assign array_update_75805[4] = add_74719 == 32'h0000_0004 ? array_update_75803 : array_update_75798[4];
  assign array_update_75805[5] = add_74719 == 32'h0000_0005 ? array_update_75803 : array_update_75798[5];
  assign array_update_75805[6] = add_74719 == 32'h0000_0006 ? array_update_75803 : array_update_75798[6];
  assign array_update_75805[7] = add_74719 == 32'h0000_0007 ? array_update_75803 : array_update_75798[7];
  assign array_update_75805[8] = add_74719 == 32'h0000_0008 ? array_update_75803 : array_update_75798[8];
  assign array_update_75805[9] = add_74719 == 32'h0000_0009 ? array_update_75803 : array_update_75798[9];
  assign array_index_75807 = array_update_72021[literal_75804 > 32'h0000_0009 ? 4'h9 : literal_75804[3:0]];
  assign array_index_75808 = array_update_75805[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_75812 = smul32b_32b_x_32b(array_index_74726[literal_75804 > 32'h0000_0009 ? 4'h9 : literal_75804[3:0]], array_index_75807[add_75802 > 32'h0000_0009 ? 4'h9 : add_75802[3:0]]);
  assign add_75814 = array_index_75808[add_75802 > 32'h0000_0009 ? 4'h9 : add_75802[3:0]] + smul_75812;
  assign array_update_75816[0] = add_75802 == 32'h0000_0000 ? add_75814 : array_index_75808[0];
  assign array_update_75816[1] = add_75802 == 32'h0000_0001 ? add_75814 : array_index_75808[1];
  assign array_update_75816[2] = add_75802 == 32'h0000_0002 ? add_75814 : array_index_75808[2];
  assign array_update_75816[3] = add_75802 == 32'h0000_0003 ? add_75814 : array_index_75808[3];
  assign array_update_75816[4] = add_75802 == 32'h0000_0004 ? add_75814 : array_index_75808[4];
  assign array_update_75816[5] = add_75802 == 32'h0000_0005 ? add_75814 : array_index_75808[5];
  assign array_update_75816[6] = add_75802 == 32'h0000_0006 ? add_75814 : array_index_75808[6];
  assign array_update_75816[7] = add_75802 == 32'h0000_0007 ? add_75814 : array_index_75808[7];
  assign array_update_75816[8] = add_75802 == 32'h0000_0008 ? add_75814 : array_index_75808[8];
  assign array_update_75816[9] = add_75802 == 32'h0000_0009 ? add_75814 : array_index_75808[9];
  assign add_75817 = literal_75804 + 32'h0000_0001;
  assign array_update_75818[0] = add_74719 == 32'h0000_0000 ? array_update_75816 : array_update_75805[0];
  assign array_update_75818[1] = add_74719 == 32'h0000_0001 ? array_update_75816 : array_update_75805[1];
  assign array_update_75818[2] = add_74719 == 32'h0000_0002 ? array_update_75816 : array_update_75805[2];
  assign array_update_75818[3] = add_74719 == 32'h0000_0003 ? array_update_75816 : array_update_75805[3];
  assign array_update_75818[4] = add_74719 == 32'h0000_0004 ? array_update_75816 : array_update_75805[4];
  assign array_update_75818[5] = add_74719 == 32'h0000_0005 ? array_update_75816 : array_update_75805[5];
  assign array_update_75818[6] = add_74719 == 32'h0000_0006 ? array_update_75816 : array_update_75805[6];
  assign array_update_75818[7] = add_74719 == 32'h0000_0007 ? array_update_75816 : array_update_75805[7];
  assign array_update_75818[8] = add_74719 == 32'h0000_0008 ? array_update_75816 : array_update_75805[8];
  assign array_update_75818[9] = add_74719 == 32'h0000_0009 ? array_update_75816 : array_update_75805[9];
  assign array_index_75820 = array_update_72021[add_75817 > 32'h0000_0009 ? 4'h9 : add_75817[3:0]];
  assign array_index_75821 = array_update_75818[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_75825 = smul32b_32b_x_32b(array_index_74726[add_75817 > 32'h0000_0009 ? 4'h9 : add_75817[3:0]], array_index_75820[add_75802 > 32'h0000_0009 ? 4'h9 : add_75802[3:0]]);
  assign add_75827 = array_index_75821[add_75802 > 32'h0000_0009 ? 4'h9 : add_75802[3:0]] + smul_75825;
  assign array_update_75829[0] = add_75802 == 32'h0000_0000 ? add_75827 : array_index_75821[0];
  assign array_update_75829[1] = add_75802 == 32'h0000_0001 ? add_75827 : array_index_75821[1];
  assign array_update_75829[2] = add_75802 == 32'h0000_0002 ? add_75827 : array_index_75821[2];
  assign array_update_75829[3] = add_75802 == 32'h0000_0003 ? add_75827 : array_index_75821[3];
  assign array_update_75829[4] = add_75802 == 32'h0000_0004 ? add_75827 : array_index_75821[4];
  assign array_update_75829[5] = add_75802 == 32'h0000_0005 ? add_75827 : array_index_75821[5];
  assign array_update_75829[6] = add_75802 == 32'h0000_0006 ? add_75827 : array_index_75821[6];
  assign array_update_75829[7] = add_75802 == 32'h0000_0007 ? add_75827 : array_index_75821[7];
  assign array_update_75829[8] = add_75802 == 32'h0000_0008 ? add_75827 : array_index_75821[8];
  assign array_update_75829[9] = add_75802 == 32'h0000_0009 ? add_75827 : array_index_75821[9];
  assign add_75830 = add_75817 + 32'h0000_0001;
  assign array_update_75831[0] = add_74719 == 32'h0000_0000 ? array_update_75829 : array_update_75818[0];
  assign array_update_75831[1] = add_74719 == 32'h0000_0001 ? array_update_75829 : array_update_75818[1];
  assign array_update_75831[2] = add_74719 == 32'h0000_0002 ? array_update_75829 : array_update_75818[2];
  assign array_update_75831[3] = add_74719 == 32'h0000_0003 ? array_update_75829 : array_update_75818[3];
  assign array_update_75831[4] = add_74719 == 32'h0000_0004 ? array_update_75829 : array_update_75818[4];
  assign array_update_75831[5] = add_74719 == 32'h0000_0005 ? array_update_75829 : array_update_75818[5];
  assign array_update_75831[6] = add_74719 == 32'h0000_0006 ? array_update_75829 : array_update_75818[6];
  assign array_update_75831[7] = add_74719 == 32'h0000_0007 ? array_update_75829 : array_update_75818[7];
  assign array_update_75831[8] = add_74719 == 32'h0000_0008 ? array_update_75829 : array_update_75818[8];
  assign array_update_75831[9] = add_74719 == 32'h0000_0009 ? array_update_75829 : array_update_75818[9];
  assign array_index_75833 = array_update_72021[add_75830 > 32'h0000_0009 ? 4'h9 : add_75830[3:0]];
  assign array_index_75834 = array_update_75831[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_75838 = smul32b_32b_x_32b(array_index_74726[add_75830 > 32'h0000_0009 ? 4'h9 : add_75830[3:0]], array_index_75833[add_75802 > 32'h0000_0009 ? 4'h9 : add_75802[3:0]]);
  assign add_75840 = array_index_75834[add_75802 > 32'h0000_0009 ? 4'h9 : add_75802[3:0]] + smul_75838;
  assign array_update_75842[0] = add_75802 == 32'h0000_0000 ? add_75840 : array_index_75834[0];
  assign array_update_75842[1] = add_75802 == 32'h0000_0001 ? add_75840 : array_index_75834[1];
  assign array_update_75842[2] = add_75802 == 32'h0000_0002 ? add_75840 : array_index_75834[2];
  assign array_update_75842[3] = add_75802 == 32'h0000_0003 ? add_75840 : array_index_75834[3];
  assign array_update_75842[4] = add_75802 == 32'h0000_0004 ? add_75840 : array_index_75834[4];
  assign array_update_75842[5] = add_75802 == 32'h0000_0005 ? add_75840 : array_index_75834[5];
  assign array_update_75842[6] = add_75802 == 32'h0000_0006 ? add_75840 : array_index_75834[6];
  assign array_update_75842[7] = add_75802 == 32'h0000_0007 ? add_75840 : array_index_75834[7];
  assign array_update_75842[8] = add_75802 == 32'h0000_0008 ? add_75840 : array_index_75834[8];
  assign array_update_75842[9] = add_75802 == 32'h0000_0009 ? add_75840 : array_index_75834[9];
  assign add_75843 = add_75830 + 32'h0000_0001;
  assign array_update_75844[0] = add_74719 == 32'h0000_0000 ? array_update_75842 : array_update_75831[0];
  assign array_update_75844[1] = add_74719 == 32'h0000_0001 ? array_update_75842 : array_update_75831[1];
  assign array_update_75844[2] = add_74719 == 32'h0000_0002 ? array_update_75842 : array_update_75831[2];
  assign array_update_75844[3] = add_74719 == 32'h0000_0003 ? array_update_75842 : array_update_75831[3];
  assign array_update_75844[4] = add_74719 == 32'h0000_0004 ? array_update_75842 : array_update_75831[4];
  assign array_update_75844[5] = add_74719 == 32'h0000_0005 ? array_update_75842 : array_update_75831[5];
  assign array_update_75844[6] = add_74719 == 32'h0000_0006 ? array_update_75842 : array_update_75831[6];
  assign array_update_75844[7] = add_74719 == 32'h0000_0007 ? array_update_75842 : array_update_75831[7];
  assign array_update_75844[8] = add_74719 == 32'h0000_0008 ? array_update_75842 : array_update_75831[8];
  assign array_update_75844[9] = add_74719 == 32'h0000_0009 ? array_update_75842 : array_update_75831[9];
  assign array_index_75846 = array_update_72021[add_75843 > 32'h0000_0009 ? 4'h9 : add_75843[3:0]];
  assign array_index_75847 = array_update_75844[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_75851 = smul32b_32b_x_32b(array_index_74726[add_75843 > 32'h0000_0009 ? 4'h9 : add_75843[3:0]], array_index_75846[add_75802 > 32'h0000_0009 ? 4'h9 : add_75802[3:0]]);
  assign add_75853 = array_index_75847[add_75802 > 32'h0000_0009 ? 4'h9 : add_75802[3:0]] + smul_75851;
  assign array_update_75855[0] = add_75802 == 32'h0000_0000 ? add_75853 : array_index_75847[0];
  assign array_update_75855[1] = add_75802 == 32'h0000_0001 ? add_75853 : array_index_75847[1];
  assign array_update_75855[2] = add_75802 == 32'h0000_0002 ? add_75853 : array_index_75847[2];
  assign array_update_75855[3] = add_75802 == 32'h0000_0003 ? add_75853 : array_index_75847[3];
  assign array_update_75855[4] = add_75802 == 32'h0000_0004 ? add_75853 : array_index_75847[4];
  assign array_update_75855[5] = add_75802 == 32'h0000_0005 ? add_75853 : array_index_75847[5];
  assign array_update_75855[6] = add_75802 == 32'h0000_0006 ? add_75853 : array_index_75847[6];
  assign array_update_75855[7] = add_75802 == 32'h0000_0007 ? add_75853 : array_index_75847[7];
  assign array_update_75855[8] = add_75802 == 32'h0000_0008 ? add_75853 : array_index_75847[8];
  assign array_update_75855[9] = add_75802 == 32'h0000_0009 ? add_75853 : array_index_75847[9];
  assign add_75856 = add_75843 + 32'h0000_0001;
  assign array_update_75857[0] = add_74719 == 32'h0000_0000 ? array_update_75855 : array_update_75844[0];
  assign array_update_75857[1] = add_74719 == 32'h0000_0001 ? array_update_75855 : array_update_75844[1];
  assign array_update_75857[2] = add_74719 == 32'h0000_0002 ? array_update_75855 : array_update_75844[2];
  assign array_update_75857[3] = add_74719 == 32'h0000_0003 ? array_update_75855 : array_update_75844[3];
  assign array_update_75857[4] = add_74719 == 32'h0000_0004 ? array_update_75855 : array_update_75844[4];
  assign array_update_75857[5] = add_74719 == 32'h0000_0005 ? array_update_75855 : array_update_75844[5];
  assign array_update_75857[6] = add_74719 == 32'h0000_0006 ? array_update_75855 : array_update_75844[6];
  assign array_update_75857[7] = add_74719 == 32'h0000_0007 ? array_update_75855 : array_update_75844[7];
  assign array_update_75857[8] = add_74719 == 32'h0000_0008 ? array_update_75855 : array_update_75844[8];
  assign array_update_75857[9] = add_74719 == 32'h0000_0009 ? array_update_75855 : array_update_75844[9];
  assign array_index_75859 = array_update_72021[add_75856 > 32'h0000_0009 ? 4'h9 : add_75856[3:0]];
  assign array_index_75860 = array_update_75857[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_75864 = smul32b_32b_x_32b(array_index_74726[add_75856 > 32'h0000_0009 ? 4'h9 : add_75856[3:0]], array_index_75859[add_75802 > 32'h0000_0009 ? 4'h9 : add_75802[3:0]]);
  assign add_75866 = array_index_75860[add_75802 > 32'h0000_0009 ? 4'h9 : add_75802[3:0]] + smul_75864;
  assign array_update_75868[0] = add_75802 == 32'h0000_0000 ? add_75866 : array_index_75860[0];
  assign array_update_75868[1] = add_75802 == 32'h0000_0001 ? add_75866 : array_index_75860[1];
  assign array_update_75868[2] = add_75802 == 32'h0000_0002 ? add_75866 : array_index_75860[2];
  assign array_update_75868[3] = add_75802 == 32'h0000_0003 ? add_75866 : array_index_75860[3];
  assign array_update_75868[4] = add_75802 == 32'h0000_0004 ? add_75866 : array_index_75860[4];
  assign array_update_75868[5] = add_75802 == 32'h0000_0005 ? add_75866 : array_index_75860[5];
  assign array_update_75868[6] = add_75802 == 32'h0000_0006 ? add_75866 : array_index_75860[6];
  assign array_update_75868[7] = add_75802 == 32'h0000_0007 ? add_75866 : array_index_75860[7];
  assign array_update_75868[8] = add_75802 == 32'h0000_0008 ? add_75866 : array_index_75860[8];
  assign array_update_75868[9] = add_75802 == 32'h0000_0009 ? add_75866 : array_index_75860[9];
  assign add_75869 = add_75856 + 32'h0000_0001;
  assign array_update_75870[0] = add_74719 == 32'h0000_0000 ? array_update_75868 : array_update_75857[0];
  assign array_update_75870[1] = add_74719 == 32'h0000_0001 ? array_update_75868 : array_update_75857[1];
  assign array_update_75870[2] = add_74719 == 32'h0000_0002 ? array_update_75868 : array_update_75857[2];
  assign array_update_75870[3] = add_74719 == 32'h0000_0003 ? array_update_75868 : array_update_75857[3];
  assign array_update_75870[4] = add_74719 == 32'h0000_0004 ? array_update_75868 : array_update_75857[4];
  assign array_update_75870[5] = add_74719 == 32'h0000_0005 ? array_update_75868 : array_update_75857[5];
  assign array_update_75870[6] = add_74719 == 32'h0000_0006 ? array_update_75868 : array_update_75857[6];
  assign array_update_75870[7] = add_74719 == 32'h0000_0007 ? array_update_75868 : array_update_75857[7];
  assign array_update_75870[8] = add_74719 == 32'h0000_0008 ? array_update_75868 : array_update_75857[8];
  assign array_update_75870[9] = add_74719 == 32'h0000_0009 ? array_update_75868 : array_update_75857[9];
  assign array_index_75872 = array_update_72021[add_75869 > 32'h0000_0009 ? 4'h9 : add_75869[3:0]];
  assign array_index_75873 = array_update_75870[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_75877 = smul32b_32b_x_32b(array_index_74726[add_75869 > 32'h0000_0009 ? 4'h9 : add_75869[3:0]], array_index_75872[add_75802 > 32'h0000_0009 ? 4'h9 : add_75802[3:0]]);
  assign add_75879 = array_index_75873[add_75802 > 32'h0000_0009 ? 4'h9 : add_75802[3:0]] + smul_75877;
  assign array_update_75881[0] = add_75802 == 32'h0000_0000 ? add_75879 : array_index_75873[0];
  assign array_update_75881[1] = add_75802 == 32'h0000_0001 ? add_75879 : array_index_75873[1];
  assign array_update_75881[2] = add_75802 == 32'h0000_0002 ? add_75879 : array_index_75873[2];
  assign array_update_75881[3] = add_75802 == 32'h0000_0003 ? add_75879 : array_index_75873[3];
  assign array_update_75881[4] = add_75802 == 32'h0000_0004 ? add_75879 : array_index_75873[4];
  assign array_update_75881[5] = add_75802 == 32'h0000_0005 ? add_75879 : array_index_75873[5];
  assign array_update_75881[6] = add_75802 == 32'h0000_0006 ? add_75879 : array_index_75873[6];
  assign array_update_75881[7] = add_75802 == 32'h0000_0007 ? add_75879 : array_index_75873[7];
  assign array_update_75881[8] = add_75802 == 32'h0000_0008 ? add_75879 : array_index_75873[8];
  assign array_update_75881[9] = add_75802 == 32'h0000_0009 ? add_75879 : array_index_75873[9];
  assign add_75882 = add_75869 + 32'h0000_0001;
  assign array_update_75883[0] = add_74719 == 32'h0000_0000 ? array_update_75881 : array_update_75870[0];
  assign array_update_75883[1] = add_74719 == 32'h0000_0001 ? array_update_75881 : array_update_75870[1];
  assign array_update_75883[2] = add_74719 == 32'h0000_0002 ? array_update_75881 : array_update_75870[2];
  assign array_update_75883[3] = add_74719 == 32'h0000_0003 ? array_update_75881 : array_update_75870[3];
  assign array_update_75883[4] = add_74719 == 32'h0000_0004 ? array_update_75881 : array_update_75870[4];
  assign array_update_75883[5] = add_74719 == 32'h0000_0005 ? array_update_75881 : array_update_75870[5];
  assign array_update_75883[6] = add_74719 == 32'h0000_0006 ? array_update_75881 : array_update_75870[6];
  assign array_update_75883[7] = add_74719 == 32'h0000_0007 ? array_update_75881 : array_update_75870[7];
  assign array_update_75883[8] = add_74719 == 32'h0000_0008 ? array_update_75881 : array_update_75870[8];
  assign array_update_75883[9] = add_74719 == 32'h0000_0009 ? array_update_75881 : array_update_75870[9];
  assign array_index_75885 = array_update_72021[add_75882 > 32'h0000_0009 ? 4'h9 : add_75882[3:0]];
  assign array_index_75886 = array_update_75883[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_75890 = smul32b_32b_x_32b(array_index_74726[add_75882 > 32'h0000_0009 ? 4'h9 : add_75882[3:0]], array_index_75885[add_75802 > 32'h0000_0009 ? 4'h9 : add_75802[3:0]]);
  assign add_75892 = array_index_75886[add_75802 > 32'h0000_0009 ? 4'h9 : add_75802[3:0]] + smul_75890;
  assign array_update_75894[0] = add_75802 == 32'h0000_0000 ? add_75892 : array_index_75886[0];
  assign array_update_75894[1] = add_75802 == 32'h0000_0001 ? add_75892 : array_index_75886[1];
  assign array_update_75894[2] = add_75802 == 32'h0000_0002 ? add_75892 : array_index_75886[2];
  assign array_update_75894[3] = add_75802 == 32'h0000_0003 ? add_75892 : array_index_75886[3];
  assign array_update_75894[4] = add_75802 == 32'h0000_0004 ? add_75892 : array_index_75886[4];
  assign array_update_75894[5] = add_75802 == 32'h0000_0005 ? add_75892 : array_index_75886[5];
  assign array_update_75894[6] = add_75802 == 32'h0000_0006 ? add_75892 : array_index_75886[6];
  assign array_update_75894[7] = add_75802 == 32'h0000_0007 ? add_75892 : array_index_75886[7];
  assign array_update_75894[8] = add_75802 == 32'h0000_0008 ? add_75892 : array_index_75886[8];
  assign array_update_75894[9] = add_75802 == 32'h0000_0009 ? add_75892 : array_index_75886[9];
  assign add_75895 = add_75882 + 32'h0000_0001;
  assign array_update_75896[0] = add_74719 == 32'h0000_0000 ? array_update_75894 : array_update_75883[0];
  assign array_update_75896[1] = add_74719 == 32'h0000_0001 ? array_update_75894 : array_update_75883[1];
  assign array_update_75896[2] = add_74719 == 32'h0000_0002 ? array_update_75894 : array_update_75883[2];
  assign array_update_75896[3] = add_74719 == 32'h0000_0003 ? array_update_75894 : array_update_75883[3];
  assign array_update_75896[4] = add_74719 == 32'h0000_0004 ? array_update_75894 : array_update_75883[4];
  assign array_update_75896[5] = add_74719 == 32'h0000_0005 ? array_update_75894 : array_update_75883[5];
  assign array_update_75896[6] = add_74719 == 32'h0000_0006 ? array_update_75894 : array_update_75883[6];
  assign array_update_75896[7] = add_74719 == 32'h0000_0007 ? array_update_75894 : array_update_75883[7];
  assign array_update_75896[8] = add_74719 == 32'h0000_0008 ? array_update_75894 : array_update_75883[8];
  assign array_update_75896[9] = add_74719 == 32'h0000_0009 ? array_update_75894 : array_update_75883[9];
  assign array_index_75898 = array_update_72021[add_75895 > 32'h0000_0009 ? 4'h9 : add_75895[3:0]];
  assign array_index_75899 = array_update_75896[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_75903 = smul32b_32b_x_32b(array_index_74726[add_75895 > 32'h0000_0009 ? 4'h9 : add_75895[3:0]], array_index_75898[add_75802 > 32'h0000_0009 ? 4'h9 : add_75802[3:0]]);
  assign add_75905 = array_index_75899[add_75802 > 32'h0000_0009 ? 4'h9 : add_75802[3:0]] + smul_75903;
  assign array_update_75907[0] = add_75802 == 32'h0000_0000 ? add_75905 : array_index_75899[0];
  assign array_update_75907[1] = add_75802 == 32'h0000_0001 ? add_75905 : array_index_75899[1];
  assign array_update_75907[2] = add_75802 == 32'h0000_0002 ? add_75905 : array_index_75899[2];
  assign array_update_75907[3] = add_75802 == 32'h0000_0003 ? add_75905 : array_index_75899[3];
  assign array_update_75907[4] = add_75802 == 32'h0000_0004 ? add_75905 : array_index_75899[4];
  assign array_update_75907[5] = add_75802 == 32'h0000_0005 ? add_75905 : array_index_75899[5];
  assign array_update_75907[6] = add_75802 == 32'h0000_0006 ? add_75905 : array_index_75899[6];
  assign array_update_75907[7] = add_75802 == 32'h0000_0007 ? add_75905 : array_index_75899[7];
  assign array_update_75907[8] = add_75802 == 32'h0000_0008 ? add_75905 : array_index_75899[8];
  assign array_update_75907[9] = add_75802 == 32'h0000_0009 ? add_75905 : array_index_75899[9];
  assign add_75908 = add_75895 + 32'h0000_0001;
  assign array_update_75909[0] = add_74719 == 32'h0000_0000 ? array_update_75907 : array_update_75896[0];
  assign array_update_75909[1] = add_74719 == 32'h0000_0001 ? array_update_75907 : array_update_75896[1];
  assign array_update_75909[2] = add_74719 == 32'h0000_0002 ? array_update_75907 : array_update_75896[2];
  assign array_update_75909[3] = add_74719 == 32'h0000_0003 ? array_update_75907 : array_update_75896[3];
  assign array_update_75909[4] = add_74719 == 32'h0000_0004 ? array_update_75907 : array_update_75896[4];
  assign array_update_75909[5] = add_74719 == 32'h0000_0005 ? array_update_75907 : array_update_75896[5];
  assign array_update_75909[6] = add_74719 == 32'h0000_0006 ? array_update_75907 : array_update_75896[6];
  assign array_update_75909[7] = add_74719 == 32'h0000_0007 ? array_update_75907 : array_update_75896[7];
  assign array_update_75909[8] = add_74719 == 32'h0000_0008 ? array_update_75907 : array_update_75896[8];
  assign array_update_75909[9] = add_74719 == 32'h0000_0009 ? array_update_75907 : array_update_75896[9];
  assign array_index_75911 = array_update_72021[add_75908 > 32'h0000_0009 ? 4'h9 : add_75908[3:0]];
  assign array_index_75912 = array_update_75909[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_75916 = smul32b_32b_x_32b(array_index_74726[add_75908 > 32'h0000_0009 ? 4'h9 : add_75908[3:0]], array_index_75911[add_75802 > 32'h0000_0009 ? 4'h9 : add_75802[3:0]]);
  assign add_75918 = array_index_75912[add_75802 > 32'h0000_0009 ? 4'h9 : add_75802[3:0]] + smul_75916;
  assign array_update_75920[0] = add_75802 == 32'h0000_0000 ? add_75918 : array_index_75912[0];
  assign array_update_75920[1] = add_75802 == 32'h0000_0001 ? add_75918 : array_index_75912[1];
  assign array_update_75920[2] = add_75802 == 32'h0000_0002 ? add_75918 : array_index_75912[2];
  assign array_update_75920[3] = add_75802 == 32'h0000_0003 ? add_75918 : array_index_75912[3];
  assign array_update_75920[4] = add_75802 == 32'h0000_0004 ? add_75918 : array_index_75912[4];
  assign array_update_75920[5] = add_75802 == 32'h0000_0005 ? add_75918 : array_index_75912[5];
  assign array_update_75920[6] = add_75802 == 32'h0000_0006 ? add_75918 : array_index_75912[6];
  assign array_update_75920[7] = add_75802 == 32'h0000_0007 ? add_75918 : array_index_75912[7];
  assign array_update_75920[8] = add_75802 == 32'h0000_0008 ? add_75918 : array_index_75912[8];
  assign array_update_75920[9] = add_75802 == 32'h0000_0009 ? add_75918 : array_index_75912[9];
  assign add_75921 = add_75908 + 32'h0000_0001;
  assign array_update_75922[0] = add_74719 == 32'h0000_0000 ? array_update_75920 : array_update_75909[0];
  assign array_update_75922[1] = add_74719 == 32'h0000_0001 ? array_update_75920 : array_update_75909[1];
  assign array_update_75922[2] = add_74719 == 32'h0000_0002 ? array_update_75920 : array_update_75909[2];
  assign array_update_75922[3] = add_74719 == 32'h0000_0003 ? array_update_75920 : array_update_75909[3];
  assign array_update_75922[4] = add_74719 == 32'h0000_0004 ? array_update_75920 : array_update_75909[4];
  assign array_update_75922[5] = add_74719 == 32'h0000_0005 ? array_update_75920 : array_update_75909[5];
  assign array_update_75922[6] = add_74719 == 32'h0000_0006 ? array_update_75920 : array_update_75909[6];
  assign array_update_75922[7] = add_74719 == 32'h0000_0007 ? array_update_75920 : array_update_75909[7];
  assign array_update_75922[8] = add_74719 == 32'h0000_0008 ? array_update_75920 : array_update_75909[8];
  assign array_update_75922[9] = add_74719 == 32'h0000_0009 ? array_update_75920 : array_update_75909[9];
  assign array_index_75924 = array_update_72021[add_75921 > 32'h0000_0009 ? 4'h9 : add_75921[3:0]];
  assign array_index_75925 = array_update_75922[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_75929 = smul32b_32b_x_32b(array_index_74726[add_75921 > 32'h0000_0009 ? 4'h9 : add_75921[3:0]], array_index_75924[add_75802 > 32'h0000_0009 ? 4'h9 : add_75802[3:0]]);
  assign add_75931 = array_index_75925[add_75802 > 32'h0000_0009 ? 4'h9 : add_75802[3:0]] + smul_75929;
  assign array_update_75932[0] = add_75802 == 32'h0000_0000 ? add_75931 : array_index_75925[0];
  assign array_update_75932[1] = add_75802 == 32'h0000_0001 ? add_75931 : array_index_75925[1];
  assign array_update_75932[2] = add_75802 == 32'h0000_0002 ? add_75931 : array_index_75925[2];
  assign array_update_75932[3] = add_75802 == 32'h0000_0003 ? add_75931 : array_index_75925[3];
  assign array_update_75932[4] = add_75802 == 32'h0000_0004 ? add_75931 : array_index_75925[4];
  assign array_update_75932[5] = add_75802 == 32'h0000_0005 ? add_75931 : array_index_75925[5];
  assign array_update_75932[6] = add_75802 == 32'h0000_0006 ? add_75931 : array_index_75925[6];
  assign array_update_75932[7] = add_75802 == 32'h0000_0007 ? add_75931 : array_index_75925[7];
  assign array_update_75932[8] = add_75802 == 32'h0000_0008 ? add_75931 : array_index_75925[8];
  assign array_update_75932[9] = add_75802 == 32'h0000_0009 ? add_75931 : array_index_75925[9];
  assign array_update_75933[0] = add_74719 == 32'h0000_0000 ? array_update_75932 : array_update_75922[0];
  assign array_update_75933[1] = add_74719 == 32'h0000_0001 ? array_update_75932 : array_update_75922[1];
  assign array_update_75933[2] = add_74719 == 32'h0000_0002 ? array_update_75932 : array_update_75922[2];
  assign array_update_75933[3] = add_74719 == 32'h0000_0003 ? array_update_75932 : array_update_75922[3];
  assign array_update_75933[4] = add_74719 == 32'h0000_0004 ? array_update_75932 : array_update_75922[4];
  assign array_update_75933[5] = add_74719 == 32'h0000_0005 ? array_update_75932 : array_update_75922[5];
  assign array_update_75933[6] = add_74719 == 32'h0000_0006 ? array_update_75932 : array_update_75922[6];
  assign array_update_75933[7] = add_74719 == 32'h0000_0007 ? array_update_75932 : array_update_75922[7];
  assign array_update_75933[8] = add_74719 == 32'h0000_0008 ? array_update_75932 : array_update_75922[8];
  assign array_update_75933[9] = add_74719 == 32'h0000_0009 ? array_update_75932 : array_update_75922[9];
  assign array_index_75935 = array_update_75933[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign add_75937 = add_75802 + 32'h0000_0001;
  assign array_update_75938[0] = add_75937 == 32'h0000_0000 ? 32'h0000_0000 : array_index_75935[0];
  assign array_update_75938[1] = add_75937 == 32'h0000_0001 ? 32'h0000_0000 : array_index_75935[1];
  assign array_update_75938[2] = add_75937 == 32'h0000_0002 ? 32'h0000_0000 : array_index_75935[2];
  assign array_update_75938[3] = add_75937 == 32'h0000_0003 ? 32'h0000_0000 : array_index_75935[3];
  assign array_update_75938[4] = add_75937 == 32'h0000_0004 ? 32'h0000_0000 : array_index_75935[4];
  assign array_update_75938[5] = add_75937 == 32'h0000_0005 ? 32'h0000_0000 : array_index_75935[5];
  assign array_update_75938[6] = add_75937 == 32'h0000_0006 ? 32'h0000_0000 : array_index_75935[6];
  assign array_update_75938[7] = add_75937 == 32'h0000_0007 ? 32'h0000_0000 : array_index_75935[7];
  assign array_update_75938[8] = add_75937 == 32'h0000_0008 ? 32'h0000_0000 : array_index_75935[8];
  assign array_update_75938[9] = add_75937 == 32'h0000_0009 ? 32'h0000_0000 : array_index_75935[9];
  assign literal_75939 = 32'h0000_0000;
  assign array_update_75940[0] = add_74719 == 32'h0000_0000 ? array_update_75938 : array_update_75933[0];
  assign array_update_75940[1] = add_74719 == 32'h0000_0001 ? array_update_75938 : array_update_75933[1];
  assign array_update_75940[2] = add_74719 == 32'h0000_0002 ? array_update_75938 : array_update_75933[2];
  assign array_update_75940[3] = add_74719 == 32'h0000_0003 ? array_update_75938 : array_update_75933[3];
  assign array_update_75940[4] = add_74719 == 32'h0000_0004 ? array_update_75938 : array_update_75933[4];
  assign array_update_75940[5] = add_74719 == 32'h0000_0005 ? array_update_75938 : array_update_75933[5];
  assign array_update_75940[6] = add_74719 == 32'h0000_0006 ? array_update_75938 : array_update_75933[6];
  assign array_update_75940[7] = add_74719 == 32'h0000_0007 ? array_update_75938 : array_update_75933[7];
  assign array_update_75940[8] = add_74719 == 32'h0000_0008 ? array_update_75938 : array_update_75933[8];
  assign array_update_75940[9] = add_74719 == 32'h0000_0009 ? array_update_75938 : array_update_75933[9];
  assign array_index_75942 = array_update_72021[literal_75939 > 32'h0000_0009 ? 4'h9 : literal_75939[3:0]];
  assign array_index_75943 = array_update_75940[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_75947 = smul32b_32b_x_32b(array_index_74726[literal_75939 > 32'h0000_0009 ? 4'h9 : literal_75939[3:0]], array_index_75942[add_75937 > 32'h0000_0009 ? 4'h9 : add_75937[3:0]]);
  assign add_75949 = array_index_75943[add_75937 > 32'h0000_0009 ? 4'h9 : add_75937[3:0]] + smul_75947;
  assign array_update_75951[0] = add_75937 == 32'h0000_0000 ? add_75949 : array_index_75943[0];
  assign array_update_75951[1] = add_75937 == 32'h0000_0001 ? add_75949 : array_index_75943[1];
  assign array_update_75951[2] = add_75937 == 32'h0000_0002 ? add_75949 : array_index_75943[2];
  assign array_update_75951[3] = add_75937 == 32'h0000_0003 ? add_75949 : array_index_75943[3];
  assign array_update_75951[4] = add_75937 == 32'h0000_0004 ? add_75949 : array_index_75943[4];
  assign array_update_75951[5] = add_75937 == 32'h0000_0005 ? add_75949 : array_index_75943[5];
  assign array_update_75951[6] = add_75937 == 32'h0000_0006 ? add_75949 : array_index_75943[6];
  assign array_update_75951[7] = add_75937 == 32'h0000_0007 ? add_75949 : array_index_75943[7];
  assign array_update_75951[8] = add_75937 == 32'h0000_0008 ? add_75949 : array_index_75943[8];
  assign array_update_75951[9] = add_75937 == 32'h0000_0009 ? add_75949 : array_index_75943[9];
  assign add_75952 = literal_75939 + 32'h0000_0001;
  assign array_update_75953[0] = add_74719 == 32'h0000_0000 ? array_update_75951 : array_update_75940[0];
  assign array_update_75953[1] = add_74719 == 32'h0000_0001 ? array_update_75951 : array_update_75940[1];
  assign array_update_75953[2] = add_74719 == 32'h0000_0002 ? array_update_75951 : array_update_75940[2];
  assign array_update_75953[3] = add_74719 == 32'h0000_0003 ? array_update_75951 : array_update_75940[3];
  assign array_update_75953[4] = add_74719 == 32'h0000_0004 ? array_update_75951 : array_update_75940[4];
  assign array_update_75953[5] = add_74719 == 32'h0000_0005 ? array_update_75951 : array_update_75940[5];
  assign array_update_75953[6] = add_74719 == 32'h0000_0006 ? array_update_75951 : array_update_75940[6];
  assign array_update_75953[7] = add_74719 == 32'h0000_0007 ? array_update_75951 : array_update_75940[7];
  assign array_update_75953[8] = add_74719 == 32'h0000_0008 ? array_update_75951 : array_update_75940[8];
  assign array_update_75953[9] = add_74719 == 32'h0000_0009 ? array_update_75951 : array_update_75940[9];
  assign array_index_75955 = array_update_72021[add_75952 > 32'h0000_0009 ? 4'h9 : add_75952[3:0]];
  assign array_index_75956 = array_update_75953[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_75960 = smul32b_32b_x_32b(array_index_74726[add_75952 > 32'h0000_0009 ? 4'h9 : add_75952[3:0]], array_index_75955[add_75937 > 32'h0000_0009 ? 4'h9 : add_75937[3:0]]);
  assign add_75962 = array_index_75956[add_75937 > 32'h0000_0009 ? 4'h9 : add_75937[3:0]] + smul_75960;
  assign array_update_75964[0] = add_75937 == 32'h0000_0000 ? add_75962 : array_index_75956[0];
  assign array_update_75964[1] = add_75937 == 32'h0000_0001 ? add_75962 : array_index_75956[1];
  assign array_update_75964[2] = add_75937 == 32'h0000_0002 ? add_75962 : array_index_75956[2];
  assign array_update_75964[3] = add_75937 == 32'h0000_0003 ? add_75962 : array_index_75956[3];
  assign array_update_75964[4] = add_75937 == 32'h0000_0004 ? add_75962 : array_index_75956[4];
  assign array_update_75964[5] = add_75937 == 32'h0000_0005 ? add_75962 : array_index_75956[5];
  assign array_update_75964[6] = add_75937 == 32'h0000_0006 ? add_75962 : array_index_75956[6];
  assign array_update_75964[7] = add_75937 == 32'h0000_0007 ? add_75962 : array_index_75956[7];
  assign array_update_75964[8] = add_75937 == 32'h0000_0008 ? add_75962 : array_index_75956[8];
  assign array_update_75964[9] = add_75937 == 32'h0000_0009 ? add_75962 : array_index_75956[9];
  assign add_75965 = add_75952 + 32'h0000_0001;
  assign array_update_75966[0] = add_74719 == 32'h0000_0000 ? array_update_75964 : array_update_75953[0];
  assign array_update_75966[1] = add_74719 == 32'h0000_0001 ? array_update_75964 : array_update_75953[1];
  assign array_update_75966[2] = add_74719 == 32'h0000_0002 ? array_update_75964 : array_update_75953[2];
  assign array_update_75966[3] = add_74719 == 32'h0000_0003 ? array_update_75964 : array_update_75953[3];
  assign array_update_75966[4] = add_74719 == 32'h0000_0004 ? array_update_75964 : array_update_75953[4];
  assign array_update_75966[5] = add_74719 == 32'h0000_0005 ? array_update_75964 : array_update_75953[5];
  assign array_update_75966[6] = add_74719 == 32'h0000_0006 ? array_update_75964 : array_update_75953[6];
  assign array_update_75966[7] = add_74719 == 32'h0000_0007 ? array_update_75964 : array_update_75953[7];
  assign array_update_75966[8] = add_74719 == 32'h0000_0008 ? array_update_75964 : array_update_75953[8];
  assign array_update_75966[9] = add_74719 == 32'h0000_0009 ? array_update_75964 : array_update_75953[9];
  assign array_index_75968 = array_update_72021[add_75965 > 32'h0000_0009 ? 4'h9 : add_75965[3:0]];
  assign array_index_75969 = array_update_75966[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_75973 = smul32b_32b_x_32b(array_index_74726[add_75965 > 32'h0000_0009 ? 4'h9 : add_75965[3:0]], array_index_75968[add_75937 > 32'h0000_0009 ? 4'h9 : add_75937[3:0]]);
  assign add_75975 = array_index_75969[add_75937 > 32'h0000_0009 ? 4'h9 : add_75937[3:0]] + smul_75973;
  assign array_update_75977[0] = add_75937 == 32'h0000_0000 ? add_75975 : array_index_75969[0];
  assign array_update_75977[1] = add_75937 == 32'h0000_0001 ? add_75975 : array_index_75969[1];
  assign array_update_75977[2] = add_75937 == 32'h0000_0002 ? add_75975 : array_index_75969[2];
  assign array_update_75977[3] = add_75937 == 32'h0000_0003 ? add_75975 : array_index_75969[3];
  assign array_update_75977[4] = add_75937 == 32'h0000_0004 ? add_75975 : array_index_75969[4];
  assign array_update_75977[5] = add_75937 == 32'h0000_0005 ? add_75975 : array_index_75969[5];
  assign array_update_75977[6] = add_75937 == 32'h0000_0006 ? add_75975 : array_index_75969[6];
  assign array_update_75977[7] = add_75937 == 32'h0000_0007 ? add_75975 : array_index_75969[7];
  assign array_update_75977[8] = add_75937 == 32'h0000_0008 ? add_75975 : array_index_75969[8];
  assign array_update_75977[9] = add_75937 == 32'h0000_0009 ? add_75975 : array_index_75969[9];
  assign add_75978 = add_75965 + 32'h0000_0001;
  assign array_update_75979[0] = add_74719 == 32'h0000_0000 ? array_update_75977 : array_update_75966[0];
  assign array_update_75979[1] = add_74719 == 32'h0000_0001 ? array_update_75977 : array_update_75966[1];
  assign array_update_75979[2] = add_74719 == 32'h0000_0002 ? array_update_75977 : array_update_75966[2];
  assign array_update_75979[3] = add_74719 == 32'h0000_0003 ? array_update_75977 : array_update_75966[3];
  assign array_update_75979[4] = add_74719 == 32'h0000_0004 ? array_update_75977 : array_update_75966[4];
  assign array_update_75979[5] = add_74719 == 32'h0000_0005 ? array_update_75977 : array_update_75966[5];
  assign array_update_75979[6] = add_74719 == 32'h0000_0006 ? array_update_75977 : array_update_75966[6];
  assign array_update_75979[7] = add_74719 == 32'h0000_0007 ? array_update_75977 : array_update_75966[7];
  assign array_update_75979[8] = add_74719 == 32'h0000_0008 ? array_update_75977 : array_update_75966[8];
  assign array_update_75979[9] = add_74719 == 32'h0000_0009 ? array_update_75977 : array_update_75966[9];
  assign array_index_75981 = array_update_72021[add_75978 > 32'h0000_0009 ? 4'h9 : add_75978[3:0]];
  assign array_index_75982 = array_update_75979[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_75986 = smul32b_32b_x_32b(array_index_74726[add_75978 > 32'h0000_0009 ? 4'h9 : add_75978[3:0]], array_index_75981[add_75937 > 32'h0000_0009 ? 4'h9 : add_75937[3:0]]);
  assign add_75988 = array_index_75982[add_75937 > 32'h0000_0009 ? 4'h9 : add_75937[3:0]] + smul_75986;
  assign array_update_75990[0] = add_75937 == 32'h0000_0000 ? add_75988 : array_index_75982[0];
  assign array_update_75990[1] = add_75937 == 32'h0000_0001 ? add_75988 : array_index_75982[1];
  assign array_update_75990[2] = add_75937 == 32'h0000_0002 ? add_75988 : array_index_75982[2];
  assign array_update_75990[3] = add_75937 == 32'h0000_0003 ? add_75988 : array_index_75982[3];
  assign array_update_75990[4] = add_75937 == 32'h0000_0004 ? add_75988 : array_index_75982[4];
  assign array_update_75990[5] = add_75937 == 32'h0000_0005 ? add_75988 : array_index_75982[5];
  assign array_update_75990[6] = add_75937 == 32'h0000_0006 ? add_75988 : array_index_75982[6];
  assign array_update_75990[7] = add_75937 == 32'h0000_0007 ? add_75988 : array_index_75982[7];
  assign array_update_75990[8] = add_75937 == 32'h0000_0008 ? add_75988 : array_index_75982[8];
  assign array_update_75990[9] = add_75937 == 32'h0000_0009 ? add_75988 : array_index_75982[9];
  assign add_75991 = add_75978 + 32'h0000_0001;
  assign array_update_75992[0] = add_74719 == 32'h0000_0000 ? array_update_75990 : array_update_75979[0];
  assign array_update_75992[1] = add_74719 == 32'h0000_0001 ? array_update_75990 : array_update_75979[1];
  assign array_update_75992[2] = add_74719 == 32'h0000_0002 ? array_update_75990 : array_update_75979[2];
  assign array_update_75992[3] = add_74719 == 32'h0000_0003 ? array_update_75990 : array_update_75979[3];
  assign array_update_75992[4] = add_74719 == 32'h0000_0004 ? array_update_75990 : array_update_75979[4];
  assign array_update_75992[5] = add_74719 == 32'h0000_0005 ? array_update_75990 : array_update_75979[5];
  assign array_update_75992[6] = add_74719 == 32'h0000_0006 ? array_update_75990 : array_update_75979[6];
  assign array_update_75992[7] = add_74719 == 32'h0000_0007 ? array_update_75990 : array_update_75979[7];
  assign array_update_75992[8] = add_74719 == 32'h0000_0008 ? array_update_75990 : array_update_75979[8];
  assign array_update_75992[9] = add_74719 == 32'h0000_0009 ? array_update_75990 : array_update_75979[9];
  assign array_index_75994 = array_update_72021[add_75991 > 32'h0000_0009 ? 4'h9 : add_75991[3:0]];
  assign array_index_75995 = array_update_75992[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_75999 = smul32b_32b_x_32b(array_index_74726[add_75991 > 32'h0000_0009 ? 4'h9 : add_75991[3:0]], array_index_75994[add_75937 > 32'h0000_0009 ? 4'h9 : add_75937[3:0]]);
  assign add_76001 = array_index_75995[add_75937 > 32'h0000_0009 ? 4'h9 : add_75937[3:0]] + smul_75999;
  assign array_update_76003[0] = add_75937 == 32'h0000_0000 ? add_76001 : array_index_75995[0];
  assign array_update_76003[1] = add_75937 == 32'h0000_0001 ? add_76001 : array_index_75995[1];
  assign array_update_76003[2] = add_75937 == 32'h0000_0002 ? add_76001 : array_index_75995[2];
  assign array_update_76003[3] = add_75937 == 32'h0000_0003 ? add_76001 : array_index_75995[3];
  assign array_update_76003[4] = add_75937 == 32'h0000_0004 ? add_76001 : array_index_75995[4];
  assign array_update_76003[5] = add_75937 == 32'h0000_0005 ? add_76001 : array_index_75995[5];
  assign array_update_76003[6] = add_75937 == 32'h0000_0006 ? add_76001 : array_index_75995[6];
  assign array_update_76003[7] = add_75937 == 32'h0000_0007 ? add_76001 : array_index_75995[7];
  assign array_update_76003[8] = add_75937 == 32'h0000_0008 ? add_76001 : array_index_75995[8];
  assign array_update_76003[9] = add_75937 == 32'h0000_0009 ? add_76001 : array_index_75995[9];
  assign add_76004 = add_75991 + 32'h0000_0001;
  assign array_update_76005[0] = add_74719 == 32'h0000_0000 ? array_update_76003 : array_update_75992[0];
  assign array_update_76005[1] = add_74719 == 32'h0000_0001 ? array_update_76003 : array_update_75992[1];
  assign array_update_76005[2] = add_74719 == 32'h0000_0002 ? array_update_76003 : array_update_75992[2];
  assign array_update_76005[3] = add_74719 == 32'h0000_0003 ? array_update_76003 : array_update_75992[3];
  assign array_update_76005[4] = add_74719 == 32'h0000_0004 ? array_update_76003 : array_update_75992[4];
  assign array_update_76005[5] = add_74719 == 32'h0000_0005 ? array_update_76003 : array_update_75992[5];
  assign array_update_76005[6] = add_74719 == 32'h0000_0006 ? array_update_76003 : array_update_75992[6];
  assign array_update_76005[7] = add_74719 == 32'h0000_0007 ? array_update_76003 : array_update_75992[7];
  assign array_update_76005[8] = add_74719 == 32'h0000_0008 ? array_update_76003 : array_update_75992[8];
  assign array_update_76005[9] = add_74719 == 32'h0000_0009 ? array_update_76003 : array_update_75992[9];
  assign array_index_76007 = array_update_72021[add_76004 > 32'h0000_0009 ? 4'h9 : add_76004[3:0]];
  assign array_index_76008 = array_update_76005[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_76012 = smul32b_32b_x_32b(array_index_74726[add_76004 > 32'h0000_0009 ? 4'h9 : add_76004[3:0]], array_index_76007[add_75937 > 32'h0000_0009 ? 4'h9 : add_75937[3:0]]);
  assign add_76014 = array_index_76008[add_75937 > 32'h0000_0009 ? 4'h9 : add_75937[3:0]] + smul_76012;
  assign array_update_76016[0] = add_75937 == 32'h0000_0000 ? add_76014 : array_index_76008[0];
  assign array_update_76016[1] = add_75937 == 32'h0000_0001 ? add_76014 : array_index_76008[1];
  assign array_update_76016[2] = add_75937 == 32'h0000_0002 ? add_76014 : array_index_76008[2];
  assign array_update_76016[3] = add_75937 == 32'h0000_0003 ? add_76014 : array_index_76008[3];
  assign array_update_76016[4] = add_75937 == 32'h0000_0004 ? add_76014 : array_index_76008[4];
  assign array_update_76016[5] = add_75937 == 32'h0000_0005 ? add_76014 : array_index_76008[5];
  assign array_update_76016[6] = add_75937 == 32'h0000_0006 ? add_76014 : array_index_76008[6];
  assign array_update_76016[7] = add_75937 == 32'h0000_0007 ? add_76014 : array_index_76008[7];
  assign array_update_76016[8] = add_75937 == 32'h0000_0008 ? add_76014 : array_index_76008[8];
  assign array_update_76016[9] = add_75937 == 32'h0000_0009 ? add_76014 : array_index_76008[9];
  assign add_76017 = add_76004 + 32'h0000_0001;
  assign array_update_76018[0] = add_74719 == 32'h0000_0000 ? array_update_76016 : array_update_76005[0];
  assign array_update_76018[1] = add_74719 == 32'h0000_0001 ? array_update_76016 : array_update_76005[1];
  assign array_update_76018[2] = add_74719 == 32'h0000_0002 ? array_update_76016 : array_update_76005[2];
  assign array_update_76018[3] = add_74719 == 32'h0000_0003 ? array_update_76016 : array_update_76005[3];
  assign array_update_76018[4] = add_74719 == 32'h0000_0004 ? array_update_76016 : array_update_76005[4];
  assign array_update_76018[5] = add_74719 == 32'h0000_0005 ? array_update_76016 : array_update_76005[5];
  assign array_update_76018[6] = add_74719 == 32'h0000_0006 ? array_update_76016 : array_update_76005[6];
  assign array_update_76018[7] = add_74719 == 32'h0000_0007 ? array_update_76016 : array_update_76005[7];
  assign array_update_76018[8] = add_74719 == 32'h0000_0008 ? array_update_76016 : array_update_76005[8];
  assign array_update_76018[9] = add_74719 == 32'h0000_0009 ? array_update_76016 : array_update_76005[9];
  assign array_index_76020 = array_update_72021[add_76017 > 32'h0000_0009 ? 4'h9 : add_76017[3:0]];
  assign array_index_76021 = array_update_76018[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_76025 = smul32b_32b_x_32b(array_index_74726[add_76017 > 32'h0000_0009 ? 4'h9 : add_76017[3:0]], array_index_76020[add_75937 > 32'h0000_0009 ? 4'h9 : add_75937[3:0]]);
  assign add_76027 = array_index_76021[add_75937 > 32'h0000_0009 ? 4'h9 : add_75937[3:0]] + smul_76025;
  assign array_update_76029[0] = add_75937 == 32'h0000_0000 ? add_76027 : array_index_76021[0];
  assign array_update_76029[1] = add_75937 == 32'h0000_0001 ? add_76027 : array_index_76021[1];
  assign array_update_76029[2] = add_75937 == 32'h0000_0002 ? add_76027 : array_index_76021[2];
  assign array_update_76029[3] = add_75937 == 32'h0000_0003 ? add_76027 : array_index_76021[3];
  assign array_update_76029[4] = add_75937 == 32'h0000_0004 ? add_76027 : array_index_76021[4];
  assign array_update_76029[5] = add_75937 == 32'h0000_0005 ? add_76027 : array_index_76021[5];
  assign array_update_76029[6] = add_75937 == 32'h0000_0006 ? add_76027 : array_index_76021[6];
  assign array_update_76029[7] = add_75937 == 32'h0000_0007 ? add_76027 : array_index_76021[7];
  assign array_update_76029[8] = add_75937 == 32'h0000_0008 ? add_76027 : array_index_76021[8];
  assign array_update_76029[9] = add_75937 == 32'h0000_0009 ? add_76027 : array_index_76021[9];
  assign add_76030 = add_76017 + 32'h0000_0001;
  assign array_update_76031[0] = add_74719 == 32'h0000_0000 ? array_update_76029 : array_update_76018[0];
  assign array_update_76031[1] = add_74719 == 32'h0000_0001 ? array_update_76029 : array_update_76018[1];
  assign array_update_76031[2] = add_74719 == 32'h0000_0002 ? array_update_76029 : array_update_76018[2];
  assign array_update_76031[3] = add_74719 == 32'h0000_0003 ? array_update_76029 : array_update_76018[3];
  assign array_update_76031[4] = add_74719 == 32'h0000_0004 ? array_update_76029 : array_update_76018[4];
  assign array_update_76031[5] = add_74719 == 32'h0000_0005 ? array_update_76029 : array_update_76018[5];
  assign array_update_76031[6] = add_74719 == 32'h0000_0006 ? array_update_76029 : array_update_76018[6];
  assign array_update_76031[7] = add_74719 == 32'h0000_0007 ? array_update_76029 : array_update_76018[7];
  assign array_update_76031[8] = add_74719 == 32'h0000_0008 ? array_update_76029 : array_update_76018[8];
  assign array_update_76031[9] = add_74719 == 32'h0000_0009 ? array_update_76029 : array_update_76018[9];
  assign array_index_76033 = array_update_72021[add_76030 > 32'h0000_0009 ? 4'h9 : add_76030[3:0]];
  assign array_index_76034 = array_update_76031[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_76038 = smul32b_32b_x_32b(array_index_74726[add_76030 > 32'h0000_0009 ? 4'h9 : add_76030[3:0]], array_index_76033[add_75937 > 32'h0000_0009 ? 4'h9 : add_75937[3:0]]);
  assign add_76040 = array_index_76034[add_75937 > 32'h0000_0009 ? 4'h9 : add_75937[3:0]] + smul_76038;
  assign array_update_76042[0] = add_75937 == 32'h0000_0000 ? add_76040 : array_index_76034[0];
  assign array_update_76042[1] = add_75937 == 32'h0000_0001 ? add_76040 : array_index_76034[1];
  assign array_update_76042[2] = add_75937 == 32'h0000_0002 ? add_76040 : array_index_76034[2];
  assign array_update_76042[3] = add_75937 == 32'h0000_0003 ? add_76040 : array_index_76034[3];
  assign array_update_76042[4] = add_75937 == 32'h0000_0004 ? add_76040 : array_index_76034[4];
  assign array_update_76042[5] = add_75937 == 32'h0000_0005 ? add_76040 : array_index_76034[5];
  assign array_update_76042[6] = add_75937 == 32'h0000_0006 ? add_76040 : array_index_76034[6];
  assign array_update_76042[7] = add_75937 == 32'h0000_0007 ? add_76040 : array_index_76034[7];
  assign array_update_76042[8] = add_75937 == 32'h0000_0008 ? add_76040 : array_index_76034[8];
  assign array_update_76042[9] = add_75937 == 32'h0000_0009 ? add_76040 : array_index_76034[9];
  assign add_76043 = add_76030 + 32'h0000_0001;
  assign array_update_76044[0] = add_74719 == 32'h0000_0000 ? array_update_76042 : array_update_76031[0];
  assign array_update_76044[1] = add_74719 == 32'h0000_0001 ? array_update_76042 : array_update_76031[1];
  assign array_update_76044[2] = add_74719 == 32'h0000_0002 ? array_update_76042 : array_update_76031[2];
  assign array_update_76044[3] = add_74719 == 32'h0000_0003 ? array_update_76042 : array_update_76031[3];
  assign array_update_76044[4] = add_74719 == 32'h0000_0004 ? array_update_76042 : array_update_76031[4];
  assign array_update_76044[5] = add_74719 == 32'h0000_0005 ? array_update_76042 : array_update_76031[5];
  assign array_update_76044[6] = add_74719 == 32'h0000_0006 ? array_update_76042 : array_update_76031[6];
  assign array_update_76044[7] = add_74719 == 32'h0000_0007 ? array_update_76042 : array_update_76031[7];
  assign array_update_76044[8] = add_74719 == 32'h0000_0008 ? array_update_76042 : array_update_76031[8];
  assign array_update_76044[9] = add_74719 == 32'h0000_0009 ? array_update_76042 : array_update_76031[9];
  assign array_index_76046 = array_update_72021[add_76043 > 32'h0000_0009 ? 4'h9 : add_76043[3:0]];
  assign array_index_76047 = array_update_76044[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_76051 = smul32b_32b_x_32b(array_index_74726[add_76043 > 32'h0000_0009 ? 4'h9 : add_76043[3:0]], array_index_76046[add_75937 > 32'h0000_0009 ? 4'h9 : add_75937[3:0]]);
  assign add_76053 = array_index_76047[add_75937 > 32'h0000_0009 ? 4'h9 : add_75937[3:0]] + smul_76051;
  assign array_update_76055[0] = add_75937 == 32'h0000_0000 ? add_76053 : array_index_76047[0];
  assign array_update_76055[1] = add_75937 == 32'h0000_0001 ? add_76053 : array_index_76047[1];
  assign array_update_76055[2] = add_75937 == 32'h0000_0002 ? add_76053 : array_index_76047[2];
  assign array_update_76055[3] = add_75937 == 32'h0000_0003 ? add_76053 : array_index_76047[3];
  assign array_update_76055[4] = add_75937 == 32'h0000_0004 ? add_76053 : array_index_76047[4];
  assign array_update_76055[5] = add_75937 == 32'h0000_0005 ? add_76053 : array_index_76047[5];
  assign array_update_76055[6] = add_75937 == 32'h0000_0006 ? add_76053 : array_index_76047[6];
  assign array_update_76055[7] = add_75937 == 32'h0000_0007 ? add_76053 : array_index_76047[7];
  assign array_update_76055[8] = add_75937 == 32'h0000_0008 ? add_76053 : array_index_76047[8];
  assign array_update_76055[9] = add_75937 == 32'h0000_0009 ? add_76053 : array_index_76047[9];
  assign add_76056 = add_76043 + 32'h0000_0001;
  assign array_update_76057[0] = add_74719 == 32'h0000_0000 ? array_update_76055 : array_update_76044[0];
  assign array_update_76057[1] = add_74719 == 32'h0000_0001 ? array_update_76055 : array_update_76044[1];
  assign array_update_76057[2] = add_74719 == 32'h0000_0002 ? array_update_76055 : array_update_76044[2];
  assign array_update_76057[3] = add_74719 == 32'h0000_0003 ? array_update_76055 : array_update_76044[3];
  assign array_update_76057[4] = add_74719 == 32'h0000_0004 ? array_update_76055 : array_update_76044[4];
  assign array_update_76057[5] = add_74719 == 32'h0000_0005 ? array_update_76055 : array_update_76044[5];
  assign array_update_76057[6] = add_74719 == 32'h0000_0006 ? array_update_76055 : array_update_76044[6];
  assign array_update_76057[7] = add_74719 == 32'h0000_0007 ? array_update_76055 : array_update_76044[7];
  assign array_update_76057[8] = add_74719 == 32'h0000_0008 ? array_update_76055 : array_update_76044[8];
  assign array_update_76057[9] = add_74719 == 32'h0000_0009 ? array_update_76055 : array_update_76044[9];
  assign array_index_76059 = array_update_72021[add_76056 > 32'h0000_0009 ? 4'h9 : add_76056[3:0]];
  assign array_index_76060 = array_update_76057[add_74719 > 32'h0000_0009 ? 4'h9 : add_74719[3:0]];
  assign smul_76064 = smul32b_32b_x_32b(array_index_74726[add_76056 > 32'h0000_0009 ? 4'h9 : add_76056[3:0]], array_index_76059[add_75937 > 32'h0000_0009 ? 4'h9 : add_75937[3:0]]);
  assign add_76066 = array_index_76060[add_75937 > 32'h0000_0009 ? 4'h9 : add_75937[3:0]] + smul_76064;
  assign array_update_76067[0] = add_75937 == 32'h0000_0000 ? add_76066 : array_index_76060[0];
  assign array_update_76067[1] = add_75937 == 32'h0000_0001 ? add_76066 : array_index_76060[1];
  assign array_update_76067[2] = add_75937 == 32'h0000_0002 ? add_76066 : array_index_76060[2];
  assign array_update_76067[3] = add_75937 == 32'h0000_0003 ? add_76066 : array_index_76060[3];
  assign array_update_76067[4] = add_75937 == 32'h0000_0004 ? add_76066 : array_index_76060[4];
  assign array_update_76067[5] = add_75937 == 32'h0000_0005 ? add_76066 : array_index_76060[5];
  assign array_update_76067[6] = add_75937 == 32'h0000_0006 ? add_76066 : array_index_76060[6];
  assign array_update_76067[7] = add_75937 == 32'h0000_0007 ? add_76066 : array_index_76060[7];
  assign array_update_76067[8] = add_75937 == 32'h0000_0008 ? add_76066 : array_index_76060[8];
  assign array_update_76067[9] = add_75937 == 32'h0000_0009 ? add_76066 : array_index_76060[9];
  assign array_update_76069[0] = add_74719 == 32'h0000_0000 ? array_update_76067 : array_update_76057[0];
  assign array_update_76069[1] = add_74719 == 32'h0000_0001 ? array_update_76067 : array_update_76057[1];
  assign array_update_76069[2] = add_74719 == 32'h0000_0002 ? array_update_76067 : array_update_76057[2];
  assign array_update_76069[3] = add_74719 == 32'h0000_0003 ? array_update_76067 : array_update_76057[3];
  assign array_update_76069[4] = add_74719 == 32'h0000_0004 ? array_update_76067 : array_update_76057[4];
  assign array_update_76069[5] = add_74719 == 32'h0000_0005 ? array_update_76067 : array_update_76057[5];
  assign array_update_76069[6] = add_74719 == 32'h0000_0006 ? array_update_76067 : array_update_76057[6];
  assign array_update_76069[7] = add_74719 == 32'h0000_0007 ? array_update_76067 : array_update_76057[7];
  assign array_update_76069[8] = add_74719 == 32'h0000_0008 ? array_update_76067 : array_update_76057[8];
  assign array_update_76069[9] = add_74719 == 32'h0000_0009 ? array_update_76067 : array_update_76057[9];
  assign add_76070 = add_74719 + 32'h0000_0001;
  assign array_index_76071 = array_update_76069[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign literal_76073 = 32'h0000_0000;
  assign array_update_76074[0] = literal_76073 == 32'h0000_0000 ? 32'h0000_0000 : array_index_76071[0];
  assign array_update_76074[1] = literal_76073 == 32'h0000_0001 ? 32'h0000_0000 : array_index_76071[1];
  assign array_update_76074[2] = literal_76073 == 32'h0000_0002 ? 32'h0000_0000 : array_index_76071[2];
  assign array_update_76074[3] = literal_76073 == 32'h0000_0003 ? 32'h0000_0000 : array_index_76071[3];
  assign array_update_76074[4] = literal_76073 == 32'h0000_0004 ? 32'h0000_0000 : array_index_76071[4];
  assign array_update_76074[5] = literal_76073 == 32'h0000_0005 ? 32'h0000_0000 : array_index_76071[5];
  assign array_update_76074[6] = literal_76073 == 32'h0000_0006 ? 32'h0000_0000 : array_index_76071[6];
  assign array_update_76074[7] = literal_76073 == 32'h0000_0007 ? 32'h0000_0000 : array_index_76071[7];
  assign array_update_76074[8] = literal_76073 == 32'h0000_0008 ? 32'h0000_0000 : array_index_76071[8];
  assign array_update_76074[9] = literal_76073 == 32'h0000_0009 ? 32'h0000_0000 : array_index_76071[9];
  assign literal_76075 = 32'h0000_0000;
  assign array_update_76076[0] = add_76070 == 32'h0000_0000 ? array_update_76074 : array_update_76069[0];
  assign array_update_76076[1] = add_76070 == 32'h0000_0001 ? array_update_76074 : array_update_76069[1];
  assign array_update_76076[2] = add_76070 == 32'h0000_0002 ? array_update_76074 : array_update_76069[2];
  assign array_update_76076[3] = add_76070 == 32'h0000_0003 ? array_update_76074 : array_update_76069[3];
  assign array_update_76076[4] = add_76070 == 32'h0000_0004 ? array_update_76074 : array_update_76069[4];
  assign array_update_76076[5] = add_76070 == 32'h0000_0005 ? array_update_76074 : array_update_76069[5];
  assign array_update_76076[6] = add_76070 == 32'h0000_0006 ? array_update_76074 : array_update_76069[6];
  assign array_update_76076[7] = add_76070 == 32'h0000_0007 ? array_update_76074 : array_update_76069[7];
  assign array_update_76076[8] = add_76070 == 32'h0000_0008 ? array_update_76074 : array_update_76069[8];
  assign array_update_76076[9] = add_76070 == 32'h0000_0009 ? array_update_76074 : array_update_76069[9];
  assign array_index_76077 = array_update_72020[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign array_index_76078 = array_update_72021[literal_76075 > 32'h0000_0009 ? 4'h9 : literal_76075[3:0]];
  assign array_index_76079 = array_update_76076[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_76083 = smul32b_32b_x_32b(array_index_76077[literal_76075 > 32'h0000_0009 ? 4'h9 : literal_76075[3:0]], array_index_76078[literal_76073 > 32'h0000_0009 ? 4'h9 : literal_76073[3:0]]);
  assign add_76085 = array_index_76079[literal_76073 > 32'h0000_0009 ? 4'h9 : literal_76073[3:0]] + smul_76083;
  assign array_update_76087[0] = literal_76073 == 32'h0000_0000 ? add_76085 : array_index_76079[0];
  assign array_update_76087[1] = literal_76073 == 32'h0000_0001 ? add_76085 : array_index_76079[1];
  assign array_update_76087[2] = literal_76073 == 32'h0000_0002 ? add_76085 : array_index_76079[2];
  assign array_update_76087[3] = literal_76073 == 32'h0000_0003 ? add_76085 : array_index_76079[3];
  assign array_update_76087[4] = literal_76073 == 32'h0000_0004 ? add_76085 : array_index_76079[4];
  assign array_update_76087[5] = literal_76073 == 32'h0000_0005 ? add_76085 : array_index_76079[5];
  assign array_update_76087[6] = literal_76073 == 32'h0000_0006 ? add_76085 : array_index_76079[6];
  assign array_update_76087[7] = literal_76073 == 32'h0000_0007 ? add_76085 : array_index_76079[7];
  assign array_update_76087[8] = literal_76073 == 32'h0000_0008 ? add_76085 : array_index_76079[8];
  assign array_update_76087[9] = literal_76073 == 32'h0000_0009 ? add_76085 : array_index_76079[9];
  assign add_76088 = literal_76075 + 32'h0000_0001;
  assign array_update_76089[0] = add_76070 == 32'h0000_0000 ? array_update_76087 : array_update_76076[0];
  assign array_update_76089[1] = add_76070 == 32'h0000_0001 ? array_update_76087 : array_update_76076[1];
  assign array_update_76089[2] = add_76070 == 32'h0000_0002 ? array_update_76087 : array_update_76076[2];
  assign array_update_76089[3] = add_76070 == 32'h0000_0003 ? array_update_76087 : array_update_76076[3];
  assign array_update_76089[4] = add_76070 == 32'h0000_0004 ? array_update_76087 : array_update_76076[4];
  assign array_update_76089[5] = add_76070 == 32'h0000_0005 ? array_update_76087 : array_update_76076[5];
  assign array_update_76089[6] = add_76070 == 32'h0000_0006 ? array_update_76087 : array_update_76076[6];
  assign array_update_76089[7] = add_76070 == 32'h0000_0007 ? array_update_76087 : array_update_76076[7];
  assign array_update_76089[8] = add_76070 == 32'h0000_0008 ? array_update_76087 : array_update_76076[8];
  assign array_update_76089[9] = add_76070 == 32'h0000_0009 ? array_update_76087 : array_update_76076[9];
  assign array_index_76091 = array_update_72021[add_76088 > 32'h0000_0009 ? 4'h9 : add_76088[3:0]];
  assign array_index_76092 = array_update_76089[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_76096 = smul32b_32b_x_32b(array_index_76077[add_76088 > 32'h0000_0009 ? 4'h9 : add_76088[3:0]], array_index_76091[literal_76073 > 32'h0000_0009 ? 4'h9 : literal_76073[3:0]]);
  assign add_76098 = array_index_76092[literal_76073 > 32'h0000_0009 ? 4'h9 : literal_76073[3:0]] + smul_76096;
  assign array_update_76100[0] = literal_76073 == 32'h0000_0000 ? add_76098 : array_index_76092[0];
  assign array_update_76100[1] = literal_76073 == 32'h0000_0001 ? add_76098 : array_index_76092[1];
  assign array_update_76100[2] = literal_76073 == 32'h0000_0002 ? add_76098 : array_index_76092[2];
  assign array_update_76100[3] = literal_76073 == 32'h0000_0003 ? add_76098 : array_index_76092[3];
  assign array_update_76100[4] = literal_76073 == 32'h0000_0004 ? add_76098 : array_index_76092[4];
  assign array_update_76100[5] = literal_76073 == 32'h0000_0005 ? add_76098 : array_index_76092[5];
  assign array_update_76100[6] = literal_76073 == 32'h0000_0006 ? add_76098 : array_index_76092[6];
  assign array_update_76100[7] = literal_76073 == 32'h0000_0007 ? add_76098 : array_index_76092[7];
  assign array_update_76100[8] = literal_76073 == 32'h0000_0008 ? add_76098 : array_index_76092[8];
  assign array_update_76100[9] = literal_76073 == 32'h0000_0009 ? add_76098 : array_index_76092[9];
  assign add_76101 = add_76088 + 32'h0000_0001;
  assign array_update_76102[0] = add_76070 == 32'h0000_0000 ? array_update_76100 : array_update_76089[0];
  assign array_update_76102[1] = add_76070 == 32'h0000_0001 ? array_update_76100 : array_update_76089[1];
  assign array_update_76102[2] = add_76070 == 32'h0000_0002 ? array_update_76100 : array_update_76089[2];
  assign array_update_76102[3] = add_76070 == 32'h0000_0003 ? array_update_76100 : array_update_76089[3];
  assign array_update_76102[4] = add_76070 == 32'h0000_0004 ? array_update_76100 : array_update_76089[4];
  assign array_update_76102[5] = add_76070 == 32'h0000_0005 ? array_update_76100 : array_update_76089[5];
  assign array_update_76102[6] = add_76070 == 32'h0000_0006 ? array_update_76100 : array_update_76089[6];
  assign array_update_76102[7] = add_76070 == 32'h0000_0007 ? array_update_76100 : array_update_76089[7];
  assign array_update_76102[8] = add_76070 == 32'h0000_0008 ? array_update_76100 : array_update_76089[8];
  assign array_update_76102[9] = add_76070 == 32'h0000_0009 ? array_update_76100 : array_update_76089[9];
  assign array_index_76104 = array_update_72021[add_76101 > 32'h0000_0009 ? 4'h9 : add_76101[3:0]];
  assign array_index_76105 = array_update_76102[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_76109 = smul32b_32b_x_32b(array_index_76077[add_76101 > 32'h0000_0009 ? 4'h9 : add_76101[3:0]], array_index_76104[literal_76073 > 32'h0000_0009 ? 4'h9 : literal_76073[3:0]]);
  assign add_76111 = array_index_76105[literal_76073 > 32'h0000_0009 ? 4'h9 : literal_76073[3:0]] + smul_76109;
  assign array_update_76113[0] = literal_76073 == 32'h0000_0000 ? add_76111 : array_index_76105[0];
  assign array_update_76113[1] = literal_76073 == 32'h0000_0001 ? add_76111 : array_index_76105[1];
  assign array_update_76113[2] = literal_76073 == 32'h0000_0002 ? add_76111 : array_index_76105[2];
  assign array_update_76113[3] = literal_76073 == 32'h0000_0003 ? add_76111 : array_index_76105[3];
  assign array_update_76113[4] = literal_76073 == 32'h0000_0004 ? add_76111 : array_index_76105[4];
  assign array_update_76113[5] = literal_76073 == 32'h0000_0005 ? add_76111 : array_index_76105[5];
  assign array_update_76113[6] = literal_76073 == 32'h0000_0006 ? add_76111 : array_index_76105[6];
  assign array_update_76113[7] = literal_76073 == 32'h0000_0007 ? add_76111 : array_index_76105[7];
  assign array_update_76113[8] = literal_76073 == 32'h0000_0008 ? add_76111 : array_index_76105[8];
  assign array_update_76113[9] = literal_76073 == 32'h0000_0009 ? add_76111 : array_index_76105[9];
  assign add_76114 = add_76101 + 32'h0000_0001;
  assign array_update_76115[0] = add_76070 == 32'h0000_0000 ? array_update_76113 : array_update_76102[0];
  assign array_update_76115[1] = add_76070 == 32'h0000_0001 ? array_update_76113 : array_update_76102[1];
  assign array_update_76115[2] = add_76070 == 32'h0000_0002 ? array_update_76113 : array_update_76102[2];
  assign array_update_76115[3] = add_76070 == 32'h0000_0003 ? array_update_76113 : array_update_76102[3];
  assign array_update_76115[4] = add_76070 == 32'h0000_0004 ? array_update_76113 : array_update_76102[4];
  assign array_update_76115[5] = add_76070 == 32'h0000_0005 ? array_update_76113 : array_update_76102[5];
  assign array_update_76115[6] = add_76070 == 32'h0000_0006 ? array_update_76113 : array_update_76102[6];
  assign array_update_76115[7] = add_76070 == 32'h0000_0007 ? array_update_76113 : array_update_76102[7];
  assign array_update_76115[8] = add_76070 == 32'h0000_0008 ? array_update_76113 : array_update_76102[8];
  assign array_update_76115[9] = add_76070 == 32'h0000_0009 ? array_update_76113 : array_update_76102[9];
  assign array_index_76117 = array_update_72021[add_76114 > 32'h0000_0009 ? 4'h9 : add_76114[3:0]];
  assign array_index_76118 = array_update_76115[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_76122 = smul32b_32b_x_32b(array_index_76077[add_76114 > 32'h0000_0009 ? 4'h9 : add_76114[3:0]], array_index_76117[literal_76073 > 32'h0000_0009 ? 4'h9 : literal_76073[3:0]]);
  assign add_76124 = array_index_76118[literal_76073 > 32'h0000_0009 ? 4'h9 : literal_76073[3:0]] + smul_76122;
  assign array_update_76126[0] = literal_76073 == 32'h0000_0000 ? add_76124 : array_index_76118[0];
  assign array_update_76126[1] = literal_76073 == 32'h0000_0001 ? add_76124 : array_index_76118[1];
  assign array_update_76126[2] = literal_76073 == 32'h0000_0002 ? add_76124 : array_index_76118[2];
  assign array_update_76126[3] = literal_76073 == 32'h0000_0003 ? add_76124 : array_index_76118[3];
  assign array_update_76126[4] = literal_76073 == 32'h0000_0004 ? add_76124 : array_index_76118[4];
  assign array_update_76126[5] = literal_76073 == 32'h0000_0005 ? add_76124 : array_index_76118[5];
  assign array_update_76126[6] = literal_76073 == 32'h0000_0006 ? add_76124 : array_index_76118[6];
  assign array_update_76126[7] = literal_76073 == 32'h0000_0007 ? add_76124 : array_index_76118[7];
  assign array_update_76126[8] = literal_76073 == 32'h0000_0008 ? add_76124 : array_index_76118[8];
  assign array_update_76126[9] = literal_76073 == 32'h0000_0009 ? add_76124 : array_index_76118[9];
  assign add_76127 = add_76114 + 32'h0000_0001;
  assign array_update_76128[0] = add_76070 == 32'h0000_0000 ? array_update_76126 : array_update_76115[0];
  assign array_update_76128[1] = add_76070 == 32'h0000_0001 ? array_update_76126 : array_update_76115[1];
  assign array_update_76128[2] = add_76070 == 32'h0000_0002 ? array_update_76126 : array_update_76115[2];
  assign array_update_76128[3] = add_76070 == 32'h0000_0003 ? array_update_76126 : array_update_76115[3];
  assign array_update_76128[4] = add_76070 == 32'h0000_0004 ? array_update_76126 : array_update_76115[4];
  assign array_update_76128[5] = add_76070 == 32'h0000_0005 ? array_update_76126 : array_update_76115[5];
  assign array_update_76128[6] = add_76070 == 32'h0000_0006 ? array_update_76126 : array_update_76115[6];
  assign array_update_76128[7] = add_76070 == 32'h0000_0007 ? array_update_76126 : array_update_76115[7];
  assign array_update_76128[8] = add_76070 == 32'h0000_0008 ? array_update_76126 : array_update_76115[8];
  assign array_update_76128[9] = add_76070 == 32'h0000_0009 ? array_update_76126 : array_update_76115[9];
  assign array_index_76130 = array_update_72021[add_76127 > 32'h0000_0009 ? 4'h9 : add_76127[3:0]];
  assign array_index_76131 = array_update_76128[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_76135 = smul32b_32b_x_32b(array_index_76077[add_76127 > 32'h0000_0009 ? 4'h9 : add_76127[3:0]], array_index_76130[literal_76073 > 32'h0000_0009 ? 4'h9 : literal_76073[3:0]]);
  assign add_76137 = array_index_76131[literal_76073 > 32'h0000_0009 ? 4'h9 : literal_76073[3:0]] + smul_76135;
  assign array_update_76139[0] = literal_76073 == 32'h0000_0000 ? add_76137 : array_index_76131[0];
  assign array_update_76139[1] = literal_76073 == 32'h0000_0001 ? add_76137 : array_index_76131[1];
  assign array_update_76139[2] = literal_76073 == 32'h0000_0002 ? add_76137 : array_index_76131[2];
  assign array_update_76139[3] = literal_76073 == 32'h0000_0003 ? add_76137 : array_index_76131[3];
  assign array_update_76139[4] = literal_76073 == 32'h0000_0004 ? add_76137 : array_index_76131[4];
  assign array_update_76139[5] = literal_76073 == 32'h0000_0005 ? add_76137 : array_index_76131[5];
  assign array_update_76139[6] = literal_76073 == 32'h0000_0006 ? add_76137 : array_index_76131[6];
  assign array_update_76139[7] = literal_76073 == 32'h0000_0007 ? add_76137 : array_index_76131[7];
  assign array_update_76139[8] = literal_76073 == 32'h0000_0008 ? add_76137 : array_index_76131[8];
  assign array_update_76139[9] = literal_76073 == 32'h0000_0009 ? add_76137 : array_index_76131[9];
  assign add_76140 = add_76127 + 32'h0000_0001;
  assign array_update_76141[0] = add_76070 == 32'h0000_0000 ? array_update_76139 : array_update_76128[0];
  assign array_update_76141[1] = add_76070 == 32'h0000_0001 ? array_update_76139 : array_update_76128[1];
  assign array_update_76141[2] = add_76070 == 32'h0000_0002 ? array_update_76139 : array_update_76128[2];
  assign array_update_76141[3] = add_76070 == 32'h0000_0003 ? array_update_76139 : array_update_76128[3];
  assign array_update_76141[4] = add_76070 == 32'h0000_0004 ? array_update_76139 : array_update_76128[4];
  assign array_update_76141[5] = add_76070 == 32'h0000_0005 ? array_update_76139 : array_update_76128[5];
  assign array_update_76141[6] = add_76070 == 32'h0000_0006 ? array_update_76139 : array_update_76128[6];
  assign array_update_76141[7] = add_76070 == 32'h0000_0007 ? array_update_76139 : array_update_76128[7];
  assign array_update_76141[8] = add_76070 == 32'h0000_0008 ? array_update_76139 : array_update_76128[8];
  assign array_update_76141[9] = add_76070 == 32'h0000_0009 ? array_update_76139 : array_update_76128[9];
  assign array_index_76143 = array_update_72021[add_76140 > 32'h0000_0009 ? 4'h9 : add_76140[3:0]];
  assign array_index_76144 = array_update_76141[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_76148 = smul32b_32b_x_32b(array_index_76077[add_76140 > 32'h0000_0009 ? 4'h9 : add_76140[3:0]], array_index_76143[literal_76073 > 32'h0000_0009 ? 4'h9 : literal_76073[3:0]]);
  assign add_76150 = array_index_76144[literal_76073 > 32'h0000_0009 ? 4'h9 : literal_76073[3:0]] + smul_76148;
  assign array_update_76152[0] = literal_76073 == 32'h0000_0000 ? add_76150 : array_index_76144[0];
  assign array_update_76152[1] = literal_76073 == 32'h0000_0001 ? add_76150 : array_index_76144[1];
  assign array_update_76152[2] = literal_76073 == 32'h0000_0002 ? add_76150 : array_index_76144[2];
  assign array_update_76152[3] = literal_76073 == 32'h0000_0003 ? add_76150 : array_index_76144[3];
  assign array_update_76152[4] = literal_76073 == 32'h0000_0004 ? add_76150 : array_index_76144[4];
  assign array_update_76152[5] = literal_76073 == 32'h0000_0005 ? add_76150 : array_index_76144[5];
  assign array_update_76152[6] = literal_76073 == 32'h0000_0006 ? add_76150 : array_index_76144[6];
  assign array_update_76152[7] = literal_76073 == 32'h0000_0007 ? add_76150 : array_index_76144[7];
  assign array_update_76152[8] = literal_76073 == 32'h0000_0008 ? add_76150 : array_index_76144[8];
  assign array_update_76152[9] = literal_76073 == 32'h0000_0009 ? add_76150 : array_index_76144[9];
  assign add_76153 = add_76140 + 32'h0000_0001;
  assign array_update_76154[0] = add_76070 == 32'h0000_0000 ? array_update_76152 : array_update_76141[0];
  assign array_update_76154[1] = add_76070 == 32'h0000_0001 ? array_update_76152 : array_update_76141[1];
  assign array_update_76154[2] = add_76070 == 32'h0000_0002 ? array_update_76152 : array_update_76141[2];
  assign array_update_76154[3] = add_76070 == 32'h0000_0003 ? array_update_76152 : array_update_76141[3];
  assign array_update_76154[4] = add_76070 == 32'h0000_0004 ? array_update_76152 : array_update_76141[4];
  assign array_update_76154[5] = add_76070 == 32'h0000_0005 ? array_update_76152 : array_update_76141[5];
  assign array_update_76154[6] = add_76070 == 32'h0000_0006 ? array_update_76152 : array_update_76141[6];
  assign array_update_76154[7] = add_76070 == 32'h0000_0007 ? array_update_76152 : array_update_76141[7];
  assign array_update_76154[8] = add_76070 == 32'h0000_0008 ? array_update_76152 : array_update_76141[8];
  assign array_update_76154[9] = add_76070 == 32'h0000_0009 ? array_update_76152 : array_update_76141[9];
  assign array_index_76156 = array_update_72021[add_76153 > 32'h0000_0009 ? 4'h9 : add_76153[3:0]];
  assign array_index_76157 = array_update_76154[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_76161 = smul32b_32b_x_32b(array_index_76077[add_76153 > 32'h0000_0009 ? 4'h9 : add_76153[3:0]], array_index_76156[literal_76073 > 32'h0000_0009 ? 4'h9 : literal_76073[3:0]]);
  assign add_76163 = array_index_76157[literal_76073 > 32'h0000_0009 ? 4'h9 : literal_76073[3:0]] + smul_76161;
  assign array_update_76165[0] = literal_76073 == 32'h0000_0000 ? add_76163 : array_index_76157[0];
  assign array_update_76165[1] = literal_76073 == 32'h0000_0001 ? add_76163 : array_index_76157[1];
  assign array_update_76165[2] = literal_76073 == 32'h0000_0002 ? add_76163 : array_index_76157[2];
  assign array_update_76165[3] = literal_76073 == 32'h0000_0003 ? add_76163 : array_index_76157[3];
  assign array_update_76165[4] = literal_76073 == 32'h0000_0004 ? add_76163 : array_index_76157[4];
  assign array_update_76165[5] = literal_76073 == 32'h0000_0005 ? add_76163 : array_index_76157[5];
  assign array_update_76165[6] = literal_76073 == 32'h0000_0006 ? add_76163 : array_index_76157[6];
  assign array_update_76165[7] = literal_76073 == 32'h0000_0007 ? add_76163 : array_index_76157[7];
  assign array_update_76165[8] = literal_76073 == 32'h0000_0008 ? add_76163 : array_index_76157[8];
  assign array_update_76165[9] = literal_76073 == 32'h0000_0009 ? add_76163 : array_index_76157[9];
  assign add_76166 = add_76153 + 32'h0000_0001;
  assign array_update_76167[0] = add_76070 == 32'h0000_0000 ? array_update_76165 : array_update_76154[0];
  assign array_update_76167[1] = add_76070 == 32'h0000_0001 ? array_update_76165 : array_update_76154[1];
  assign array_update_76167[2] = add_76070 == 32'h0000_0002 ? array_update_76165 : array_update_76154[2];
  assign array_update_76167[3] = add_76070 == 32'h0000_0003 ? array_update_76165 : array_update_76154[3];
  assign array_update_76167[4] = add_76070 == 32'h0000_0004 ? array_update_76165 : array_update_76154[4];
  assign array_update_76167[5] = add_76070 == 32'h0000_0005 ? array_update_76165 : array_update_76154[5];
  assign array_update_76167[6] = add_76070 == 32'h0000_0006 ? array_update_76165 : array_update_76154[6];
  assign array_update_76167[7] = add_76070 == 32'h0000_0007 ? array_update_76165 : array_update_76154[7];
  assign array_update_76167[8] = add_76070 == 32'h0000_0008 ? array_update_76165 : array_update_76154[8];
  assign array_update_76167[9] = add_76070 == 32'h0000_0009 ? array_update_76165 : array_update_76154[9];
  assign array_index_76169 = array_update_72021[add_76166 > 32'h0000_0009 ? 4'h9 : add_76166[3:0]];
  assign array_index_76170 = array_update_76167[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_76174 = smul32b_32b_x_32b(array_index_76077[add_76166 > 32'h0000_0009 ? 4'h9 : add_76166[3:0]], array_index_76169[literal_76073 > 32'h0000_0009 ? 4'h9 : literal_76073[3:0]]);
  assign add_76176 = array_index_76170[literal_76073 > 32'h0000_0009 ? 4'h9 : literal_76073[3:0]] + smul_76174;
  assign array_update_76178[0] = literal_76073 == 32'h0000_0000 ? add_76176 : array_index_76170[0];
  assign array_update_76178[1] = literal_76073 == 32'h0000_0001 ? add_76176 : array_index_76170[1];
  assign array_update_76178[2] = literal_76073 == 32'h0000_0002 ? add_76176 : array_index_76170[2];
  assign array_update_76178[3] = literal_76073 == 32'h0000_0003 ? add_76176 : array_index_76170[3];
  assign array_update_76178[4] = literal_76073 == 32'h0000_0004 ? add_76176 : array_index_76170[4];
  assign array_update_76178[5] = literal_76073 == 32'h0000_0005 ? add_76176 : array_index_76170[5];
  assign array_update_76178[6] = literal_76073 == 32'h0000_0006 ? add_76176 : array_index_76170[6];
  assign array_update_76178[7] = literal_76073 == 32'h0000_0007 ? add_76176 : array_index_76170[7];
  assign array_update_76178[8] = literal_76073 == 32'h0000_0008 ? add_76176 : array_index_76170[8];
  assign array_update_76178[9] = literal_76073 == 32'h0000_0009 ? add_76176 : array_index_76170[9];
  assign add_76179 = add_76166 + 32'h0000_0001;
  assign array_update_76180[0] = add_76070 == 32'h0000_0000 ? array_update_76178 : array_update_76167[0];
  assign array_update_76180[1] = add_76070 == 32'h0000_0001 ? array_update_76178 : array_update_76167[1];
  assign array_update_76180[2] = add_76070 == 32'h0000_0002 ? array_update_76178 : array_update_76167[2];
  assign array_update_76180[3] = add_76070 == 32'h0000_0003 ? array_update_76178 : array_update_76167[3];
  assign array_update_76180[4] = add_76070 == 32'h0000_0004 ? array_update_76178 : array_update_76167[4];
  assign array_update_76180[5] = add_76070 == 32'h0000_0005 ? array_update_76178 : array_update_76167[5];
  assign array_update_76180[6] = add_76070 == 32'h0000_0006 ? array_update_76178 : array_update_76167[6];
  assign array_update_76180[7] = add_76070 == 32'h0000_0007 ? array_update_76178 : array_update_76167[7];
  assign array_update_76180[8] = add_76070 == 32'h0000_0008 ? array_update_76178 : array_update_76167[8];
  assign array_update_76180[9] = add_76070 == 32'h0000_0009 ? array_update_76178 : array_update_76167[9];
  assign array_index_76182 = array_update_72021[add_76179 > 32'h0000_0009 ? 4'h9 : add_76179[3:0]];
  assign array_index_76183 = array_update_76180[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_76187 = smul32b_32b_x_32b(array_index_76077[add_76179 > 32'h0000_0009 ? 4'h9 : add_76179[3:0]], array_index_76182[literal_76073 > 32'h0000_0009 ? 4'h9 : literal_76073[3:0]]);
  assign add_76189 = array_index_76183[literal_76073 > 32'h0000_0009 ? 4'h9 : literal_76073[3:0]] + smul_76187;
  assign array_update_76191[0] = literal_76073 == 32'h0000_0000 ? add_76189 : array_index_76183[0];
  assign array_update_76191[1] = literal_76073 == 32'h0000_0001 ? add_76189 : array_index_76183[1];
  assign array_update_76191[2] = literal_76073 == 32'h0000_0002 ? add_76189 : array_index_76183[2];
  assign array_update_76191[3] = literal_76073 == 32'h0000_0003 ? add_76189 : array_index_76183[3];
  assign array_update_76191[4] = literal_76073 == 32'h0000_0004 ? add_76189 : array_index_76183[4];
  assign array_update_76191[5] = literal_76073 == 32'h0000_0005 ? add_76189 : array_index_76183[5];
  assign array_update_76191[6] = literal_76073 == 32'h0000_0006 ? add_76189 : array_index_76183[6];
  assign array_update_76191[7] = literal_76073 == 32'h0000_0007 ? add_76189 : array_index_76183[7];
  assign array_update_76191[8] = literal_76073 == 32'h0000_0008 ? add_76189 : array_index_76183[8];
  assign array_update_76191[9] = literal_76073 == 32'h0000_0009 ? add_76189 : array_index_76183[9];
  assign add_76192 = add_76179 + 32'h0000_0001;
  assign array_update_76193[0] = add_76070 == 32'h0000_0000 ? array_update_76191 : array_update_76180[0];
  assign array_update_76193[1] = add_76070 == 32'h0000_0001 ? array_update_76191 : array_update_76180[1];
  assign array_update_76193[2] = add_76070 == 32'h0000_0002 ? array_update_76191 : array_update_76180[2];
  assign array_update_76193[3] = add_76070 == 32'h0000_0003 ? array_update_76191 : array_update_76180[3];
  assign array_update_76193[4] = add_76070 == 32'h0000_0004 ? array_update_76191 : array_update_76180[4];
  assign array_update_76193[5] = add_76070 == 32'h0000_0005 ? array_update_76191 : array_update_76180[5];
  assign array_update_76193[6] = add_76070 == 32'h0000_0006 ? array_update_76191 : array_update_76180[6];
  assign array_update_76193[7] = add_76070 == 32'h0000_0007 ? array_update_76191 : array_update_76180[7];
  assign array_update_76193[8] = add_76070 == 32'h0000_0008 ? array_update_76191 : array_update_76180[8];
  assign array_update_76193[9] = add_76070 == 32'h0000_0009 ? array_update_76191 : array_update_76180[9];
  assign array_index_76195 = array_update_72021[add_76192 > 32'h0000_0009 ? 4'h9 : add_76192[3:0]];
  assign array_index_76196 = array_update_76193[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_76200 = smul32b_32b_x_32b(array_index_76077[add_76192 > 32'h0000_0009 ? 4'h9 : add_76192[3:0]], array_index_76195[literal_76073 > 32'h0000_0009 ? 4'h9 : literal_76073[3:0]]);
  assign add_76202 = array_index_76196[literal_76073 > 32'h0000_0009 ? 4'h9 : literal_76073[3:0]] + smul_76200;
  assign array_update_76203[0] = literal_76073 == 32'h0000_0000 ? add_76202 : array_index_76196[0];
  assign array_update_76203[1] = literal_76073 == 32'h0000_0001 ? add_76202 : array_index_76196[1];
  assign array_update_76203[2] = literal_76073 == 32'h0000_0002 ? add_76202 : array_index_76196[2];
  assign array_update_76203[3] = literal_76073 == 32'h0000_0003 ? add_76202 : array_index_76196[3];
  assign array_update_76203[4] = literal_76073 == 32'h0000_0004 ? add_76202 : array_index_76196[4];
  assign array_update_76203[5] = literal_76073 == 32'h0000_0005 ? add_76202 : array_index_76196[5];
  assign array_update_76203[6] = literal_76073 == 32'h0000_0006 ? add_76202 : array_index_76196[6];
  assign array_update_76203[7] = literal_76073 == 32'h0000_0007 ? add_76202 : array_index_76196[7];
  assign array_update_76203[8] = literal_76073 == 32'h0000_0008 ? add_76202 : array_index_76196[8];
  assign array_update_76203[9] = literal_76073 == 32'h0000_0009 ? add_76202 : array_index_76196[9];
  assign array_update_76204[0] = add_76070 == 32'h0000_0000 ? array_update_76203 : array_update_76193[0];
  assign array_update_76204[1] = add_76070 == 32'h0000_0001 ? array_update_76203 : array_update_76193[1];
  assign array_update_76204[2] = add_76070 == 32'h0000_0002 ? array_update_76203 : array_update_76193[2];
  assign array_update_76204[3] = add_76070 == 32'h0000_0003 ? array_update_76203 : array_update_76193[3];
  assign array_update_76204[4] = add_76070 == 32'h0000_0004 ? array_update_76203 : array_update_76193[4];
  assign array_update_76204[5] = add_76070 == 32'h0000_0005 ? array_update_76203 : array_update_76193[5];
  assign array_update_76204[6] = add_76070 == 32'h0000_0006 ? array_update_76203 : array_update_76193[6];
  assign array_update_76204[7] = add_76070 == 32'h0000_0007 ? array_update_76203 : array_update_76193[7];
  assign array_update_76204[8] = add_76070 == 32'h0000_0008 ? array_update_76203 : array_update_76193[8];
  assign array_update_76204[9] = add_76070 == 32'h0000_0009 ? array_update_76203 : array_update_76193[9];
  assign array_index_76206 = array_update_76204[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign add_76208 = literal_76073 + 32'h0000_0001;
  assign array_update_76209[0] = add_76208 == 32'h0000_0000 ? 32'h0000_0000 : array_index_76206[0];
  assign array_update_76209[1] = add_76208 == 32'h0000_0001 ? 32'h0000_0000 : array_index_76206[1];
  assign array_update_76209[2] = add_76208 == 32'h0000_0002 ? 32'h0000_0000 : array_index_76206[2];
  assign array_update_76209[3] = add_76208 == 32'h0000_0003 ? 32'h0000_0000 : array_index_76206[3];
  assign array_update_76209[4] = add_76208 == 32'h0000_0004 ? 32'h0000_0000 : array_index_76206[4];
  assign array_update_76209[5] = add_76208 == 32'h0000_0005 ? 32'h0000_0000 : array_index_76206[5];
  assign array_update_76209[6] = add_76208 == 32'h0000_0006 ? 32'h0000_0000 : array_index_76206[6];
  assign array_update_76209[7] = add_76208 == 32'h0000_0007 ? 32'h0000_0000 : array_index_76206[7];
  assign array_update_76209[8] = add_76208 == 32'h0000_0008 ? 32'h0000_0000 : array_index_76206[8];
  assign array_update_76209[9] = add_76208 == 32'h0000_0009 ? 32'h0000_0000 : array_index_76206[9];
  assign literal_76210 = 32'h0000_0000;
  assign array_update_76211[0] = add_76070 == 32'h0000_0000 ? array_update_76209 : array_update_76204[0];
  assign array_update_76211[1] = add_76070 == 32'h0000_0001 ? array_update_76209 : array_update_76204[1];
  assign array_update_76211[2] = add_76070 == 32'h0000_0002 ? array_update_76209 : array_update_76204[2];
  assign array_update_76211[3] = add_76070 == 32'h0000_0003 ? array_update_76209 : array_update_76204[3];
  assign array_update_76211[4] = add_76070 == 32'h0000_0004 ? array_update_76209 : array_update_76204[4];
  assign array_update_76211[5] = add_76070 == 32'h0000_0005 ? array_update_76209 : array_update_76204[5];
  assign array_update_76211[6] = add_76070 == 32'h0000_0006 ? array_update_76209 : array_update_76204[6];
  assign array_update_76211[7] = add_76070 == 32'h0000_0007 ? array_update_76209 : array_update_76204[7];
  assign array_update_76211[8] = add_76070 == 32'h0000_0008 ? array_update_76209 : array_update_76204[8];
  assign array_update_76211[9] = add_76070 == 32'h0000_0009 ? array_update_76209 : array_update_76204[9];
  assign array_index_76213 = array_update_72021[literal_76210 > 32'h0000_0009 ? 4'h9 : literal_76210[3:0]];
  assign array_index_76214 = array_update_76211[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_76218 = smul32b_32b_x_32b(array_index_76077[literal_76210 > 32'h0000_0009 ? 4'h9 : literal_76210[3:0]], array_index_76213[add_76208 > 32'h0000_0009 ? 4'h9 : add_76208[3:0]]);
  assign add_76220 = array_index_76214[add_76208 > 32'h0000_0009 ? 4'h9 : add_76208[3:0]] + smul_76218;
  assign array_update_76222[0] = add_76208 == 32'h0000_0000 ? add_76220 : array_index_76214[0];
  assign array_update_76222[1] = add_76208 == 32'h0000_0001 ? add_76220 : array_index_76214[1];
  assign array_update_76222[2] = add_76208 == 32'h0000_0002 ? add_76220 : array_index_76214[2];
  assign array_update_76222[3] = add_76208 == 32'h0000_0003 ? add_76220 : array_index_76214[3];
  assign array_update_76222[4] = add_76208 == 32'h0000_0004 ? add_76220 : array_index_76214[4];
  assign array_update_76222[5] = add_76208 == 32'h0000_0005 ? add_76220 : array_index_76214[5];
  assign array_update_76222[6] = add_76208 == 32'h0000_0006 ? add_76220 : array_index_76214[6];
  assign array_update_76222[7] = add_76208 == 32'h0000_0007 ? add_76220 : array_index_76214[7];
  assign array_update_76222[8] = add_76208 == 32'h0000_0008 ? add_76220 : array_index_76214[8];
  assign array_update_76222[9] = add_76208 == 32'h0000_0009 ? add_76220 : array_index_76214[9];
  assign add_76223 = literal_76210 + 32'h0000_0001;
  assign array_update_76224[0] = add_76070 == 32'h0000_0000 ? array_update_76222 : array_update_76211[0];
  assign array_update_76224[1] = add_76070 == 32'h0000_0001 ? array_update_76222 : array_update_76211[1];
  assign array_update_76224[2] = add_76070 == 32'h0000_0002 ? array_update_76222 : array_update_76211[2];
  assign array_update_76224[3] = add_76070 == 32'h0000_0003 ? array_update_76222 : array_update_76211[3];
  assign array_update_76224[4] = add_76070 == 32'h0000_0004 ? array_update_76222 : array_update_76211[4];
  assign array_update_76224[5] = add_76070 == 32'h0000_0005 ? array_update_76222 : array_update_76211[5];
  assign array_update_76224[6] = add_76070 == 32'h0000_0006 ? array_update_76222 : array_update_76211[6];
  assign array_update_76224[7] = add_76070 == 32'h0000_0007 ? array_update_76222 : array_update_76211[7];
  assign array_update_76224[8] = add_76070 == 32'h0000_0008 ? array_update_76222 : array_update_76211[8];
  assign array_update_76224[9] = add_76070 == 32'h0000_0009 ? array_update_76222 : array_update_76211[9];
  assign array_index_76226 = array_update_72021[add_76223 > 32'h0000_0009 ? 4'h9 : add_76223[3:0]];
  assign array_index_76227 = array_update_76224[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_76231 = smul32b_32b_x_32b(array_index_76077[add_76223 > 32'h0000_0009 ? 4'h9 : add_76223[3:0]], array_index_76226[add_76208 > 32'h0000_0009 ? 4'h9 : add_76208[3:0]]);
  assign add_76233 = array_index_76227[add_76208 > 32'h0000_0009 ? 4'h9 : add_76208[3:0]] + smul_76231;
  assign array_update_76235[0] = add_76208 == 32'h0000_0000 ? add_76233 : array_index_76227[0];
  assign array_update_76235[1] = add_76208 == 32'h0000_0001 ? add_76233 : array_index_76227[1];
  assign array_update_76235[2] = add_76208 == 32'h0000_0002 ? add_76233 : array_index_76227[2];
  assign array_update_76235[3] = add_76208 == 32'h0000_0003 ? add_76233 : array_index_76227[3];
  assign array_update_76235[4] = add_76208 == 32'h0000_0004 ? add_76233 : array_index_76227[4];
  assign array_update_76235[5] = add_76208 == 32'h0000_0005 ? add_76233 : array_index_76227[5];
  assign array_update_76235[6] = add_76208 == 32'h0000_0006 ? add_76233 : array_index_76227[6];
  assign array_update_76235[7] = add_76208 == 32'h0000_0007 ? add_76233 : array_index_76227[7];
  assign array_update_76235[8] = add_76208 == 32'h0000_0008 ? add_76233 : array_index_76227[8];
  assign array_update_76235[9] = add_76208 == 32'h0000_0009 ? add_76233 : array_index_76227[9];
  assign add_76236 = add_76223 + 32'h0000_0001;
  assign array_update_76237[0] = add_76070 == 32'h0000_0000 ? array_update_76235 : array_update_76224[0];
  assign array_update_76237[1] = add_76070 == 32'h0000_0001 ? array_update_76235 : array_update_76224[1];
  assign array_update_76237[2] = add_76070 == 32'h0000_0002 ? array_update_76235 : array_update_76224[2];
  assign array_update_76237[3] = add_76070 == 32'h0000_0003 ? array_update_76235 : array_update_76224[3];
  assign array_update_76237[4] = add_76070 == 32'h0000_0004 ? array_update_76235 : array_update_76224[4];
  assign array_update_76237[5] = add_76070 == 32'h0000_0005 ? array_update_76235 : array_update_76224[5];
  assign array_update_76237[6] = add_76070 == 32'h0000_0006 ? array_update_76235 : array_update_76224[6];
  assign array_update_76237[7] = add_76070 == 32'h0000_0007 ? array_update_76235 : array_update_76224[7];
  assign array_update_76237[8] = add_76070 == 32'h0000_0008 ? array_update_76235 : array_update_76224[8];
  assign array_update_76237[9] = add_76070 == 32'h0000_0009 ? array_update_76235 : array_update_76224[9];
  assign array_index_76239 = array_update_72021[add_76236 > 32'h0000_0009 ? 4'h9 : add_76236[3:0]];
  assign array_index_76240 = array_update_76237[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_76244 = smul32b_32b_x_32b(array_index_76077[add_76236 > 32'h0000_0009 ? 4'h9 : add_76236[3:0]], array_index_76239[add_76208 > 32'h0000_0009 ? 4'h9 : add_76208[3:0]]);
  assign add_76246 = array_index_76240[add_76208 > 32'h0000_0009 ? 4'h9 : add_76208[3:0]] + smul_76244;
  assign array_update_76248[0] = add_76208 == 32'h0000_0000 ? add_76246 : array_index_76240[0];
  assign array_update_76248[1] = add_76208 == 32'h0000_0001 ? add_76246 : array_index_76240[1];
  assign array_update_76248[2] = add_76208 == 32'h0000_0002 ? add_76246 : array_index_76240[2];
  assign array_update_76248[3] = add_76208 == 32'h0000_0003 ? add_76246 : array_index_76240[3];
  assign array_update_76248[4] = add_76208 == 32'h0000_0004 ? add_76246 : array_index_76240[4];
  assign array_update_76248[5] = add_76208 == 32'h0000_0005 ? add_76246 : array_index_76240[5];
  assign array_update_76248[6] = add_76208 == 32'h0000_0006 ? add_76246 : array_index_76240[6];
  assign array_update_76248[7] = add_76208 == 32'h0000_0007 ? add_76246 : array_index_76240[7];
  assign array_update_76248[8] = add_76208 == 32'h0000_0008 ? add_76246 : array_index_76240[8];
  assign array_update_76248[9] = add_76208 == 32'h0000_0009 ? add_76246 : array_index_76240[9];
  assign add_76249 = add_76236 + 32'h0000_0001;
  assign array_update_76250[0] = add_76070 == 32'h0000_0000 ? array_update_76248 : array_update_76237[0];
  assign array_update_76250[1] = add_76070 == 32'h0000_0001 ? array_update_76248 : array_update_76237[1];
  assign array_update_76250[2] = add_76070 == 32'h0000_0002 ? array_update_76248 : array_update_76237[2];
  assign array_update_76250[3] = add_76070 == 32'h0000_0003 ? array_update_76248 : array_update_76237[3];
  assign array_update_76250[4] = add_76070 == 32'h0000_0004 ? array_update_76248 : array_update_76237[4];
  assign array_update_76250[5] = add_76070 == 32'h0000_0005 ? array_update_76248 : array_update_76237[5];
  assign array_update_76250[6] = add_76070 == 32'h0000_0006 ? array_update_76248 : array_update_76237[6];
  assign array_update_76250[7] = add_76070 == 32'h0000_0007 ? array_update_76248 : array_update_76237[7];
  assign array_update_76250[8] = add_76070 == 32'h0000_0008 ? array_update_76248 : array_update_76237[8];
  assign array_update_76250[9] = add_76070 == 32'h0000_0009 ? array_update_76248 : array_update_76237[9];
  assign array_index_76252 = array_update_72021[add_76249 > 32'h0000_0009 ? 4'h9 : add_76249[3:0]];
  assign array_index_76253 = array_update_76250[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_76257 = smul32b_32b_x_32b(array_index_76077[add_76249 > 32'h0000_0009 ? 4'h9 : add_76249[3:0]], array_index_76252[add_76208 > 32'h0000_0009 ? 4'h9 : add_76208[3:0]]);
  assign add_76259 = array_index_76253[add_76208 > 32'h0000_0009 ? 4'h9 : add_76208[3:0]] + smul_76257;
  assign array_update_76261[0] = add_76208 == 32'h0000_0000 ? add_76259 : array_index_76253[0];
  assign array_update_76261[1] = add_76208 == 32'h0000_0001 ? add_76259 : array_index_76253[1];
  assign array_update_76261[2] = add_76208 == 32'h0000_0002 ? add_76259 : array_index_76253[2];
  assign array_update_76261[3] = add_76208 == 32'h0000_0003 ? add_76259 : array_index_76253[3];
  assign array_update_76261[4] = add_76208 == 32'h0000_0004 ? add_76259 : array_index_76253[4];
  assign array_update_76261[5] = add_76208 == 32'h0000_0005 ? add_76259 : array_index_76253[5];
  assign array_update_76261[6] = add_76208 == 32'h0000_0006 ? add_76259 : array_index_76253[6];
  assign array_update_76261[7] = add_76208 == 32'h0000_0007 ? add_76259 : array_index_76253[7];
  assign array_update_76261[8] = add_76208 == 32'h0000_0008 ? add_76259 : array_index_76253[8];
  assign array_update_76261[9] = add_76208 == 32'h0000_0009 ? add_76259 : array_index_76253[9];
  assign add_76262 = add_76249 + 32'h0000_0001;
  assign array_update_76263[0] = add_76070 == 32'h0000_0000 ? array_update_76261 : array_update_76250[0];
  assign array_update_76263[1] = add_76070 == 32'h0000_0001 ? array_update_76261 : array_update_76250[1];
  assign array_update_76263[2] = add_76070 == 32'h0000_0002 ? array_update_76261 : array_update_76250[2];
  assign array_update_76263[3] = add_76070 == 32'h0000_0003 ? array_update_76261 : array_update_76250[3];
  assign array_update_76263[4] = add_76070 == 32'h0000_0004 ? array_update_76261 : array_update_76250[4];
  assign array_update_76263[5] = add_76070 == 32'h0000_0005 ? array_update_76261 : array_update_76250[5];
  assign array_update_76263[6] = add_76070 == 32'h0000_0006 ? array_update_76261 : array_update_76250[6];
  assign array_update_76263[7] = add_76070 == 32'h0000_0007 ? array_update_76261 : array_update_76250[7];
  assign array_update_76263[8] = add_76070 == 32'h0000_0008 ? array_update_76261 : array_update_76250[8];
  assign array_update_76263[9] = add_76070 == 32'h0000_0009 ? array_update_76261 : array_update_76250[9];
  assign array_index_76265 = array_update_72021[add_76262 > 32'h0000_0009 ? 4'h9 : add_76262[3:0]];
  assign array_index_76266 = array_update_76263[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_76270 = smul32b_32b_x_32b(array_index_76077[add_76262 > 32'h0000_0009 ? 4'h9 : add_76262[3:0]], array_index_76265[add_76208 > 32'h0000_0009 ? 4'h9 : add_76208[3:0]]);
  assign add_76272 = array_index_76266[add_76208 > 32'h0000_0009 ? 4'h9 : add_76208[3:0]] + smul_76270;
  assign array_update_76274[0] = add_76208 == 32'h0000_0000 ? add_76272 : array_index_76266[0];
  assign array_update_76274[1] = add_76208 == 32'h0000_0001 ? add_76272 : array_index_76266[1];
  assign array_update_76274[2] = add_76208 == 32'h0000_0002 ? add_76272 : array_index_76266[2];
  assign array_update_76274[3] = add_76208 == 32'h0000_0003 ? add_76272 : array_index_76266[3];
  assign array_update_76274[4] = add_76208 == 32'h0000_0004 ? add_76272 : array_index_76266[4];
  assign array_update_76274[5] = add_76208 == 32'h0000_0005 ? add_76272 : array_index_76266[5];
  assign array_update_76274[6] = add_76208 == 32'h0000_0006 ? add_76272 : array_index_76266[6];
  assign array_update_76274[7] = add_76208 == 32'h0000_0007 ? add_76272 : array_index_76266[7];
  assign array_update_76274[8] = add_76208 == 32'h0000_0008 ? add_76272 : array_index_76266[8];
  assign array_update_76274[9] = add_76208 == 32'h0000_0009 ? add_76272 : array_index_76266[9];
  assign add_76275 = add_76262 + 32'h0000_0001;
  assign array_update_76276[0] = add_76070 == 32'h0000_0000 ? array_update_76274 : array_update_76263[0];
  assign array_update_76276[1] = add_76070 == 32'h0000_0001 ? array_update_76274 : array_update_76263[1];
  assign array_update_76276[2] = add_76070 == 32'h0000_0002 ? array_update_76274 : array_update_76263[2];
  assign array_update_76276[3] = add_76070 == 32'h0000_0003 ? array_update_76274 : array_update_76263[3];
  assign array_update_76276[4] = add_76070 == 32'h0000_0004 ? array_update_76274 : array_update_76263[4];
  assign array_update_76276[5] = add_76070 == 32'h0000_0005 ? array_update_76274 : array_update_76263[5];
  assign array_update_76276[6] = add_76070 == 32'h0000_0006 ? array_update_76274 : array_update_76263[6];
  assign array_update_76276[7] = add_76070 == 32'h0000_0007 ? array_update_76274 : array_update_76263[7];
  assign array_update_76276[8] = add_76070 == 32'h0000_0008 ? array_update_76274 : array_update_76263[8];
  assign array_update_76276[9] = add_76070 == 32'h0000_0009 ? array_update_76274 : array_update_76263[9];
  assign array_index_76278 = array_update_72021[add_76275 > 32'h0000_0009 ? 4'h9 : add_76275[3:0]];
  assign array_index_76279 = array_update_76276[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_76283 = smul32b_32b_x_32b(array_index_76077[add_76275 > 32'h0000_0009 ? 4'h9 : add_76275[3:0]], array_index_76278[add_76208 > 32'h0000_0009 ? 4'h9 : add_76208[3:0]]);
  assign add_76285 = array_index_76279[add_76208 > 32'h0000_0009 ? 4'h9 : add_76208[3:0]] + smul_76283;
  assign array_update_76287[0] = add_76208 == 32'h0000_0000 ? add_76285 : array_index_76279[0];
  assign array_update_76287[1] = add_76208 == 32'h0000_0001 ? add_76285 : array_index_76279[1];
  assign array_update_76287[2] = add_76208 == 32'h0000_0002 ? add_76285 : array_index_76279[2];
  assign array_update_76287[3] = add_76208 == 32'h0000_0003 ? add_76285 : array_index_76279[3];
  assign array_update_76287[4] = add_76208 == 32'h0000_0004 ? add_76285 : array_index_76279[4];
  assign array_update_76287[5] = add_76208 == 32'h0000_0005 ? add_76285 : array_index_76279[5];
  assign array_update_76287[6] = add_76208 == 32'h0000_0006 ? add_76285 : array_index_76279[6];
  assign array_update_76287[7] = add_76208 == 32'h0000_0007 ? add_76285 : array_index_76279[7];
  assign array_update_76287[8] = add_76208 == 32'h0000_0008 ? add_76285 : array_index_76279[8];
  assign array_update_76287[9] = add_76208 == 32'h0000_0009 ? add_76285 : array_index_76279[9];
  assign add_76288 = add_76275 + 32'h0000_0001;
  assign array_update_76289[0] = add_76070 == 32'h0000_0000 ? array_update_76287 : array_update_76276[0];
  assign array_update_76289[1] = add_76070 == 32'h0000_0001 ? array_update_76287 : array_update_76276[1];
  assign array_update_76289[2] = add_76070 == 32'h0000_0002 ? array_update_76287 : array_update_76276[2];
  assign array_update_76289[3] = add_76070 == 32'h0000_0003 ? array_update_76287 : array_update_76276[3];
  assign array_update_76289[4] = add_76070 == 32'h0000_0004 ? array_update_76287 : array_update_76276[4];
  assign array_update_76289[5] = add_76070 == 32'h0000_0005 ? array_update_76287 : array_update_76276[5];
  assign array_update_76289[6] = add_76070 == 32'h0000_0006 ? array_update_76287 : array_update_76276[6];
  assign array_update_76289[7] = add_76070 == 32'h0000_0007 ? array_update_76287 : array_update_76276[7];
  assign array_update_76289[8] = add_76070 == 32'h0000_0008 ? array_update_76287 : array_update_76276[8];
  assign array_update_76289[9] = add_76070 == 32'h0000_0009 ? array_update_76287 : array_update_76276[9];
  assign array_index_76291 = array_update_72021[add_76288 > 32'h0000_0009 ? 4'h9 : add_76288[3:0]];
  assign array_index_76292 = array_update_76289[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_76296 = smul32b_32b_x_32b(array_index_76077[add_76288 > 32'h0000_0009 ? 4'h9 : add_76288[3:0]], array_index_76291[add_76208 > 32'h0000_0009 ? 4'h9 : add_76208[3:0]]);
  assign add_76298 = array_index_76292[add_76208 > 32'h0000_0009 ? 4'h9 : add_76208[3:0]] + smul_76296;
  assign array_update_76300[0] = add_76208 == 32'h0000_0000 ? add_76298 : array_index_76292[0];
  assign array_update_76300[1] = add_76208 == 32'h0000_0001 ? add_76298 : array_index_76292[1];
  assign array_update_76300[2] = add_76208 == 32'h0000_0002 ? add_76298 : array_index_76292[2];
  assign array_update_76300[3] = add_76208 == 32'h0000_0003 ? add_76298 : array_index_76292[3];
  assign array_update_76300[4] = add_76208 == 32'h0000_0004 ? add_76298 : array_index_76292[4];
  assign array_update_76300[5] = add_76208 == 32'h0000_0005 ? add_76298 : array_index_76292[5];
  assign array_update_76300[6] = add_76208 == 32'h0000_0006 ? add_76298 : array_index_76292[6];
  assign array_update_76300[7] = add_76208 == 32'h0000_0007 ? add_76298 : array_index_76292[7];
  assign array_update_76300[8] = add_76208 == 32'h0000_0008 ? add_76298 : array_index_76292[8];
  assign array_update_76300[9] = add_76208 == 32'h0000_0009 ? add_76298 : array_index_76292[9];
  assign add_76301 = add_76288 + 32'h0000_0001;
  assign array_update_76302[0] = add_76070 == 32'h0000_0000 ? array_update_76300 : array_update_76289[0];
  assign array_update_76302[1] = add_76070 == 32'h0000_0001 ? array_update_76300 : array_update_76289[1];
  assign array_update_76302[2] = add_76070 == 32'h0000_0002 ? array_update_76300 : array_update_76289[2];
  assign array_update_76302[3] = add_76070 == 32'h0000_0003 ? array_update_76300 : array_update_76289[3];
  assign array_update_76302[4] = add_76070 == 32'h0000_0004 ? array_update_76300 : array_update_76289[4];
  assign array_update_76302[5] = add_76070 == 32'h0000_0005 ? array_update_76300 : array_update_76289[5];
  assign array_update_76302[6] = add_76070 == 32'h0000_0006 ? array_update_76300 : array_update_76289[6];
  assign array_update_76302[7] = add_76070 == 32'h0000_0007 ? array_update_76300 : array_update_76289[7];
  assign array_update_76302[8] = add_76070 == 32'h0000_0008 ? array_update_76300 : array_update_76289[8];
  assign array_update_76302[9] = add_76070 == 32'h0000_0009 ? array_update_76300 : array_update_76289[9];
  assign array_index_76304 = array_update_72021[add_76301 > 32'h0000_0009 ? 4'h9 : add_76301[3:0]];
  assign array_index_76305 = array_update_76302[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_76309 = smul32b_32b_x_32b(array_index_76077[add_76301 > 32'h0000_0009 ? 4'h9 : add_76301[3:0]], array_index_76304[add_76208 > 32'h0000_0009 ? 4'h9 : add_76208[3:0]]);
  assign add_76311 = array_index_76305[add_76208 > 32'h0000_0009 ? 4'h9 : add_76208[3:0]] + smul_76309;
  assign array_update_76313[0] = add_76208 == 32'h0000_0000 ? add_76311 : array_index_76305[0];
  assign array_update_76313[1] = add_76208 == 32'h0000_0001 ? add_76311 : array_index_76305[1];
  assign array_update_76313[2] = add_76208 == 32'h0000_0002 ? add_76311 : array_index_76305[2];
  assign array_update_76313[3] = add_76208 == 32'h0000_0003 ? add_76311 : array_index_76305[3];
  assign array_update_76313[4] = add_76208 == 32'h0000_0004 ? add_76311 : array_index_76305[4];
  assign array_update_76313[5] = add_76208 == 32'h0000_0005 ? add_76311 : array_index_76305[5];
  assign array_update_76313[6] = add_76208 == 32'h0000_0006 ? add_76311 : array_index_76305[6];
  assign array_update_76313[7] = add_76208 == 32'h0000_0007 ? add_76311 : array_index_76305[7];
  assign array_update_76313[8] = add_76208 == 32'h0000_0008 ? add_76311 : array_index_76305[8];
  assign array_update_76313[9] = add_76208 == 32'h0000_0009 ? add_76311 : array_index_76305[9];
  assign add_76314 = add_76301 + 32'h0000_0001;
  assign array_update_76315[0] = add_76070 == 32'h0000_0000 ? array_update_76313 : array_update_76302[0];
  assign array_update_76315[1] = add_76070 == 32'h0000_0001 ? array_update_76313 : array_update_76302[1];
  assign array_update_76315[2] = add_76070 == 32'h0000_0002 ? array_update_76313 : array_update_76302[2];
  assign array_update_76315[3] = add_76070 == 32'h0000_0003 ? array_update_76313 : array_update_76302[3];
  assign array_update_76315[4] = add_76070 == 32'h0000_0004 ? array_update_76313 : array_update_76302[4];
  assign array_update_76315[5] = add_76070 == 32'h0000_0005 ? array_update_76313 : array_update_76302[5];
  assign array_update_76315[6] = add_76070 == 32'h0000_0006 ? array_update_76313 : array_update_76302[6];
  assign array_update_76315[7] = add_76070 == 32'h0000_0007 ? array_update_76313 : array_update_76302[7];
  assign array_update_76315[8] = add_76070 == 32'h0000_0008 ? array_update_76313 : array_update_76302[8];
  assign array_update_76315[9] = add_76070 == 32'h0000_0009 ? array_update_76313 : array_update_76302[9];
  assign array_index_76317 = array_update_72021[add_76314 > 32'h0000_0009 ? 4'h9 : add_76314[3:0]];
  assign array_index_76318 = array_update_76315[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_76322 = smul32b_32b_x_32b(array_index_76077[add_76314 > 32'h0000_0009 ? 4'h9 : add_76314[3:0]], array_index_76317[add_76208 > 32'h0000_0009 ? 4'h9 : add_76208[3:0]]);
  assign add_76324 = array_index_76318[add_76208 > 32'h0000_0009 ? 4'h9 : add_76208[3:0]] + smul_76322;
  assign array_update_76326[0] = add_76208 == 32'h0000_0000 ? add_76324 : array_index_76318[0];
  assign array_update_76326[1] = add_76208 == 32'h0000_0001 ? add_76324 : array_index_76318[1];
  assign array_update_76326[2] = add_76208 == 32'h0000_0002 ? add_76324 : array_index_76318[2];
  assign array_update_76326[3] = add_76208 == 32'h0000_0003 ? add_76324 : array_index_76318[3];
  assign array_update_76326[4] = add_76208 == 32'h0000_0004 ? add_76324 : array_index_76318[4];
  assign array_update_76326[5] = add_76208 == 32'h0000_0005 ? add_76324 : array_index_76318[5];
  assign array_update_76326[6] = add_76208 == 32'h0000_0006 ? add_76324 : array_index_76318[6];
  assign array_update_76326[7] = add_76208 == 32'h0000_0007 ? add_76324 : array_index_76318[7];
  assign array_update_76326[8] = add_76208 == 32'h0000_0008 ? add_76324 : array_index_76318[8];
  assign array_update_76326[9] = add_76208 == 32'h0000_0009 ? add_76324 : array_index_76318[9];
  assign add_76327 = add_76314 + 32'h0000_0001;
  assign array_update_76328[0] = add_76070 == 32'h0000_0000 ? array_update_76326 : array_update_76315[0];
  assign array_update_76328[1] = add_76070 == 32'h0000_0001 ? array_update_76326 : array_update_76315[1];
  assign array_update_76328[2] = add_76070 == 32'h0000_0002 ? array_update_76326 : array_update_76315[2];
  assign array_update_76328[3] = add_76070 == 32'h0000_0003 ? array_update_76326 : array_update_76315[3];
  assign array_update_76328[4] = add_76070 == 32'h0000_0004 ? array_update_76326 : array_update_76315[4];
  assign array_update_76328[5] = add_76070 == 32'h0000_0005 ? array_update_76326 : array_update_76315[5];
  assign array_update_76328[6] = add_76070 == 32'h0000_0006 ? array_update_76326 : array_update_76315[6];
  assign array_update_76328[7] = add_76070 == 32'h0000_0007 ? array_update_76326 : array_update_76315[7];
  assign array_update_76328[8] = add_76070 == 32'h0000_0008 ? array_update_76326 : array_update_76315[8];
  assign array_update_76328[9] = add_76070 == 32'h0000_0009 ? array_update_76326 : array_update_76315[9];
  assign array_index_76330 = array_update_72021[add_76327 > 32'h0000_0009 ? 4'h9 : add_76327[3:0]];
  assign array_index_76331 = array_update_76328[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_76335 = smul32b_32b_x_32b(array_index_76077[add_76327 > 32'h0000_0009 ? 4'h9 : add_76327[3:0]], array_index_76330[add_76208 > 32'h0000_0009 ? 4'h9 : add_76208[3:0]]);
  assign add_76337 = array_index_76331[add_76208 > 32'h0000_0009 ? 4'h9 : add_76208[3:0]] + smul_76335;
  assign array_update_76338[0] = add_76208 == 32'h0000_0000 ? add_76337 : array_index_76331[0];
  assign array_update_76338[1] = add_76208 == 32'h0000_0001 ? add_76337 : array_index_76331[1];
  assign array_update_76338[2] = add_76208 == 32'h0000_0002 ? add_76337 : array_index_76331[2];
  assign array_update_76338[3] = add_76208 == 32'h0000_0003 ? add_76337 : array_index_76331[3];
  assign array_update_76338[4] = add_76208 == 32'h0000_0004 ? add_76337 : array_index_76331[4];
  assign array_update_76338[5] = add_76208 == 32'h0000_0005 ? add_76337 : array_index_76331[5];
  assign array_update_76338[6] = add_76208 == 32'h0000_0006 ? add_76337 : array_index_76331[6];
  assign array_update_76338[7] = add_76208 == 32'h0000_0007 ? add_76337 : array_index_76331[7];
  assign array_update_76338[8] = add_76208 == 32'h0000_0008 ? add_76337 : array_index_76331[8];
  assign array_update_76338[9] = add_76208 == 32'h0000_0009 ? add_76337 : array_index_76331[9];
  assign array_update_76339[0] = add_76070 == 32'h0000_0000 ? array_update_76338 : array_update_76328[0];
  assign array_update_76339[1] = add_76070 == 32'h0000_0001 ? array_update_76338 : array_update_76328[1];
  assign array_update_76339[2] = add_76070 == 32'h0000_0002 ? array_update_76338 : array_update_76328[2];
  assign array_update_76339[3] = add_76070 == 32'h0000_0003 ? array_update_76338 : array_update_76328[3];
  assign array_update_76339[4] = add_76070 == 32'h0000_0004 ? array_update_76338 : array_update_76328[4];
  assign array_update_76339[5] = add_76070 == 32'h0000_0005 ? array_update_76338 : array_update_76328[5];
  assign array_update_76339[6] = add_76070 == 32'h0000_0006 ? array_update_76338 : array_update_76328[6];
  assign array_update_76339[7] = add_76070 == 32'h0000_0007 ? array_update_76338 : array_update_76328[7];
  assign array_update_76339[8] = add_76070 == 32'h0000_0008 ? array_update_76338 : array_update_76328[8];
  assign array_update_76339[9] = add_76070 == 32'h0000_0009 ? array_update_76338 : array_update_76328[9];
  assign array_index_76341 = array_update_76339[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign add_76343 = add_76208 + 32'h0000_0001;
  assign array_update_76344[0] = add_76343 == 32'h0000_0000 ? 32'h0000_0000 : array_index_76341[0];
  assign array_update_76344[1] = add_76343 == 32'h0000_0001 ? 32'h0000_0000 : array_index_76341[1];
  assign array_update_76344[2] = add_76343 == 32'h0000_0002 ? 32'h0000_0000 : array_index_76341[2];
  assign array_update_76344[3] = add_76343 == 32'h0000_0003 ? 32'h0000_0000 : array_index_76341[3];
  assign array_update_76344[4] = add_76343 == 32'h0000_0004 ? 32'h0000_0000 : array_index_76341[4];
  assign array_update_76344[5] = add_76343 == 32'h0000_0005 ? 32'h0000_0000 : array_index_76341[5];
  assign array_update_76344[6] = add_76343 == 32'h0000_0006 ? 32'h0000_0000 : array_index_76341[6];
  assign array_update_76344[7] = add_76343 == 32'h0000_0007 ? 32'h0000_0000 : array_index_76341[7];
  assign array_update_76344[8] = add_76343 == 32'h0000_0008 ? 32'h0000_0000 : array_index_76341[8];
  assign array_update_76344[9] = add_76343 == 32'h0000_0009 ? 32'h0000_0000 : array_index_76341[9];
  assign literal_76345 = 32'h0000_0000;
  assign array_update_76346[0] = add_76070 == 32'h0000_0000 ? array_update_76344 : array_update_76339[0];
  assign array_update_76346[1] = add_76070 == 32'h0000_0001 ? array_update_76344 : array_update_76339[1];
  assign array_update_76346[2] = add_76070 == 32'h0000_0002 ? array_update_76344 : array_update_76339[2];
  assign array_update_76346[3] = add_76070 == 32'h0000_0003 ? array_update_76344 : array_update_76339[3];
  assign array_update_76346[4] = add_76070 == 32'h0000_0004 ? array_update_76344 : array_update_76339[4];
  assign array_update_76346[5] = add_76070 == 32'h0000_0005 ? array_update_76344 : array_update_76339[5];
  assign array_update_76346[6] = add_76070 == 32'h0000_0006 ? array_update_76344 : array_update_76339[6];
  assign array_update_76346[7] = add_76070 == 32'h0000_0007 ? array_update_76344 : array_update_76339[7];
  assign array_update_76346[8] = add_76070 == 32'h0000_0008 ? array_update_76344 : array_update_76339[8];
  assign array_update_76346[9] = add_76070 == 32'h0000_0009 ? array_update_76344 : array_update_76339[9];
  assign array_index_76348 = array_update_72021[literal_76345 > 32'h0000_0009 ? 4'h9 : literal_76345[3:0]];
  assign array_index_76349 = array_update_76346[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_76353 = smul32b_32b_x_32b(array_index_76077[literal_76345 > 32'h0000_0009 ? 4'h9 : literal_76345[3:0]], array_index_76348[add_76343 > 32'h0000_0009 ? 4'h9 : add_76343[3:0]]);
  assign add_76355 = array_index_76349[add_76343 > 32'h0000_0009 ? 4'h9 : add_76343[3:0]] + smul_76353;
  assign array_update_76357[0] = add_76343 == 32'h0000_0000 ? add_76355 : array_index_76349[0];
  assign array_update_76357[1] = add_76343 == 32'h0000_0001 ? add_76355 : array_index_76349[1];
  assign array_update_76357[2] = add_76343 == 32'h0000_0002 ? add_76355 : array_index_76349[2];
  assign array_update_76357[3] = add_76343 == 32'h0000_0003 ? add_76355 : array_index_76349[3];
  assign array_update_76357[4] = add_76343 == 32'h0000_0004 ? add_76355 : array_index_76349[4];
  assign array_update_76357[5] = add_76343 == 32'h0000_0005 ? add_76355 : array_index_76349[5];
  assign array_update_76357[6] = add_76343 == 32'h0000_0006 ? add_76355 : array_index_76349[6];
  assign array_update_76357[7] = add_76343 == 32'h0000_0007 ? add_76355 : array_index_76349[7];
  assign array_update_76357[8] = add_76343 == 32'h0000_0008 ? add_76355 : array_index_76349[8];
  assign array_update_76357[9] = add_76343 == 32'h0000_0009 ? add_76355 : array_index_76349[9];
  assign add_76358 = literal_76345 + 32'h0000_0001;
  assign array_update_76359[0] = add_76070 == 32'h0000_0000 ? array_update_76357 : array_update_76346[0];
  assign array_update_76359[1] = add_76070 == 32'h0000_0001 ? array_update_76357 : array_update_76346[1];
  assign array_update_76359[2] = add_76070 == 32'h0000_0002 ? array_update_76357 : array_update_76346[2];
  assign array_update_76359[3] = add_76070 == 32'h0000_0003 ? array_update_76357 : array_update_76346[3];
  assign array_update_76359[4] = add_76070 == 32'h0000_0004 ? array_update_76357 : array_update_76346[4];
  assign array_update_76359[5] = add_76070 == 32'h0000_0005 ? array_update_76357 : array_update_76346[5];
  assign array_update_76359[6] = add_76070 == 32'h0000_0006 ? array_update_76357 : array_update_76346[6];
  assign array_update_76359[7] = add_76070 == 32'h0000_0007 ? array_update_76357 : array_update_76346[7];
  assign array_update_76359[8] = add_76070 == 32'h0000_0008 ? array_update_76357 : array_update_76346[8];
  assign array_update_76359[9] = add_76070 == 32'h0000_0009 ? array_update_76357 : array_update_76346[9];
  assign array_index_76361 = array_update_72021[add_76358 > 32'h0000_0009 ? 4'h9 : add_76358[3:0]];
  assign array_index_76362 = array_update_76359[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_76366 = smul32b_32b_x_32b(array_index_76077[add_76358 > 32'h0000_0009 ? 4'h9 : add_76358[3:0]], array_index_76361[add_76343 > 32'h0000_0009 ? 4'h9 : add_76343[3:0]]);
  assign add_76368 = array_index_76362[add_76343 > 32'h0000_0009 ? 4'h9 : add_76343[3:0]] + smul_76366;
  assign array_update_76370[0] = add_76343 == 32'h0000_0000 ? add_76368 : array_index_76362[0];
  assign array_update_76370[1] = add_76343 == 32'h0000_0001 ? add_76368 : array_index_76362[1];
  assign array_update_76370[2] = add_76343 == 32'h0000_0002 ? add_76368 : array_index_76362[2];
  assign array_update_76370[3] = add_76343 == 32'h0000_0003 ? add_76368 : array_index_76362[3];
  assign array_update_76370[4] = add_76343 == 32'h0000_0004 ? add_76368 : array_index_76362[4];
  assign array_update_76370[5] = add_76343 == 32'h0000_0005 ? add_76368 : array_index_76362[5];
  assign array_update_76370[6] = add_76343 == 32'h0000_0006 ? add_76368 : array_index_76362[6];
  assign array_update_76370[7] = add_76343 == 32'h0000_0007 ? add_76368 : array_index_76362[7];
  assign array_update_76370[8] = add_76343 == 32'h0000_0008 ? add_76368 : array_index_76362[8];
  assign array_update_76370[9] = add_76343 == 32'h0000_0009 ? add_76368 : array_index_76362[9];
  assign add_76371 = add_76358 + 32'h0000_0001;
  assign array_update_76372[0] = add_76070 == 32'h0000_0000 ? array_update_76370 : array_update_76359[0];
  assign array_update_76372[1] = add_76070 == 32'h0000_0001 ? array_update_76370 : array_update_76359[1];
  assign array_update_76372[2] = add_76070 == 32'h0000_0002 ? array_update_76370 : array_update_76359[2];
  assign array_update_76372[3] = add_76070 == 32'h0000_0003 ? array_update_76370 : array_update_76359[3];
  assign array_update_76372[4] = add_76070 == 32'h0000_0004 ? array_update_76370 : array_update_76359[4];
  assign array_update_76372[5] = add_76070 == 32'h0000_0005 ? array_update_76370 : array_update_76359[5];
  assign array_update_76372[6] = add_76070 == 32'h0000_0006 ? array_update_76370 : array_update_76359[6];
  assign array_update_76372[7] = add_76070 == 32'h0000_0007 ? array_update_76370 : array_update_76359[7];
  assign array_update_76372[8] = add_76070 == 32'h0000_0008 ? array_update_76370 : array_update_76359[8];
  assign array_update_76372[9] = add_76070 == 32'h0000_0009 ? array_update_76370 : array_update_76359[9];
  assign array_index_76374 = array_update_72021[add_76371 > 32'h0000_0009 ? 4'h9 : add_76371[3:0]];
  assign array_index_76375 = array_update_76372[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_76379 = smul32b_32b_x_32b(array_index_76077[add_76371 > 32'h0000_0009 ? 4'h9 : add_76371[3:0]], array_index_76374[add_76343 > 32'h0000_0009 ? 4'h9 : add_76343[3:0]]);
  assign add_76381 = array_index_76375[add_76343 > 32'h0000_0009 ? 4'h9 : add_76343[3:0]] + smul_76379;
  assign array_update_76383[0] = add_76343 == 32'h0000_0000 ? add_76381 : array_index_76375[0];
  assign array_update_76383[1] = add_76343 == 32'h0000_0001 ? add_76381 : array_index_76375[1];
  assign array_update_76383[2] = add_76343 == 32'h0000_0002 ? add_76381 : array_index_76375[2];
  assign array_update_76383[3] = add_76343 == 32'h0000_0003 ? add_76381 : array_index_76375[3];
  assign array_update_76383[4] = add_76343 == 32'h0000_0004 ? add_76381 : array_index_76375[4];
  assign array_update_76383[5] = add_76343 == 32'h0000_0005 ? add_76381 : array_index_76375[5];
  assign array_update_76383[6] = add_76343 == 32'h0000_0006 ? add_76381 : array_index_76375[6];
  assign array_update_76383[7] = add_76343 == 32'h0000_0007 ? add_76381 : array_index_76375[7];
  assign array_update_76383[8] = add_76343 == 32'h0000_0008 ? add_76381 : array_index_76375[8];
  assign array_update_76383[9] = add_76343 == 32'h0000_0009 ? add_76381 : array_index_76375[9];
  assign add_76384 = add_76371 + 32'h0000_0001;
  assign array_update_76385[0] = add_76070 == 32'h0000_0000 ? array_update_76383 : array_update_76372[0];
  assign array_update_76385[1] = add_76070 == 32'h0000_0001 ? array_update_76383 : array_update_76372[1];
  assign array_update_76385[2] = add_76070 == 32'h0000_0002 ? array_update_76383 : array_update_76372[2];
  assign array_update_76385[3] = add_76070 == 32'h0000_0003 ? array_update_76383 : array_update_76372[3];
  assign array_update_76385[4] = add_76070 == 32'h0000_0004 ? array_update_76383 : array_update_76372[4];
  assign array_update_76385[5] = add_76070 == 32'h0000_0005 ? array_update_76383 : array_update_76372[5];
  assign array_update_76385[6] = add_76070 == 32'h0000_0006 ? array_update_76383 : array_update_76372[6];
  assign array_update_76385[7] = add_76070 == 32'h0000_0007 ? array_update_76383 : array_update_76372[7];
  assign array_update_76385[8] = add_76070 == 32'h0000_0008 ? array_update_76383 : array_update_76372[8];
  assign array_update_76385[9] = add_76070 == 32'h0000_0009 ? array_update_76383 : array_update_76372[9];
  assign array_index_76387 = array_update_72021[add_76384 > 32'h0000_0009 ? 4'h9 : add_76384[3:0]];
  assign array_index_76388 = array_update_76385[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_76392 = smul32b_32b_x_32b(array_index_76077[add_76384 > 32'h0000_0009 ? 4'h9 : add_76384[3:0]], array_index_76387[add_76343 > 32'h0000_0009 ? 4'h9 : add_76343[3:0]]);
  assign add_76394 = array_index_76388[add_76343 > 32'h0000_0009 ? 4'h9 : add_76343[3:0]] + smul_76392;
  assign array_update_76396[0] = add_76343 == 32'h0000_0000 ? add_76394 : array_index_76388[0];
  assign array_update_76396[1] = add_76343 == 32'h0000_0001 ? add_76394 : array_index_76388[1];
  assign array_update_76396[2] = add_76343 == 32'h0000_0002 ? add_76394 : array_index_76388[2];
  assign array_update_76396[3] = add_76343 == 32'h0000_0003 ? add_76394 : array_index_76388[3];
  assign array_update_76396[4] = add_76343 == 32'h0000_0004 ? add_76394 : array_index_76388[4];
  assign array_update_76396[5] = add_76343 == 32'h0000_0005 ? add_76394 : array_index_76388[5];
  assign array_update_76396[6] = add_76343 == 32'h0000_0006 ? add_76394 : array_index_76388[6];
  assign array_update_76396[7] = add_76343 == 32'h0000_0007 ? add_76394 : array_index_76388[7];
  assign array_update_76396[8] = add_76343 == 32'h0000_0008 ? add_76394 : array_index_76388[8];
  assign array_update_76396[9] = add_76343 == 32'h0000_0009 ? add_76394 : array_index_76388[9];
  assign add_76397 = add_76384 + 32'h0000_0001;
  assign array_update_76398[0] = add_76070 == 32'h0000_0000 ? array_update_76396 : array_update_76385[0];
  assign array_update_76398[1] = add_76070 == 32'h0000_0001 ? array_update_76396 : array_update_76385[1];
  assign array_update_76398[2] = add_76070 == 32'h0000_0002 ? array_update_76396 : array_update_76385[2];
  assign array_update_76398[3] = add_76070 == 32'h0000_0003 ? array_update_76396 : array_update_76385[3];
  assign array_update_76398[4] = add_76070 == 32'h0000_0004 ? array_update_76396 : array_update_76385[4];
  assign array_update_76398[5] = add_76070 == 32'h0000_0005 ? array_update_76396 : array_update_76385[5];
  assign array_update_76398[6] = add_76070 == 32'h0000_0006 ? array_update_76396 : array_update_76385[6];
  assign array_update_76398[7] = add_76070 == 32'h0000_0007 ? array_update_76396 : array_update_76385[7];
  assign array_update_76398[8] = add_76070 == 32'h0000_0008 ? array_update_76396 : array_update_76385[8];
  assign array_update_76398[9] = add_76070 == 32'h0000_0009 ? array_update_76396 : array_update_76385[9];
  assign array_index_76400 = array_update_72021[add_76397 > 32'h0000_0009 ? 4'h9 : add_76397[3:0]];
  assign array_index_76401 = array_update_76398[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_76405 = smul32b_32b_x_32b(array_index_76077[add_76397 > 32'h0000_0009 ? 4'h9 : add_76397[3:0]], array_index_76400[add_76343 > 32'h0000_0009 ? 4'h9 : add_76343[3:0]]);
  assign add_76407 = array_index_76401[add_76343 > 32'h0000_0009 ? 4'h9 : add_76343[3:0]] + smul_76405;
  assign array_update_76409[0] = add_76343 == 32'h0000_0000 ? add_76407 : array_index_76401[0];
  assign array_update_76409[1] = add_76343 == 32'h0000_0001 ? add_76407 : array_index_76401[1];
  assign array_update_76409[2] = add_76343 == 32'h0000_0002 ? add_76407 : array_index_76401[2];
  assign array_update_76409[3] = add_76343 == 32'h0000_0003 ? add_76407 : array_index_76401[3];
  assign array_update_76409[4] = add_76343 == 32'h0000_0004 ? add_76407 : array_index_76401[4];
  assign array_update_76409[5] = add_76343 == 32'h0000_0005 ? add_76407 : array_index_76401[5];
  assign array_update_76409[6] = add_76343 == 32'h0000_0006 ? add_76407 : array_index_76401[6];
  assign array_update_76409[7] = add_76343 == 32'h0000_0007 ? add_76407 : array_index_76401[7];
  assign array_update_76409[8] = add_76343 == 32'h0000_0008 ? add_76407 : array_index_76401[8];
  assign array_update_76409[9] = add_76343 == 32'h0000_0009 ? add_76407 : array_index_76401[9];
  assign add_76410 = add_76397 + 32'h0000_0001;
  assign array_update_76411[0] = add_76070 == 32'h0000_0000 ? array_update_76409 : array_update_76398[0];
  assign array_update_76411[1] = add_76070 == 32'h0000_0001 ? array_update_76409 : array_update_76398[1];
  assign array_update_76411[2] = add_76070 == 32'h0000_0002 ? array_update_76409 : array_update_76398[2];
  assign array_update_76411[3] = add_76070 == 32'h0000_0003 ? array_update_76409 : array_update_76398[3];
  assign array_update_76411[4] = add_76070 == 32'h0000_0004 ? array_update_76409 : array_update_76398[4];
  assign array_update_76411[5] = add_76070 == 32'h0000_0005 ? array_update_76409 : array_update_76398[5];
  assign array_update_76411[6] = add_76070 == 32'h0000_0006 ? array_update_76409 : array_update_76398[6];
  assign array_update_76411[7] = add_76070 == 32'h0000_0007 ? array_update_76409 : array_update_76398[7];
  assign array_update_76411[8] = add_76070 == 32'h0000_0008 ? array_update_76409 : array_update_76398[8];
  assign array_update_76411[9] = add_76070 == 32'h0000_0009 ? array_update_76409 : array_update_76398[9];
  assign array_index_76413 = array_update_72021[add_76410 > 32'h0000_0009 ? 4'h9 : add_76410[3:0]];
  assign array_index_76414 = array_update_76411[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_76418 = smul32b_32b_x_32b(array_index_76077[add_76410 > 32'h0000_0009 ? 4'h9 : add_76410[3:0]], array_index_76413[add_76343 > 32'h0000_0009 ? 4'h9 : add_76343[3:0]]);
  assign add_76420 = array_index_76414[add_76343 > 32'h0000_0009 ? 4'h9 : add_76343[3:0]] + smul_76418;
  assign array_update_76422[0] = add_76343 == 32'h0000_0000 ? add_76420 : array_index_76414[0];
  assign array_update_76422[1] = add_76343 == 32'h0000_0001 ? add_76420 : array_index_76414[1];
  assign array_update_76422[2] = add_76343 == 32'h0000_0002 ? add_76420 : array_index_76414[2];
  assign array_update_76422[3] = add_76343 == 32'h0000_0003 ? add_76420 : array_index_76414[3];
  assign array_update_76422[4] = add_76343 == 32'h0000_0004 ? add_76420 : array_index_76414[4];
  assign array_update_76422[5] = add_76343 == 32'h0000_0005 ? add_76420 : array_index_76414[5];
  assign array_update_76422[6] = add_76343 == 32'h0000_0006 ? add_76420 : array_index_76414[6];
  assign array_update_76422[7] = add_76343 == 32'h0000_0007 ? add_76420 : array_index_76414[7];
  assign array_update_76422[8] = add_76343 == 32'h0000_0008 ? add_76420 : array_index_76414[8];
  assign array_update_76422[9] = add_76343 == 32'h0000_0009 ? add_76420 : array_index_76414[9];
  assign add_76423 = add_76410 + 32'h0000_0001;
  assign array_update_76424[0] = add_76070 == 32'h0000_0000 ? array_update_76422 : array_update_76411[0];
  assign array_update_76424[1] = add_76070 == 32'h0000_0001 ? array_update_76422 : array_update_76411[1];
  assign array_update_76424[2] = add_76070 == 32'h0000_0002 ? array_update_76422 : array_update_76411[2];
  assign array_update_76424[3] = add_76070 == 32'h0000_0003 ? array_update_76422 : array_update_76411[3];
  assign array_update_76424[4] = add_76070 == 32'h0000_0004 ? array_update_76422 : array_update_76411[4];
  assign array_update_76424[5] = add_76070 == 32'h0000_0005 ? array_update_76422 : array_update_76411[5];
  assign array_update_76424[6] = add_76070 == 32'h0000_0006 ? array_update_76422 : array_update_76411[6];
  assign array_update_76424[7] = add_76070 == 32'h0000_0007 ? array_update_76422 : array_update_76411[7];
  assign array_update_76424[8] = add_76070 == 32'h0000_0008 ? array_update_76422 : array_update_76411[8];
  assign array_update_76424[9] = add_76070 == 32'h0000_0009 ? array_update_76422 : array_update_76411[9];
  assign array_index_76426 = array_update_72021[add_76423 > 32'h0000_0009 ? 4'h9 : add_76423[3:0]];
  assign array_index_76427 = array_update_76424[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_76431 = smul32b_32b_x_32b(array_index_76077[add_76423 > 32'h0000_0009 ? 4'h9 : add_76423[3:0]], array_index_76426[add_76343 > 32'h0000_0009 ? 4'h9 : add_76343[3:0]]);
  assign add_76433 = array_index_76427[add_76343 > 32'h0000_0009 ? 4'h9 : add_76343[3:0]] + smul_76431;
  assign array_update_76435[0] = add_76343 == 32'h0000_0000 ? add_76433 : array_index_76427[0];
  assign array_update_76435[1] = add_76343 == 32'h0000_0001 ? add_76433 : array_index_76427[1];
  assign array_update_76435[2] = add_76343 == 32'h0000_0002 ? add_76433 : array_index_76427[2];
  assign array_update_76435[3] = add_76343 == 32'h0000_0003 ? add_76433 : array_index_76427[3];
  assign array_update_76435[4] = add_76343 == 32'h0000_0004 ? add_76433 : array_index_76427[4];
  assign array_update_76435[5] = add_76343 == 32'h0000_0005 ? add_76433 : array_index_76427[5];
  assign array_update_76435[6] = add_76343 == 32'h0000_0006 ? add_76433 : array_index_76427[6];
  assign array_update_76435[7] = add_76343 == 32'h0000_0007 ? add_76433 : array_index_76427[7];
  assign array_update_76435[8] = add_76343 == 32'h0000_0008 ? add_76433 : array_index_76427[8];
  assign array_update_76435[9] = add_76343 == 32'h0000_0009 ? add_76433 : array_index_76427[9];
  assign add_76436 = add_76423 + 32'h0000_0001;
  assign array_update_76437[0] = add_76070 == 32'h0000_0000 ? array_update_76435 : array_update_76424[0];
  assign array_update_76437[1] = add_76070 == 32'h0000_0001 ? array_update_76435 : array_update_76424[1];
  assign array_update_76437[2] = add_76070 == 32'h0000_0002 ? array_update_76435 : array_update_76424[2];
  assign array_update_76437[3] = add_76070 == 32'h0000_0003 ? array_update_76435 : array_update_76424[3];
  assign array_update_76437[4] = add_76070 == 32'h0000_0004 ? array_update_76435 : array_update_76424[4];
  assign array_update_76437[5] = add_76070 == 32'h0000_0005 ? array_update_76435 : array_update_76424[5];
  assign array_update_76437[6] = add_76070 == 32'h0000_0006 ? array_update_76435 : array_update_76424[6];
  assign array_update_76437[7] = add_76070 == 32'h0000_0007 ? array_update_76435 : array_update_76424[7];
  assign array_update_76437[8] = add_76070 == 32'h0000_0008 ? array_update_76435 : array_update_76424[8];
  assign array_update_76437[9] = add_76070 == 32'h0000_0009 ? array_update_76435 : array_update_76424[9];
  assign array_index_76439 = array_update_72021[add_76436 > 32'h0000_0009 ? 4'h9 : add_76436[3:0]];
  assign array_index_76440 = array_update_76437[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_76444 = smul32b_32b_x_32b(array_index_76077[add_76436 > 32'h0000_0009 ? 4'h9 : add_76436[3:0]], array_index_76439[add_76343 > 32'h0000_0009 ? 4'h9 : add_76343[3:0]]);
  assign add_76446 = array_index_76440[add_76343 > 32'h0000_0009 ? 4'h9 : add_76343[3:0]] + smul_76444;
  assign array_update_76448[0] = add_76343 == 32'h0000_0000 ? add_76446 : array_index_76440[0];
  assign array_update_76448[1] = add_76343 == 32'h0000_0001 ? add_76446 : array_index_76440[1];
  assign array_update_76448[2] = add_76343 == 32'h0000_0002 ? add_76446 : array_index_76440[2];
  assign array_update_76448[3] = add_76343 == 32'h0000_0003 ? add_76446 : array_index_76440[3];
  assign array_update_76448[4] = add_76343 == 32'h0000_0004 ? add_76446 : array_index_76440[4];
  assign array_update_76448[5] = add_76343 == 32'h0000_0005 ? add_76446 : array_index_76440[5];
  assign array_update_76448[6] = add_76343 == 32'h0000_0006 ? add_76446 : array_index_76440[6];
  assign array_update_76448[7] = add_76343 == 32'h0000_0007 ? add_76446 : array_index_76440[7];
  assign array_update_76448[8] = add_76343 == 32'h0000_0008 ? add_76446 : array_index_76440[8];
  assign array_update_76448[9] = add_76343 == 32'h0000_0009 ? add_76446 : array_index_76440[9];
  assign add_76449 = add_76436 + 32'h0000_0001;
  assign array_update_76450[0] = add_76070 == 32'h0000_0000 ? array_update_76448 : array_update_76437[0];
  assign array_update_76450[1] = add_76070 == 32'h0000_0001 ? array_update_76448 : array_update_76437[1];
  assign array_update_76450[2] = add_76070 == 32'h0000_0002 ? array_update_76448 : array_update_76437[2];
  assign array_update_76450[3] = add_76070 == 32'h0000_0003 ? array_update_76448 : array_update_76437[3];
  assign array_update_76450[4] = add_76070 == 32'h0000_0004 ? array_update_76448 : array_update_76437[4];
  assign array_update_76450[5] = add_76070 == 32'h0000_0005 ? array_update_76448 : array_update_76437[5];
  assign array_update_76450[6] = add_76070 == 32'h0000_0006 ? array_update_76448 : array_update_76437[6];
  assign array_update_76450[7] = add_76070 == 32'h0000_0007 ? array_update_76448 : array_update_76437[7];
  assign array_update_76450[8] = add_76070 == 32'h0000_0008 ? array_update_76448 : array_update_76437[8];
  assign array_update_76450[9] = add_76070 == 32'h0000_0009 ? array_update_76448 : array_update_76437[9];
  assign array_index_76452 = array_update_72021[add_76449 > 32'h0000_0009 ? 4'h9 : add_76449[3:0]];
  assign array_index_76453 = array_update_76450[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_76457 = smul32b_32b_x_32b(array_index_76077[add_76449 > 32'h0000_0009 ? 4'h9 : add_76449[3:0]], array_index_76452[add_76343 > 32'h0000_0009 ? 4'h9 : add_76343[3:0]]);
  assign add_76459 = array_index_76453[add_76343 > 32'h0000_0009 ? 4'h9 : add_76343[3:0]] + smul_76457;
  assign array_update_76461[0] = add_76343 == 32'h0000_0000 ? add_76459 : array_index_76453[0];
  assign array_update_76461[1] = add_76343 == 32'h0000_0001 ? add_76459 : array_index_76453[1];
  assign array_update_76461[2] = add_76343 == 32'h0000_0002 ? add_76459 : array_index_76453[2];
  assign array_update_76461[3] = add_76343 == 32'h0000_0003 ? add_76459 : array_index_76453[3];
  assign array_update_76461[4] = add_76343 == 32'h0000_0004 ? add_76459 : array_index_76453[4];
  assign array_update_76461[5] = add_76343 == 32'h0000_0005 ? add_76459 : array_index_76453[5];
  assign array_update_76461[6] = add_76343 == 32'h0000_0006 ? add_76459 : array_index_76453[6];
  assign array_update_76461[7] = add_76343 == 32'h0000_0007 ? add_76459 : array_index_76453[7];
  assign array_update_76461[8] = add_76343 == 32'h0000_0008 ? add_76459 : array_index_76453[8];
  assign array_update_76461[9] = add_76343 == 32'h0000_0009 ? add_76459 : array_index_76453[9];
  assign add_76462 = add_76449 + 32'h0000_0001;
  assign array_update_76463[0] = add_76070 == 32'h0000_0000 ? array_update_76461 : array_update_76450[0];
  assign array_update_76463[1] = add_76070 == 32'h0000_0001 ? array_update_76461 : array_update_76450[1];
  assign array_update_76463[2] = add_76070 == 32'h0000_0002 ? array_update_76461 : array_update_76450[2];
  assign array_update_76463[3] = add_76070 == 32'h0000_0003 ? array_update_76461 : array_update_76450[3];
  assign array_update_76463[4] = add_76070 == 32'h0000_0004 ? array_update_76461 : array_update_76450[4];
  assign array_update_76463[5] = add_76070 == 32'h0000_0005 ? array_update_76461 : array_update_76450[5];
  assign array_update_76463[6] = add_76070 == 32'h0000_0006 ? array_update_76461 : array_update_76450[6];
  assign array_update_76463[7] = add_76070 == 32'h0000_0007 ? array_update_76461 : array_update_76450[7];
  assign array_update_76463[8] = add_76070 == 32'h0000_0008 ? array_update_76461 : array_update_76450[8];
  assign array_update_76463[9] = add_76070 == 32'h0000_0009 ? array_update_76461 : array_update_76450[9];
  assign array_index_76465 = array_update_72021[add_76462 > 32'h0000_0009 ? 4'h9 : add_76462[3:0]];
  assign array_index_76466 = array_update_76463[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_76470 = smul32b_32b_x_32b(array_index_76077[add_76462 > 32'h0000_0009 ? 4'h9 : add_76462[3:0]], array_index_76465[add_76343 > 32'h0000_0009 ? 4'h9 : add_76343[3:0]]);
  assign add_76472 = array_index_76466[add_76343 > 32'h0000_0009 ? 4'h9 : add_76343[3:0]] + smul_76470;
  assign array_update_76473[0] = add_76343 == 32'h0000_0000 ? add_76472 : array_index_76466[0];
  assign array_update_76473[1] = add_76343 == 32'h0000_0001 ? add_76472 : array_index_76466[1];
  assign array_update_76473[2] = add_76343 == 32'h0000_0002 ? add_76472 : array_index_76466[2];
  assign array_update_76473[3] = add_76343 == 32'h0000_0003 ? add_76472 : array_index_76466[3];
  assign array_update_76473[4] = add_76343 == 32'h0000_0004 ? add_76472 : array_index_76466[4];
  assign array_update_76473[5] = add_76343 == 32'h0000_0005 ? add_76472 : array_index_76466[5];
  assign array_update_76473[6] = add_76343 == 32'h0000_0006 ? add_76472 : array_index_76466[6];
  assign array_update_76473[7] = add_76343 == 32'h0000_0007 ? add_76472 : array_index_76466[7];
  assign array_update_76473[8] = add_76343 == 32'h0000_0008 ? add_76472 : array_index_76466[8];
  assign array_update_76473[9] = add_76343 == 32'h0000_0009 ? add_76472 : array_index_76466[9];
  assign array_update_76474[0] = add_76070 == 32'h0000_0000 ? array_update_76473 : array_update_76463[0];
  assign array_update_76474[1] = add_76070 == 32'h0000_0001 ? array_update_76473 : array_update_76463[1];
  assign array_update_76474[2] = add_76070 == 32'h0000_0002 ? array_update_76473 : array_update_76463[2];
  assign array_update_76474[3] = add_76070 == 32'h0000_0003 ? array_update_76473 : array_update_76463[3];
  assign array_update_76474[4] = add_76070 == 32'h0000_0004 ? array_update_76473 : array_update_76463[4];
  assign array_update_76474[5] = add_76070 == 32'h0000_0005 ? array_update_76473 : array_update_76463[5];
  assign array_update_76474[6] = add_76070 == 32'h0000_0006 ? array_update_76473 : array_update_76463[6];
  assign array_update_76474[7] = add_76070 == 32'h0000_0007 ? array_update_76473 : array_update_76463[7];
  assign array_update_76474[8] = add_76070 == 32'h0000_0008 ? array_update_76473 : array_update_76463[8];
  assign array_update_76474[9] = add_76070 == 32'h0000_0009 ? array_update_76473 : array_update_76463[9];
  assign array_index_76476 = array_update_76474[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign add_76478 = add_76343 + 32'h0000_0001;
  assign array_update_76479[0] = add_76478 == 32'h0000_0000 ? 32'h0000_0000 : array_index_76476[0];
  assign array_update_76479[1] = add_76478 == 32'h0000_0001 ? 32'h0000_0000 : array_index_76476[1];
  assign array_update_76479[2] = add_76478 == 32'h0000_0002 ? 32'h0000_0000 : array_index_76476[2];
  assign array_update_76479[3] = add_76478 == 32'h0000_0003 ? 32'h0000_0000 : array_index_76476[3];
  assign array_update_76479[4] = add_76478 == 32'h0000_0004 ? 32'h0000_0000 : array_index_76476[4];
  assign array_update_76479[5] = add_76478 == 32'h0000_0005 ? 32'h0000_0000 : array_index_76476[5];
  assign array_update_76479[6] = add_76478 == 32'h0000_0006 ? 32'h0000_0000 : array_index_76476[6];
  assign array_update_76479[7] = add_76478 == 32'h0000_0007 ? 32'h0000_0000 : array_index_76476[7];
  assign array_update_76479[8] = add_76478 == 32'h0000_0008 ? 32'h0000_0000 : array_index_76476[8];
  assign array_update_76479[9] = add_76478 == 32'h0000_0009 ? 32'h0000_0000 : array_index_76476[9];
  assign literal_76480 = 32'h0000_0000;
  assign array_update_76481[0] = add_76070 == 32'h0000_0000 ? array_update_76479 : array_update_76474[0];
  assign array_update_76481[1] = add_76070 == 32'h0000_0001 ? array_update_76479 : array_update_76474[1];
  assign array_update_76481[2] = add_76070 == 32'h0000_0002 ? array_update_76479 : array_update_76474[2];
  assign array_update_76481[3] = add_76070 == 32'h0000_0003 ? array_update_76479 : array_update_76474[3];
  assign array_update_76481[4] = add_76070 == 32'h0000_0004 ? array_update_76479 : array_update_76474[4];
  assign array_update_76481[5] = add_76070 == 32'h0000_0005 ? array_update_76479 : array_update_76474[5];
  assign array_update_76481[6] = add_76070 == 32'h0000_0006 ? array_update_76479 : array_update_76474[6];
  assign array_update_76481[7] = add_76070 == 32'h0000_0007 ? array_update_76479 : array_update_76474[7];
  assign array_update_76481[8] = add_76070 == 32'h0000_0008 ? array_update_76479 : array_update_76474[8];
  assign array_update_76481[9] = add_76070 == 32'h0000_0009 ? array_update_76479 : array_update_76474[9];
  assign array_index_76483 = array_update_72021[literal_76480 > 32'h0000_0009 ? 4'h9 : literal_76480[3:0]];
  assign array_index_76484 = array_update_76481[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_76488 = smul32b_32b_x_32b(array_index_76077[literal_76480 > 32'h0000_0009 ? 4'h9 : literal_76480[3:0]], array_index_76483[add_76478 > 32'h0000_0009 ? 4'h9 : add_76478[3:0]]);
  assign add_76490 = array_index_76484[add_76478 > 32'h0000_0009 ? 4'h9 : add_76478[3:0]] + smul_76488;
  assign array_update_76492[0] = add_76478 == 32'h0000_0000 ? add_76490 : array_index_76484[0];
  assign array_update_76492[1] = add_76478 == 32'h0000_0001 ? add_76490 : array_index_76484[1];
  assign array_update_76492[2] = add_76478 == 32'h0000_0002 ? add_76490 : array_index_76484[2];
  assign array_update_76492[3] = add_76478 == 32'h0000_0003 ? add_76490 : array_index_76484[3];
  assign array_update_76492[4] = add_76478 == 32'h0000_0004 ? add_76490 : array_index_76484[4];
  assign array_update_76492[5] = add_76478 == 32'h0000_0005 ? add_76490 : array_index_76484[5];
  assign array_update_76492[6] = add_76478 == 32'h0000_0006 ? add_76490 : array_index_76484[6];
  assign array_update_76492[7] = add_76478 == 32'h0000_0007 ? add_76490 : array_index_76484[7];
  assign array_update_76492[8] = add_76478 == 32'h0000_0008 ? add_76490 : array_index_76484[8];
  assign array_update_76492[9] = add_76478 == 32'h0000_0009 ? add_76490 : array_index_76484[9];
  assign add_76493 = literal_76480 + 32'h0000_0001;
  assign array_update_76494[0] = add_76070 == 32'h0000_0000 ? array_update_76492 : array_update_76481[0];
  assign array_update_76494[1] = add_76070 == 32'h0000_0001 ? array_update_76492 : array_update_76481[1];
  assign array_update_76494[2] = add_76070 == 32'h0000_0002 ? array_update_76492 : array_update_76481[2];
  assign array_update_76494[3] = add_76070 == 32'h0000_0003 ? array_update_76492 : array_update_76481[3];
  assign array_update_76494[4] = add_76070 == 32'h0000_0004 ? array_update_76492 : array_update_76481[4];
  assign array_update_76494[5] = add_76070 == 32'h0000_0005 ? array_update_76492 : array_update_76481[5];
  assign array_update_76494[6] = add_76070 == 32'h0000_0006 ? array_update_76492 : array_update_76481[6];
  assign array_update_76494[7] = add_76070 == 32'h0000_0007 ? array_update_76492 : array_update_76481[7];
  assign array_update_76494[8] = add_76070 == 32'h0000_0008 ? array_update_76492 : array_update_76481[8];
  assign array_update_76494[9] = add_76070 == 32'h0000_0009 ? array_update_76492 : array_update_76481[9];
  assign array_index_76496 = array_update_72021[add_76493 > 32'h0000_0009 ? 4'h9 : add_76493[3:0]];
  assign array_index_76497 = array_update_76494[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_76501 = smul32b_32b_x_32b(array_index_76077[add_76493 > 32'h0000_0009 ? 4'h9 : add_76493[3:0]], array_index_76496[add_76478 > 32'h0000_0009 ? 4'h9 : add_76478[3:0]]);
  assign add_76503 = array_index_76497[add_76478 > 32'h0000_0009 ? 4'h9 : add_76478[3:0]] + smul_76501;
  assign array_update_76505[0] = add_76478 == 32'h0000_0000 ? add_76503 : array_index_76497[0];
  assign array_update_76505[1] = add_76478 == 32'h0000_0001 ? add_76503 : array_index_76497[1];
  assign array_update_76505[2] = add_76478 == 32'h0000_0002 ? add_76503 : array_index_76497[2];
  assign array_update_76505[3] = add_76478 == 32'h0000_0003 ? add_76503 : array_index_76497[3];
  assign array_update_76505[4] = add_76478 == 32'h0000_0004 ? add_76503 : array_index_76497[4];
  assign array_update_76505[5] = add_76478 == 32'h0000_0005 ? add_76503 : array_index_76497[5];
  assign array_update_76505[6] = add_76478 == 32'h0000_0006 ? add_76503 : array_index_76497[6];
  assign array_update_76505[7] = add_76478 == 32'h0000_0007 ? add_76503 : array_index_76497[7];
  assign array_update_76505[8] = add_76478 == 32'h0000_0008 ? add_76503 : array_index_76497[8];
  assign array_update_76505[9] = add_76478 == 32'h0000_0009 ? add_76503 : array_index_76497[9];
  assign add_76506 = add_76493 + 32'h0000_0001;
  assign array_update_76507[0] = add_76070 == 32'h0000_0000 ? array_update_76505 : array_update_76494[0];
  assign array_update_76507[1] = add_76070 == 32'h0000_0001 ? array_update_76505 : array_update_76494[1];
  assign array_update_76507[2] = add_76070 == 32'h0000_0002 ? array_update_76505 : array_update_76494[2];
  assign array_update_76507[3] = add_76070 == 32'h0000_0003 ? array_update_76505 : array_update_76494[3];
  assign array_update_76507[4] = add_76070 == 32'h0000_0004 ? array_update_76505 : array_update_76494[4];
  assign array_update_76507[5] = add_76070 == 32'h0000_0005 ? array_update_76505 : array_update_76494[5];
  assign array_update_76507[6] = add_76070 == 32'h0000_0006 ? array_update_76505 : array_update_76494[6];
  assign array_update_76507[7] = add_76070 == 32'h0000_0007 ? array_update_76505 : array_update_76494[7];
  assign array_update_76507[8] = add_76070 == 32'h0000_0008 ? array_update_76505 : array_update_76494[8];
  assign array_update_76507[9] = add_76070 == 32'h0000_0009 ? array_update_76505 : array_update_76494[9];
  assign array_index_76509 = array_update_72021[add_76506 > 32'h0000_0009 ? 4'h9 : add_76506[3:0]];
  assign array_index_76510 = array_update_76507[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_76514 = smul32b_32b_x_32b(array_index_76077[add_76506 > 32'h0000_0009 ? 4'h9 : add_76506[3:0]], array_index_76509[add_76478 > 32'h0000_0009 ? 4'h9 : add_76478[3:0]]);
  assign add_76516 = array_index_76510[add_76478 > 32'h0000_0009 ? 4'h9 : add_76478[3:0]] + smul_76514;
  assign array_update_76518[0] = add_76478 == 32'h0000_0000 ? add_76516 : array_index_76510[0];
  assign array_update_76518[1] = add_76478 == 32'h0000_0001 ? add_76516 : array_index_76510[1];
  assign array_update_76518[2] = add_76478 == 32'h0000_0002 ? add_76516 : array_index_76510[2];
  assign array_update_76518[3] = add_76478 == 32'h0000_0003 ? add_76516 : array_index_76510[3];
  assign array_update_76518[4] = add_76478 == 32'h0000_0004 ? add_76516 : array_index_76510[4];
  assign array_update_76518[5] = add_76478 == 32'h0000_0005 ? add_76516 : array_index_76510[5];
  assign array_update_76518[6] = add_76478 == 32'h0000_0006 ? add_76516 : array_index_76510[6];
  assign array_update_76518[7] = add_76478 == 32'h0000_0007 ? add_76516 : array_index_76510[7];
  assign array_update_76518[8] = add_76478 == 32'h0000_0008 ? add_76516 : array_index_76510[8];
  assign array_update_76518[9] = add_76478 == 32'h0000_0009 ? add_76516 : array_index_76510[9];
  assign add_76519 = add_76506 + 32'h0000_0001;
  assign array_update_76520[0] = add_76070 == 32'h0000_0000 ? array_update_76518 : array_update_76507[0];
  assign array_update_76520[1] = add_76070 == 32'h0000_0001 ? array_update_76518 : array_update_76507[1];
  assign array_update_76520[2] = add_76070 == 32'h0000_0002 ? array_update_76518 : array_update_76507[2];
  assign array_update_76520[3] = add_76070 == 32'h0000_0003 ? array_update_76518 : array_update_76507[3];
  assign array_update_76520[4] = add_76070 == 32'h0000_0004 ? array_update_76518 : array_update_76507[4];
  assign array_update_76520[5] = add_76070 == 32'h0000_0005 ? array_update_76518 : array_update_76507[5];
  assign array_update_76520[6] = add_76070 == 32'h0000_0006 ? array_update_76518 : array_update_76507[6];
  assign array_update_76520[7] = add_76070 == 32'h0000_0007 ? array_update_76518 : array_update_76507[7];
  assign array_update_76520[8] = add_76070 == 32'h0000_0008 ? array_update_76518 : array_update_76507[8];
  assign array_update_76520[9] = add_76070 == 32'h0000_0009 ? array_update_76518 : array_update_76507[9];
  assign array_index_76522 = array_update_72021[add_76519 > 32'h0000_0009 ? 4'h9 : add_76519[3:0]];
  assign array_index_76523 = array_update_76520[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_76527 = smul32b_32b_x_32b(array_index_76077[add_76519 > 32'h0000_0009 ? 4'h9 : add_76519[3:0]], array_index_76522[add_76478 > 32'h0000_0009 ? 4'h9 : add_76478[3:0]]);
  assign add_76529 = array_index_76523[add_76478 > 32'h0000_0009 ? 4'h9 : add_76478[3:0]] + smul_76527;
  assign array_update_76531[0] = add_76478 == 32'h0000_0000 ? add_76529 : array_index_76523[0];
  assign array_update_76531[1] = add_76478 == 32'h0000_0001 ? add_76529 : array_index_76523[1];
  assign array_update_76531[2] = add_76478 == 32'h0000_0002 ? add_76529 : array_index_76523[2];
  assign array_update_76531[3] = add_76478 == 32'h0000_0003 ? add_76529 : array_index_76523[3];
  assign array_update_76531[4] = add_76478 == 32'h0000_0004 ? add_76529 : array_index_76523[4];
  assign array_update_76531[5] = add_76478 == 32'h0000_0005 ? add_76529 : array_index_76523[5];
  assign array_update_76531[6] = add_76478 == 32'h0000_0006 ? add_76529 : array_index_76523[6];
  assign array_update_76531[7] = add_76478 == 32'h0000_0007 ? add_76529 : array_index_76523[7];
  assign array_update_76531[8] = add_76478 == 32'h0000_0008 ? add_76529 : array_index_76523[8];
  assign array_update_76531[9] = add_76478 == 32'h0000_0009 ? add_76529 : array_index_76523[9];
  assign add_76532 = add_76519 + 32'h0000_0001;
  assign array_update_76533[0] = add_76070 == 32'h0000_0000 ? array_update_76531 : array_update_76520[0];
  assign array_update_76533[1] = add_76070 == 32'h0000_0001 ? array_update_76531 : array_update_76520[1];
  assign array_update_76533[2] = add_76070 == 32'h0000_0002 ? array_update_76531 : array_update_76520[2];
  assign array_update_76533[3] = add_76070 == 32'h0000_0003 ? array_update_76531 : array_update_76520[3];
  assign array_update_76533[4] = add_76070 == 32'h0000_0004 ? array_update_76531 : array_update_76520[4];
  assign array_update_76533[5] = add_76070 == 32'h0000_0005 ? array_update_76531 : array_update_76520[5];
  assign array_update_76533[6] = add_76070 == 32'h0000_0006 ? array_update_76531 : array_update_76520[6];
  assign array_update_76533[7] = add_76070 == 32'h0000_0007 ? array_update_76531 : array_update_76520[7];
  assign array_update_76533[8] = add_76070 == 32'h0000_0008 ? array_update_76531 : array_update_76520[8];
  assign array_update_76533[9] = add_76070 == 32'h0000_0009 ? array_update_76531 : array_update_76520[9];
  assign array_index_76535 = array_update_72021[add_76532 > 32'h0000_0009 ? 4'h9 : add_76532[3:0]];
  assign array_index_76536 = array_update_76533[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_76540 = smul32b_32b_x_32b(array_index_76077[add_76532 > 32'h0000_0009 ? 4'h9 : add_76532[3:0]], array_index_76535[add_76478 > 32'h0000_0009 ? 4'h9 : add_76478[3:0]]);
  assign add_76542 = array_index_76536[add_76478 > 32'h0000_0009 ? 4'h9 : add_76478[3:0]] + smul_76540;
  assign array_update_76544[0] = add_76478 == 32'h0000_0000 ? add_76542 : array_index_76536[0];
  assign array_update_76544[1] = add_76478 == 32'h0000_0001 ? add_76542 : array_index_76536[1];
  assign array_update_76544[2] = add_76478 == 32'h0000_0002 ? add_76542 : array_index_76536[2];
  assign array_update_76544[3] = add_76478 == 32'h0000_0003 ? add_76542 : array_index_76536[3];
  assign array_update_76544[4] = add_76478 == 32'h0000_0004 ? add_76542 : array_index_76536[4];
  assign array_update_76544[5] = add_76478 == 32'h0000_0005 ? add_76542 : array_index_76536[5];
  assign array_update_76544[6] = add_76478 == 32'h0000_0006 ? add_76542 : array_index_76536[6];
  assign array_update_76544[7] = add_76478 == 32'h0000_0007 ? add_76542 : array_index_76536[7];
  assign array_update_76544[8] = add_76478 == 32'h0000_0008 ? add_76542 : array_index_76536[8];
  assign array_update_76544[9] = add_76478 == 32'h0000_0009 ? add_76542 : array_index_76536[9];
  assign add_76545 = add_76532 + 32'h0000_0001;
  assign array_update_76546[0] = add_76070 == 32'h0000_0000 ? array_update_76544 : array_update_76533[0];
  assign array_update_76546[1] = add_76070 == 32'h0000_0001 ? array_update_76544 : array_update_76533[1];
  assign array_update_76546[2] = add_76070 == 32'h0000_0002 ? array_update_76544 : array_update_76533[2];
  assign array_update_76546[3] = add_76070 == 32'h0000_0003 ? array_update_76544 : array_update_76533[3];
  assign array_update_76546[4] = add_76070 == 32'h0000_0004 ? array_update_76544 : array_update_76533[4];
  assign array_update_76546[5] = add_76070 == 32'h0000_0005 ? array_update_76544 : array_update_76533[5];
  assign array_update_76546[6] = add_76070 == 32'h0000_0006 ? array_update_76544 : array_update_76533[6];
  assign array_update_76546[7] = add_76070 == 32'h0000_0007 ? array_update_76544 : array_update_76533[7];
  assign array_update_76546[8] = add_76070 == 32'h0000_0008 ? array_update_76544 : array_update_76533[8];
  assign array_update_76546[9] = add_76070 == 32'h0000_0009 ? array_update_76544 : array_update_76533[9];
  assign array_index_76548 = array_update_72021[add_76545 > 32'h0000_0009 ? 4'h9 : add_76545[3:0]];
  assign array_index_76549 = array_update_76546[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_76553 = smul32b_32b_x_32b(array_index_76077[add_76545 > 32'h0000_0009 ? 4'h9 : add_76545[3:0]], array_index_76548[add_76478 > 32'h0000_0009 ? 4'h9 : add_76478[3:0]]);
  assign add_76555 = array_index_76549[add_76478 > 32'h0000_0009 ? 4'h9 : add_76478[3:0]] + smul_76553;
  assign array_update_76557[0] = add_76478 == 32'h0000_0000 ? add_76555 : array_index_76549[0];
  assign array_update_76557[1] = add_76478 == 32'h0000_0001 ? add_76555 : array_index_76549[1];
  assign array_update_76557[2] = add_76478 == 32'h0000_0002 ? add_76555 : array_index_76549[2];
  assign array_update_76557[3] = add_76478 == 32'h0000_0003 ? add_76555 : array_index_76549[3];
  assign array_update_76557[4] = add_76478 == 32'h0000_0004 ? add_76555 : array_index_76549[4];
  assign array_update_76557[5] = add_76478 == 32'h0000_0005 ? add_76555 : array_index_76549[5];
  assign array_update_76557[6] = add_76478 == 32'h0000_0006 ? add_76555 : array_index_76549[6];
  assign array_update_76557[7] = add_76478 == 32'h0000_0007 ? add_76555 : array_index_76549[7];
  assign array_update_76557[8] = add_76478 == 32'h0000_0008 ? add_76555 : array_index_76549[8];
  assign array_update_76557[9] = add_76478 == 32'h0000_0009 ? add_76555 : array_index_76549[9];
  assign add_76558 = add_76545 + 32'h0000_0001;
  assign array_update_76559[0] = add_76070 == 32'h0000_0000 ? array_update_76557 : array_update_76546[0];
  assign array_update_76559[1] = add_76070 == 32'h0000_0001 ? array_update_76557 : array_update_76546[1];
  assign array_update_76559[2] = add_76070 == 32'h0000_0002 ? array_update_76557 : array_update_76546[2];
  assign array_update_76559[3] = add_76070 == 32'h0000_0003 ? array_update_76557 : array_update_76546[3];
  assign array_update_76559[4] = add_76070 == 32'h0000_0004 ? array_update_76557 : array_update_76546[4];
  assign array_update_76559[5] = add_76070 == 32'h0000_0005 ? array_update_76557 : array_update_76546[5];
  assign array_update_76559[6] = add_76070 == 32'h0000_0006 ? array_update_76557 : array_update_76546[6];
  assign array_update_76559[7] = add_76070 == 32'h0000_0007 ? array_update_76557 : array_update_76546[7];
  assign array_update_76559[8] = add_76070 == 32'h0000_0008 ? array_update_76557 : array_update_76546[8];
  assign array_update_76559[9] = add_76070 == 32'h0000_0009 ? array_update_76557 : array_update_76546[9];
  assign array_index_76561 = array_update_72021[add_76558 > 32'h0000_0009 ? 4'h9 : add_76558[3:0]];
  assign array_index_76562 = array_update_76559[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_76566 = smul32b_32b_x_32b(array_index_76077[add_76558 > 32'h0000_0009 ? 4'h9 : add_76558[3:0]], array_index_76561[add_76478 > 32'h0000_0009 ? 4'h9 : add_76478[3:0]]);
  assign add_76568 = array_index_76562[add_76478 > 32'h0000_0009 ? 4'h9 : add_76478[3:0]] + smul_76566;
  assign array_update_76570[0] = add_76478 == 32'h0000_0000 ? add_76568 : array_index_76562[0];
  assign array_update_76570[1] = add_76478 == 32'h0000_0001 ? add_76568 : array_index_76562[1];
  assign array_update_76570[2] = add_76478 == 32'h0000_0002 ? add_76568 : array_index_76562[2];
  assign array_update_76570[3] = add_76478 == 32'h0000_0003 ? add_76568 : array_index_76562[3];
  assign array_update_76570[4] = add_76478 == 32'h0000_0004 ? add_76568 : array_index_76562[4];
  assign array_update_76570[5] = add_76478 == 32'h0000_0005 ? add_76568 : array_index_76562[5];
  assign array_update_76570[6] = add_76478 == 32'h0000_0006 ? add_76568 : array_index_76562[6];
  assign array_update_76570[7] = add_76478 == 32'h0000_0007 ? add_76568 : array_index_76562[7];
  assign array_update_76570[8] = add_76478 == 32'h0000_0008 ? add_76568 : array_index_76562[8];
  assign array_update_76570[9] = add_76478 == 32'h0000_0009 ? add_76568 : array_index_76562[9];
  assign add_76571 = add_76558 + 32'h0000_0001;
  assign array_update_76572[0] = add_76070 == 32'h0000_0000 ? array_update_76570 : array_update_76559[0];
  assign array_update_76572[1] = add_76070 == 32'h0000_0001 ? array_update_76570 : array_update_76559[1];
  assign array_update_76572[2] = add_76070 == 32'h0000_0002 ? array_update_76570 : array_update_76559[2];
  assign array_update_76572[3] = add_76070 == 32'h0000_0003 ? array_update_76570 : array_update_76559[3];
  assign array_update_76572[4] = add_76070 == 32'h0000_0004 ? array_update_76570 : array_update_76559[4];
  assign array_update_76572[5] = add_76070 == 32'h0000_0005 ? array_update_76570 : array_update_76559[5];
  assign array_update_76572[6] = add_76070 == 32'h0000_0006 ? array_update_76570 : array_update_76559[6];
  assign array_update_76572[7] = add_76070 == 32'h0000_0007 ? array_update_76570 : array_update_76559[7];
  assign array_update_76572[8] = add_76070 == 32'h0000_0008 ? array_update_76570 : array_update_76559[8];
  assign array_update_76572[9] = add_76070 == 32'h0000_0009 ? array_update_76570 : array_update_76559[9];
  assign array_index_76574 = array_update_72021[add_76571 > 32'h0000_0009 ? 4'h9 : add_76571[3:0]];
  assign array_index_76575 = array_update_76572[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_76579 = smul32b_32b_x_32b(array_index_76077[add_76571 > 32'h0000_0009 ? 4'h9 : add_76571[3:0]], array_index_76574[add_76478 > 32'h0000_0009 ? 4'h9 : add_76478[3:0]]);
  assign add_76581 = array_index_76575[add_76478 > 32'h0000_0009 ? 4'h9 : add_76478[3:0]] + smul_76579;
  assign array_update_76583[0] = add_76478 == 32'h0000_0000 ? add_76581 : array_index_76575[0];
  assign array_update_76583[1] = add_76478 == 32'h0000_0001 ? add_76581 : array_index_76575[1];
  assign array_update_76583[2] = add_76478 == 32'h0000_0002 ? add_76581 : array_index_76575[2];
  assign array_update_76583[3] = add_76478 == 32'h0000_0003 ? add_76581 : array_index_76575[3];
  assign array_update_76583[4] = add_76478 == 32'h0000_0004 ? add_76581 : array_index_76575[4];
  assign array_update_76583[5] = add_76478 == 32'h0000_0005 ? add_76581 : array_index_76575[5];
  assign array_update_76583[6] = add_76478 == 32'h0000_0006 ? add_76581 : array_index_76575[6];
  assign array_update_76583[7] = add_76478 == 32'h0000_0007 ? add_76581 : array_index_76575[7];
  assign array_update_76583[8] = add_76478 == 32'h0000_0008 ? add_76581 : array_index_76575[8];
  assign array_update_76583[9] = add_76478 == 32'h0000_0009 ? add_76581 : array_index_76575[9];
  assign add_76584 = add_76571 + 32'h0000_0001;
  assign array_update_76585[0] = add_76070 == 32'h0000_0000 ? array_update_76583 : array_update_76572[0];
  assign array_update_76585[1] = add_76070 == 32'h0000_0001 ? array_update_76583 : array_update_76572[1];
  assign array_update_76585[2] = add_76070 == 32'h0000_0002 ? array_update_76583 : array_update_76572[2];
  assign array_update_76585[3] = add_76070 == 32'h0000_0003 ? array_update_76583 : array_update_76572[3];
  assign array_update_76585[4] = add_76070 == 32'h0000_0004 ? array_update_76583 : array_update_76572[4];
  assign array_update_76585[5] = add_76070 == 32'h0000_0005 ? array_update_76583 : array_update_76572[5];
  assign array_update_76585[6] = add_76070 == 32'h0000_0006 ? array_update_76583 : array_update_76572[6];
  assign array_update_76585[7] = add_76070 == 32'h0000_0007 ? array_update_76583 : array_update_76572[7];
  assign array_update_76585[8] = add_76070 == 32'h0000_0008 ? array_update_76583 : array_update_76572[8];
  assign array_update_76585[9] = add_76070 == 32'h0000_0009 ? array_update_76583 : array_update_76572[9];
  assign array_index_76587 = array_update_72021[add_76584 > 32'h0000_0009 ? 4'h9 : add_76584[3:0]];
  assign array_index_76588 = array_update_76585[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_76592 = smul32b_32b_x_32b(array_index_76077[add_76584 > 32'h0000_0009 ? 4'h9 : add_76584[3:0]], array_index_76587[add_76478 > 32'h0000_0009 ? 4'h9 : add_76478[3:0]]);
  assign add_76594 = array_index_76588[add_76478 > 32'h0000_0009 ? 4'h9 : add_76478[3:0]] + smul_76592;
  assign array_update_76596[0] = add_76478 == 32'h0000_0000 ? add_76594 : array_index_76588[0];
  assign array_update_76596[1] = add_76478 == 32'h0000_0001 ? add_76594 : array_index_76588[1];
  assign array_update_76596[2] = add_76478 == 32'h0000_0002 ? add_76594 : array_index_76588[2];
  assign array_update_76596[3] = add_76478 == 32'h0000_0003 ? add_76594 : array_index_76588[3];
  assign array_update_76596[4] = add_76478 == 32'h0000_0004 ? add_76594 : array_index_76588[4];
  assign array_update_76596[5] = add_76478 == 32'h0000_0005 ? add_76594 : array_index_76588[5];
  assign array_update_76596[6] = add_76478 == 32'h0000_0006 ? add_76594 : array_index_76588[6];
  assign array_update_76596[7] = add_76478 == 32'h0000_0007 ? add_76594 : array_index_76588[7];
  assign array_update_76596[8] = add_76478 == 32'h0000_0008 ? add_76594 : array_index_76588[8];
  assign array_update_76596[9] = add_76478 == 32'h0000_0009 ? add_76594 : array_index_76588[9];
  assign add_76597 = add_76584 + 32'h0000_0001;
  assign array_update_76598[0] = add_76070 == 32'h0000_0000 ? array_update_76596 : array_update_76585[0];
  assign array_update_76598[1] = add_76070 == 32'h0000_0001 ? array_update_76596 : array_update_76585[1];
  assign array_update_76598[2] = add_76070 == 32'h0000_0002 ? array_update_76596 : array_update_76585[2];
  assign array_update_76598[3] = add_76070 == 32'h0000_0003 ? array_update_76596 : array_update_76585[3];
  assign array_update_76598[4] = add_76070 == 32'h0000_0004 ? array_update_76596 : array_update_76585[4];
  assign array_update_76598[5] = add_76070 == 32'h0000_0005 ? array_update_76596 : array_update_76585[5];
  assign array_update_76598[6] = add_76070 == 32'h0000_0006 ? array_update_76596 : array_update_76585[6];
  assign array_update_76598[7] = add_76070 == 32'h0000_0007 ? array_update_76596 : array_update_76585[7];
  assign array_update_76598[8] = add_76070 == 32'h0000_0008 ? array_update_76596 : array_update_76585[8];
  assign array_update_76598[9] = add_76070 == 32'h0000_0009 ? array_update_76596 : array_update_76585[9];
  assign array_index_76600 = array_update_72021[add_76597 > 32'h0000_0009 ? 4'h9 : add_76597[3:0]];
  assign array_index_76601 = array_update_76598[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_76605 = smul32b_32b_x_32b(array_index_76077[add_76597 > 32'h0000_0009 ? 4'h9 : add_76597[3:0]], array_index_76600[add_76478 > 32'h0000_0009 ? 4'h9 : add_76478[3:0]]);
  assign add_76607 = array_index_76601[add_76478 > 32'h0000_0009 ? 4'h9 : add_76478[3:0]] + smul_76605;
  assign array_update_76608[0] = add_76478 == 32'h0000_0000 ? add_76607 : array_index_76601[0];
  assign array_update_76608[1] = add_76478 == 32'h0000_0001 ? add_76607 : array_index_76601[1];
  assign array_update_76608[2] = add_76478 == 32'h0000_0002 ? add_76607 : array_index_76601[2];
  assign array_update_76608[3] = add_76478 == 32'h0000_0003 ? add_76607 : array_index_76601[3];
  assign array_update_76608[4] = add_76478 == 32'h0000_0004 ? add_76607 : array_index_76601[4];
  assign array_update_76608[5] = add_76478 == 32'h0000_0005 ? add_76607 : array_index_76601[5];
  assign array_update_76608[6] = add_76478 == 32'h0000_0006 ? add_76607 : array_index_76601[6];
  assign array_update_76608[7] = add_76478 == 32'h0000_0007 ? add_76607 : array_index_76601[7];
  assign array_update_76608[8] = add_76478 == 32'h0000_0008 ? add_76607 : array_index_76601[8];
  assign array_update_76608[9] = add_76478 == 32'h0000_0009 ? add_76607 : array_index_76601[9];
  assign array_update_76609[0] = add_76070 == 32'h0000_0000 ? array_update_76608 : array_update_76598[0];
  assign array_update_76609[1] = add_76070 == 32'h0000_0001 ? array_update_76608 : array_update_76598[1];
  assign array_update_76609[2] = add_76070 == 32'h0000_0002 ? array_update_76608 : array_update_76598[2];
  assign array_update_76609[3] = add_76070 == 32'h0000_0003 ? array_update_76608 : array_update_76598[3];
  assign array_update_76609[4] = add_76070 == 32'h0000_0004 ? array_update_76608 : array_update_76598[4];
  assign array_update_76609[5] = add_76070 == 32'h0000_0005 ? array_update_76608 : array_update_76598[5];
  assign array_update_76609[6] = add_76070 == 32'h0000_0006 ? array_update_76608 : array_update_76598[6];
  assign array_update_76609[7] = add_76070 == 32'h0000_0007 ? array_update_76608 : array_update_76598[7];
  assign array_update_76609[8] = add_76070 == 32'h0000_0008 ? array_update_76608 : array_update_76598[8];
  assign array_update_76609[9] = add_76070 == 32'h0000_0009 ? array_update_76608 : array_update_76598[9];
  assign array_index_76611 = array_update_76609[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign add_76613 = add_76478 + 32'h0000_0001;
  assign array_update_76614[0] = add_76613 == 32'h0000_0000 ? 32'h0000_0000 : array_index_76611[0];
  assign array_update_76614[1] = add_76613 == 32'h0000_0001 ? 32'h0000_0000 : array_index_76611[1];
  assign array_update_76614[2] = add_76613 == 32'h0000_0002 ? 32'h0000_0000 : array_index_76611[2];
  assign array_update_76614[3] = add_76613 == 32'h0000_0003 ? 32'h0000_0000 : array_index_76611[3];
  assign array_update_76614[4] = add_76613 == 32'h0000_0004 ? 32'h0000_0000 : array_index_76611[4];
  assign array_update_76614[5] = add_76613 == 32'h0000_0005 ? 32'h0000_0000 : array_index_76611[5];
  assign array_update_76614[6] = add_76613 == 32'h0000_0006 ? 32'h0000_0000 : array_index_76611[6];
  assign array_update_76614[7] = add_76613 == 32'h0000_0007 ? 32'h0000_0000 : array_index_76611[7];
  assign array_update_76614[8] = add_76613 == 32'h0000_0008 ? 32'h0000_0000 : array_index_76611[8];
  assign array_update_76614[9] = add_76613 == 32'h0000_0009 ? 32'h0000_0000 : array_index_76611[9];
  assign literal_76615 = 32'h0000_0000;
  assign array_update_76616[0] = add_76070 == 32'h0000_0000 ? array_update_76614 : array_update_76609[0];
  assign array_update_76616[1] = add_76070 == 32'h0000_0001 ? array_update_76614 : array_update_76609[1];
  assign array_update_76616[2] = add_76070 == 32'h0000_0002 ? array_update_76614 : array_update_76609[2];
  assign array_update_76616[3] = add_76070 == 32'h0000_0003 ? array_update_76614 : array_update_76609[3];
  assign array_update_76616[4] = add_76070 == 32'h0000_0004 ? array_update_76614 : array_update_76609[4];
  assign array_update_76616[5] = add_76070 == 32'h0000_0005 ? array_update_76614 : array_update_76609[5];
  assign array_update_76616[6] = add_76070 == 32'h0000_0006 ? array_update_76614 : array_update_76609[6];
  assign array_update_76616[7] = add_76070 == 32'h0000_0007 ? array_update_76614 : array_update_76609[7];
  assign array_update_76616[8] = add_76070 == 32'h0000_0008 ? array_update_76614 : array_update_76609[8];
  assign array_update_76616[9] = add_76070 == 32'h0000_0009 ? array_update_76614 : array_update_76609[9];
  assign array_index_76618 = array_update_72021[literal_76615 > 32'h0000_0009 ? 4'h9 : literal_76615[3:0]];
  assign array_index_76619 = array_update_76616[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_76623 = smul32b_32b_x_32b(array_index_76077[literal_76615 > 32'h0000_0009 ? 4'h9 : literal_76615[3:0]], array_index_76618[add_76613 > 32'h0000_0009 ? 4'h9 : add_76613[3:0]]);
  assign add_76625 = array_index_76619[add_76613 > 32'h0000_0009 ? 4'h9 : add_76613[3:0]] + smul_76623;
  assign array_update_76627[0] = add_76613 == 32'h0000_0000 ? add_76625 : array_index_76619[0];
  assign array_update_76627[1] = add_76613 == 32'h0000_0001 ? add_76625 : array_index_76619[1];
  assign array_update_76627[2] = add_76613 == 32'h0000_0002 ? add_76625 : array_index_76619[2];
  assign array_update_76627[3] = add_76613 == 32'h0000_0003 ? add_76625 : array_index_76619[3];
  assign array_update_76627[4] = add_76613 == 32'h0000_0004 ? add_76625 : array_index_76619[4];
  assign array_update_76627[5] = add_76613 == 32'h0000_0005 ? add_76625 : array_index_76619[5];
  assign array_update_76627[6] = add_76613 == 32'h0000_0006 ? add_76625 : array_index_76619[6];
  assign array_update_76627[7] = add_76613 == 32'h0000_0007 ? add_76625 : array_index_76619[7];
  assign array_update_76627[8] = add_76613 == 32'h0000_0008 ? add_76625 : array_index_76619[8];
  assign array_update_76627[9] = add_76613 == 32'h0000_0009 ? add_76625 : array_index_76619[9];
  assign add_76628 = literal_76615 + 32'h0000_0001;
  assign array_update_76629[0] = add_76070 == 32'h0000_0000 ? array_update_76627 : array_update_76616[0];
  assign array_update_76629[1] = add_76070 == 32'h0000_0001 ? array_update_76627 : array_update_76616[1];
  assign array_update_76629[2] = add_76070 == 32'h0000_0002 ? array_update_76627 : array_update_76616[2];
  assign array_update_76629[3] = add_76070 == 32'h0000_0003 ? array_update_76627 : array_update_76616[3];
  assign array_update_76629[4] = add_76070 == 32'h0000_0004 ? array_update_76627 : array_update_76616[4];
  assign array_update_76629[5] = add_76070 == 32'h0000_0005 ? array_update_76627 : array_update_76616[5];
  assign array_update_76629[6] = add_76070 == 32'h0000_0006 ? array_update_76627 : array_update_76616[6];
  assign array_update_76629[7] = add_76070 == 32'h0000_0007 ? array_update_76627 : array_update_76616[7];
  assign array_update_76629[8] = add_76070 == 32'h0000_0008 ? array_update_76627 : array_update_76616[8];
  assign array_update_76629[9] = add_76070 == 32'h0000_0009 ? array_update_76627 : array_update_76616[9];
  assign array_index_76631 = array_update_72021[add_76628 > 32'h0000_0009 ? 4'h9 : add_76628[3:0]];
  assign array_index_76632 = array_update_76629[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_76636 = smul32b_32b_x_32b(array_index_76077[add_76628 > 32'h0000_0009 ? 4'h9 : add_76628[3:0]], array_index_76631[add_76613 > 32'h0000_0009 ? 4'h9 : add_76613[3:0]]);
  assign add_76638 = array_index_76632[add_76613 > 32'h0000_0009 ? 4'h9 : add_76613[3:0]] + smul_76636;
  assign array_update_76640[0] = add_76613 == 32'h0000_0000 ? add_76638 : array_index_76632[0];
  assign array_update_76640[1] = add_76613 == 32'h0000_0001 ? add_76638 : array_index_76632[1];
  assign array_update_76640[2] = add_76613 == 32'h0000_0002 ? add_76638 : array_index_76632[2];
  assign array_update_76640[3] = add_76613 == 32'h0000_0003 ? add_76638 : array_index_76632[3];
  assign array_update_76640[4] = add_76613 == 32'h0000_0004 ? add_76638 : array_index_76632[4];
  assign array_update_76640[5] = add_76613 == 32'h0000_0005 ? add_76638 : array_index_76632[5];
  assign array_update_76640[6] = add_76613 == 32'h0000_0006 ? add_76638 : array_index_76632[6];
  assign array_update_76640[7] = add_76613 == 32'h0000_0007 ? add_76638 : array_index_76632[7];
  assign array_update_76640[8] = add_76613 == 32'h0000_0008 ? add_76638 : array_index_76632[8];
  assign array_update_76640[9] = add_76613 == 32'h0000_0009 ? add_76638 : array_index_76632[9];
  assign add_76641 = add_76628 + 32'h0000_0001;
  assign array_update_76642[0] = add_76070 == 32'h0000_0000 ? array_update_76640 : array_update_76629[0];
  assign array_update_76642[1] = add_76070 == 32'h0000_0001 ? array_update_76640 : array_update_76629[1];
  assign array_update_76642[2] = add_76070 == 32'h0000_0002 ? array_update_76640 : array_update_76629[2];
  assign array_update_76642[3] = add_76070 == 32'h0000_0003 ? array_update_76640 : array_update_76629[3];
  assign array_update_76642[4] = add_76070 == 32'h0000_0004 ? array_update_76640 : array_update_76629[4];
  assign array_update_76642[5] = add_76070 == 32'h0000_0005 ? array_update_76640 : array_update_76629[5];
  assign array_update_76642[6] = add_76070 == 32'h0000_0006 ? array_update_76640 : array_update_76629[6];
  assign array_update_76642[7] = add_76070 == 32'h0000_0007 ? array_update_76640 : array_update_76629[7];
  assign array_update_76642[8] = add_76070 == 32'h0000_0008 ? array_update_76640 : array_update_76629[8];
  assign array_update_76642[9] = add_76070 == 32'h0000_0009 ? array_update_76640 : array_update_76629[9];
  assign array_index_76644 = array_update_72021[add_76641 > 32'h0000_0009 ? 4'h9 : add_76641[3:0]];
  assign array_index_76645 = array_update_76642[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_76649 = smul32b_32b_x_32b(array_index_76077[add_76641 > 32'h0000_0009 ? 4'h9 : add_76641[3:0]], array_index_76644[add_76613 > 32'h0000_0009 ? 4'h9 : add_76613[3:0]]);
  assign add_76651 = array_index_76645[add_76613 > 32'h0000_0009 ? 4'h9 : add_76613[3:0]] + smul_76649;
  assign array_update_76653[0] = add_76613 == 32'h0000_0000 ? add_76651 : array_index_76645[0];
  assign array_update_76653[1] = add_76613 == 32'h0000_0001 ? add_76651 : array_index_76645[1];
  assign array_update_76653[2] = add_76613 == 32'h0000_0002 ? add_76651 : array_index_76645[2];
  assign array_update_76653[3] = add_76613 == 32'h0000_0003 ? add_76651 : array_index_76645[3];
  assign array_update_76653[4] = add_76613 == 32'h0000_0004 ? add_76651 : array_index_76645[4];
  assign array_update_76653[5] = add_76613 == 32'h0000_0005 ? add_76651 : array_index_76645[5];
  assign array_update_76653[6] = add_76613 == 32'h0000_0006 ? add_76651 : array_index_76645[6];
  assign array_update_76653[7] = add_76613 == 32'h0000_0007 ? add_76651 : array_index_76645[7];
  assign array_update_76653[8] = add_76613 == 32'h0000_0008 ? add_76651 : array_index_76645[8];
  assign array_update_76653[9] = add_76613 == 32'h0000_0009 ? add_76651 : array_index_76645[9];
  assign add_76654 = add_76641 + 32'h0000_0001;
  assign array_update_76655[0] = add_76070 == 32'h0000_0000 ? array_update_76653 : array_update_76642[0];
  assign array_update_76655[1] = add_76070 == 32'h0000_0001 ? array_update_76653 : array_update_76642[1];
  assign array_update_76655[2] = add_76070 == 32'h0000_0002 ? array_update_76653 : array_update_76642[2];
  assign array_update_76655[3] = add_76070 == 32'h0000_0003 ? array_update_76653 : array_update_76642[3];
  assign array_update_76655[4] = add_76070 == 32'h0000_0004 ? array_update_76653 : array_update_76642[4];
  assign array_update_76655[5] = add_76070 == 32'h0000_0005 ? array_update_76653 : array_update_76642[5];
  assign array_update_76655[6] = add_76070 == 32'h0000_0006 ? array_update_76653 : array_update_76642[6];
  assign array_update_76655[7] = add_76070 == 32'h0000_0007 ? array_update_76653 : array_update_76642[7];
  assign array_update_76655[8] = add_76070 == 32'h0000_0008 ? array_update_76653 : array_update_76642[8];
  assign array_update_76655[9] = add_76070 == 32'h0000_0009 ? array_update_76653 : array_update_76642[9];
  assign array_index_76657 = array_update_72021[add_76654 > 32'h0000_0009 ? 4'h9 : add_76654[3:0]];
  assign array_index_76658 = array_update_76655[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_76662 = smul32b_32b_x_32b(array_index_76077[add_76654 > 32'h0000_0009 ? 4'h9 : add_76654[3:0]], array_index_76657[add_76613 > 32'h0000_0009 ? 4'h9 : add_76613[3:0]]);
  assign add_76664 = array_index_76658[add_76613 > 32'h0000_0009 ? 4'h9 : add_76613[3:0]] + smul_76662;
  assign array_update_76666[0] = add_76613 == 32'h0000_0000 ? add_76664 : array_index_76658[0];
  assign array_update_76666[1] = add_76613 == 32'h0000_0001 ? add_76664 : array_index_76658[1];
  assign array_update_76666[2] = add_76613 == 32'h0000_0002 ? add_76664 : array_index_76658[2];
  assign array_update_76666[3] = add_76613 == 32'h0000_0003 ? add_76664 : array_index_76658[3];
  assign array_update_76666[4] = add_76613 == 32'h0000_0004 ? add_76664 : array_index_76658[4];
  assign array_update_76666[5] = add_76613 == 32'h0000_0005 ? add_76664 : array_index_76658[5];
  assign array_update_76666[6] = add_76613 == 32'h0000_0006 ? add_76664 : array_index_76658[6];
  assign array_update_76666[7] = add_76613 == 32'h0000_0007 ? add_76664 : array_index_76658[7];
  assign array_update_76666[8] = add_76613 == 32'h0000_0008 ? add_76664 : array_index_76658[8];
  assign array_update_76666[9] = add_76613 == 32'h0000_0009 ? add_76664 : array_index_76658[9];
  assign add_76667 = add_76654 + 32'h0000_0001;
  assign array_update_76668[0] = add_76070 == 32'h0000_0000 ? array_update_76666 : array_update_76655[0];
  assign array_update_76668[1] = add_76070 == 32'h0000_0001 ? array_update_76666 : array_update_76655[1];
  assign array_update_76668[2] = add_76070 == 32'h0000_0002 ? array_update_76666 : array_update_76655[2];
  assign array_update_76668[3] = add_76070 == 32'h0000_0003 ? array_update_76666 : array_update_76655[3];
  assign array_update_76668[4] = add_76070 == 32'h0000_0004 ? array_update_76666 : array_update_76655[4];
  assign array_update_76668[5] = add_76070 == 32'h0000_0005 ? array_update_76666 : array_update_76655[5];
  assign array_update_76668[6] = add_76070 == 32'h0000_0006 ? array_update_76666 : array_update_76655[6];
  assign array_update_76668[7] = add_76070 == 32'h0000_0007 ? array_update_76666 : array_update_76655[7];
  assign array_update_76668[8] = add_76070 == 32'h0000_0008 ? array_update_76666 : array_update_76655[8];
  assign array_update_76668[9] = add_76070 == 32'h0000_0009 ? array_update_76666 : array_update_76655[9];
  assign array_index_76670 = array_update_72021[add_76667 > 32'h0000_0009 ? 4'h9 : add_76667[3:0]];
  assign array_index_76671 = array_update_76668[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_76675 = smul32b_32b_x_32b(array_index_76077[add_76667 > 32'h0000_0009 ? 4'h9 : add_76667[3:0]], array_index_76670[add_76613 > 32'h0000_0009 ? 4'h9 : add_76613[3:0]]);
  assign add_76677 = array_index_76671[add_76613 > 32'h0000_0009 ? 4'h9 : add_76613[3:0]] + smul_76675;
  assign array_update_76679[0] = add_76613 == 32'h0000_0000 ? add_76677 : array_index_76671[0];
  assign array_update_76679[1] = add_76613 == 32'h0000_0001 ? add_76677 : array_index_76671[1];
  assign array_update_76679[2] = add_76613 == 32'h0000_0002 ? add_76677 : array_index_76671[2];
  assign array_update_76679[3] = add_76613 == 32'h0000_0003 ? add_76677 : array_index_76671[3];
  assign array_update_76679[4] = add_76613 == 32'h0000_0004 ? add_76677 : array_index_76671[4];
  assign array_update_76679[5] = add_76613 == 32'h0000_0005 ? add_76677 : array_index_76671[5];
  assign array_update_76679[6] = add_76613 == 32'h0000_0006 ? add_76677 : array_index_76671[6];
  assign array_update_76679[7] = add_76613 == 32'h0000_0007 ? add_76677 : array_index_76671[7];
  assign array_update_76679[8] = add_76613 == 32'h0000_0008 ? add_76677 : array_index_76671[8];
  assign array_update_76679[9] = add_76613 == 32'h0000_0009 ? add_76677 : array_index_76671[9];
  assign add_76680 = add_76667 + 32'h0000_0001;
  assign array_update_76681[0] = add_76070 == 32'h0000_0000 ? array_update_76679 : array_update_76668[0];
  assign array_update_76681[1] = add_76070 == 32'h0000_0001 ? array_update_76679 : array_update_76668[1];
  assign array_update_76681[2] = add_76070 == 32'h0000_0002 ? array_update_76679 : array_update_76668[2];
  assign array_update_76681[3] = add_76070 == 32'h0000_0003 ? array_update_76679 : array_update_76668[3];
  assign array_update_76681[4] = add_76070 == 32'h0000_0004 ? array_update_76679 : array_update_76668[4];
  assign array_update_76681[5] = add_76070 == 32'h0000_0005 ? array_update_76679 : array_update_76668[5];
  assign array_update_76681[6] = add_76070 == 32'h0000_0006 ? array_update_76679 : array_update_76668[6];
  assign array_update_76681[7] = add_76070 == 32'h0000_0007 ? array_update_76679 : array_update_76668[7];
  assign array_update_76681[8] = add_76070 == 32'h0000_0008 ? array_update_76679 : array_update_76668[8];
  assign array_update_76681[9] = add_76070 == 32'h0000_0009 ? array_update_76679 : array_update_76668[9];
  assign array_index_76683 = array_update_72021[add_76680 > 32'h0000_0009 ? 4'h9 : add_76680[3:0]];
  assign array_index_76684 = array_update_76681[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_76688 = smul32b_32b_x_32b(array_index_76077[add_76680 > 32'h0000_0009 ? 4'h9 : add_76680[3:0]], array_index_76683[add_76613 > 32'h0000_0009 ? 4'h9 : add_76613[3:0]]);
  assign add_76690 = array_index_76684[add_76613 > 32'h0000_0009 ? 4'h9 : add_76613[3:0]] + smul_76688;
  assign array_update_76692[0] = add_76613 == 32'h0000_0000 ? add_76690 : array_index_76684[0];
  assign array_update_76692[1] = add_76613 == 32'h0000_0001 ? add_76690 : array_index_76684[1];
  assign array_update_76692[2] = add_76613 == 32'h0000_0002 ? add_76690 : array_index_76684[2];
  assign array_update_76692[3] = add_76613 == 32'h0000_0003 ? add_76690 : array_index_76684[3];
  assign array_update_76692[4] = add_76613 == 32'h0000_0004 ? add_76690 : array_index_76684[4];
  assign array_update_76692[5] = add_76613 == 32'h0000_0005 ? add_76690 : array_index_76684[5];
  assign array_update_76692[6] = add_76613 == 32'h0000_0006 ? add_76690 : array_index_76684[6];
  assign array_update_76692[7] = add_76613 == 32'h0000_0007 ? add_76690 : array_index_76684[7];
  assign array_update_76692[8] = add_76613 == 32'h0000_0008 ? add_76690 : array_index_76684[8];
  assign array_update_76692[9] = add_76613 == 32'h0000_0009 ? add_76690 : array_index_76684[9];
  assign add_76693 = add_76680 + 32'h0000_0001;
  assign array_update_76694[0] = add_76070 == 32'h0000_0000 ? array_update_76692 : array_update_76681[0];
  assign array_update_76694[1] = add_76070 == 32'h0000_0001 ? array_update_76692 : array_update_76681[1];
  assign array_update_76694[2] = add_76070 == 32'h0000_0002 ? array_update_76692 : array_update_76681[2];
  assign array_update_76694[3] = add_76070 == 32'h0000_0003 ? array_update_76692 : array_update_76681[3];
  assign array_update_76694[4] = add_76070 == 32'h0000_0004 ? array_update_76692 : array_update_76681[4];
  assign array_update_76694[5] = add_76070 == 32'h0000_0005 ? array_update_76692 : array_update_76681[5];
  assign array_update_76694[6] = add_76070 == 32'h0000_0006 ? array_update_76692 : array_update_76681[6];
  assign array_update_76694[7] = add_76070 == 32'h0000_0007 ? array_update_76692 : array_update_76681[7];
  assign array_update_76694[8] = add_76070 == 32'h0000_0008 ? array_update_76692 : array_update_76681[8];
  assign array_update_76694[9] = add_76070 == 32'h0000_0009 ? array_update_76692 : array_update_76681[9];
  assign array_index_76696 = array_update_72021[add_76693 > 32'h0000_0009 ? 4'h9 : add_76693[3:0]];
  assign array_index_76697 = array_update_76694[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_76701 = smul32b_32b_x_32b(array_index_76077[add_76693 > 32'h0000_0009 ? 4'h9 : add_76693[3:0]], array_index_76696[add_76613 > 32'h0000_0009 ? 4'h9 : add_76613[3:0]]);
  assign add_76703 = array_index_76697[add_76613 > 32'h0000_0009 ? 4'h9 : add_76613[3:0]] + smul_76701;
  assign array_update_76705[0] = add_76613 == 32'h0000_0000 ? add_76703 : array_index_76697[0];
  assign array_update_76705[1] = add_76613 == 32'h0000_0001 ? add_76703 : array_index_76697[1];
  assign array_update_76705[2] = add_76613 == 32'h0000_0002 ? add_76703 : array_index_76697[2];
  assign array_update_76705[3] = add_76613 == 32'h0000_0003 ? add_76703 : array_index_76697[3];
  assign array_update_76705[4] = add_76613 == 32'h0000_0004 ? add_76703 : array_index_76697[4];
  assign array_update_76705[5] = add_76613 == 32'h0000_0005 ? add_76703 : array_index_76697[5];
  assign array_update_76705[6] = add_76613 == 32'h0000_0006 ? add_76703 : array_index_76697[6];
  assign array_update_76705[7] = add_76613 == 32'h0000_0007 ? add_76703 : array_index_76697[7];
  assign array_update_76705[8] = add_76613 == 32'h0000_0008 ? add_76703 : array_index_76697[8];
  assign array_update_76705[9] = add_76613 == 32'h0000_0009 ? add_76703 : array_index_76697[9];
  assign add_76706 = add_76693 + 32'h0000_0001;
  assign array_update_76707[0] = add_76070 == 32'h0000_0000 ? array_update_76705 : array_update_76694[0];
  assign array_update_76707[1] = add_76070 == 32'h0000_0001 ? array_update_76705 : array_update_76694[1];
  assign array_update_76707[2] = add_76070 == 32'h0000_0002 ? array_update_76705 : array_update_76694[2];
  assign array_update_76707[3] = add_76070 == 32'h0000_0003 ? array_update_76705 : array_update_76694[3];
  assign array_update_76707[4] = add_76070 == 32'h0000_0004 ? array_update_76705 : array_update_76694[4];
  assign array_update_76707[5] = add_76070 == 32'h0000_0005 ? array_update_76705 : array_update_76694[5];
  assign array_update_76707[6] = add_76070 == 32'h0000_0006 ? array_update_76705 : array_update_76694[6];
  assign array_update_76707[7] = add_76070 == 32'h0000_0007 ? array_update_76705 : array_update_76694[7];
  assign array_update_76707[8] = add_76070 == 32'h0000_0008 ? array_update_76705 : array_update_76694[8];
  assign array_update_76707[9] = add_76070 == 32'h0000_0009 ? array_update_76705 : array_update_76694[9];
  assign array_index_76709 = array_update_72021[add_76706 > 32'h0000_0009 ? 4'h9 : add_76706[3:0]];
  assign array_index_76710 = array_update_76707[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_76714 = smul32b_32b_x_32b(array_index_76077[add_76706 > 32'h0000_0009 ? 4'h9 : add_76706[3:0]], array_index_76709[add_76613 > 32'h0000_0009 ? 4'h9 : add_76613[3:0]]);
  assign add_76716 = array_index_76710[add_76613 > 32'h0000_0009 ? 4'h9 : add_76613[3:0]] + smul_76714;
  assign array_update_76718[0] = add_76613 == 32'h0000_0000 ? add_76716 : array_index_76710[0];
  assign array_update_76718[1] = add_76613 == 32'h0000_0001 ? add_76716 : array_index_76710[1];
  assign array_update_76718[2] = add_76613 == 32'h0000_0002 ? add_76716 : array_index_76710[2];
  assign array_update_76718[3] = add_76613 == 32'h0000_0003 ? add_76716 : array_index_76710[3];
  assign array_update_76718[4] = add_76613 == 32'h0000_0004 ? add_76716 : array_index_76710[4];
  assign array_update_76718[5] = add_76613 == 32'h0000_0005 ? add_76716 : array_index_76710[5];
  assign array_update_76718[6] = add_76613 == 32'h0000_0006 ? add_76716 : array_index_76710[6];
  assign array_update_76718[7] = add_76613 == 32'h0000_0007 ? add_76716 : array_index_76710[7];
  assign array_update_76718[8] = add_76613 == 32'h0000_0008 ? add_76716 : array_index_76710[8];
  assign array_update_76718[9] = add_76613 == 32'h0000_0009 ? add_76716 : array_index_76710[9];
  assign add_76719 = add_76706 + 32'h0000_0001;
  assign array_update_76720[0] = add_76070 == 32'h0000_0000 ? array_update_76718 : array_update_76707[0];
  assign array_update_76720[1] = add_76070 == 32'h0000_0001 ? array_update_76718 : array_update_76707[1];
  assign array_update_76720[2] = add_76070 == 32'h0000_0002 ? array_update_76718 : array_update_76707[2];
  assign array_update_76720[3] = add_76070 == 32'h0000_0003 ? array_update_76718 : array_update_76707[3];
  assign array_update_76720[4] = add_76070 == 32'h0000_0004 ? array_update_76718 : array_update_76707[4];
  assign array_update_76720[5] = add_76070 == 32'h0000_0005 ? array_update_76718 : array_update_76707[5];
  assign array_update_76720[6] = add_76070 == 32'h0000_0006 ? array_update_76718 : array_update_76707[6];
  assign array_update_76720[7] = add_76070 == 32'h0000_0007 ? array_update_76718 : array_update_76707[7];
  assign array_update_76720[8] = add_76070 == 32'h0000_0008 ? array_update_76718 : array_update_76707[8];
  assign array_update_76720[9] = add_76070 == 32'h0000_0009 ? array_update_76718 : array_update_76707[9];
  assign array_index_76722 = array_update_72021[add_76719 > 32'h0000_0009 ? 4'h9 : add_76719[3:0]];
  assign array_index_76723 = array_update_76720[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_76727 = smul32b_32b_x_32b(array_index_76077[add_76719 > 32'h0000_0009 ? 4'h9 : add_76719[3:0]], array_index_76722[add_76613 > 32'h0000_0009 ? 4'h9 : add_76613[3:0]]);
  assign add_76729 = array_index_76723[add_76613 > 32'h0000_0009 ? 4'h9 : add_76613[3:0]] + smul_76727;
  assign array_update_76731[0] = add_76613 == 32'h0000_0000 ? add_76729 : array_index_76723[0];
  assign array_update_76731[1] = add_76613 == 32'h0000_0001 ? add_76729 : array_index_76723[1];
  assign array_update_76731[2] = add_76613 == 32'h0000_0002 ? add_76729 : array_index_76723[2];
  assign array_update_76731[3] = add_76613 == 32'h0000_0003 ? add_76729 : array_index_76723[3];
  assign array_update_76731[4] = add_76613 == 32'h0000_0004 ? add_76729 : array_index_76723[4];
  assign array_update_76731[5] = add_76613 == 32'h0000_0005 ? add_76729 : array_index_76723[5];
  assign array_update_76731[6] = add_76613 == 32'h0000_0006 ? add_76729 : array_index_76723[6];
  assign array_update_76731[7] = add_76613 == 32'h0000_0007 ? add_76729 : array_index_76723[7];
  assign array_update_76731[8] = add_76613 == 32'h0000_0008 ? add_76729 : array_index_76723[8];
  assign array_update_76731[9] = add_76613 == 32'h0000_0009 ? add_76729 : array_index_76723[9];
  assign add_76732 = add_76719 + 32'h0000_0001;
  assign array_update_76733[0] = add_76070 == 32'h0000_0000 ? array_update_76731 : array_update_76720[0];
  assign array_update_76733[1] = add_76070 == 32'h0000_0001 ? array_update_76731 : array_update_76720[1];
  assign array_update_76733[2] = add_76070 == 32'h0000_0002 ? array_update_76731 : array_update_76720[2];
  assign array_update_76733[3] = add_76070 == 32'h0000_0003 ? array_update_76731 : array_update_76720[3];
  assign array_update_76733[4] = add_76070 == 32'h0000_0004 ? array_update_76731 : array_update_76720[4];
  assign array_update_76733[5] = add_76070 == 32'h0000_0005 ? array_update_76731 : array_update_76720[5];
  assign array_update_76733[6] = add_76070 == 32'h0000_0006 ? array_update_76731 : array_update_76720[6];
  assign array_update_76733[7] = add_76070 == 32'h0000_0007 ? array_update_76731 : array_update_76720[7];
  assign array_update_76733[8] = add_76070 == 32'h0000_0008 ? array_update_76731 : array_update_76720[8];
  assign array_update_76733[9] = add_76070 == 32'h0000_0009 ? array_update_76731 : array_update_76720[9];
  assign array_index_76735 = array_update_72021[add_76732 > 32'h0000_0009 ? 4'h9 : add_76732[3:0]];
  assign array_index_76736 = array_update_76733[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_76740 = smul32b_32b_x_32b(array_index_76077[add_76732 > 32'h0000_0009 ? 4'h9 : add_76732[3:0]], array_index_76735[add_76613 > 32'h0000_0009 ? 4'h9 : add_76613[3:0]]);
  assign add_76742 = array_index_76736[add_76613 > 32'h0000_0009 ? 4'h9 : add_76613[3:0]] + smul_76740;
  assign array_update_76743[0] = add_76613 == 32'h0000_0000 ? add_76742 : array_index_76736[0];
  assign array_update_76743[1] = add_76613 == 32'h0000_0001 ? add_76742 : array_index_76736[1];
  assign array_update_76743[2] = add_76613 == 32'h0000_0002 ? add_76742 : array_index_76736[2];
  assign array_update_76743[3] = add_76613 == 32'h0000_0003 ? add_76742 : array_index_76736[3];
  assign array_update_76743[4] = add_76613 == 32'h0000_0004 ? add_76742 : array_index_76736[4];
  assign array_update_76743[5] = add_76613 == 32'h0000_0005 ? add_76742 : array_index_76736[5];
  assign array_update_76743[6] = add_76613 == 32'h0000_0006 ? add_76742 : array_index_76736[6];
  assign array_update_76743[7] = add_76613 == 32'h0000_0007 ? add_76742 : array_index_76736[7];
  assign array_update_76743[8] = add_76613 == 32'h0000_0008 ? add_76742 : array_index_76736[8];
  assign array_update_76743[9] = add_76613 == 32'h0000_0009 ? add_76742 : array_index_76736[9];
  assign array_update_76744[0] = add_76070 == 32'h0000_0000 ? array_update_76743 : array_update_76733[0];
  assign array_update_76744[1] = add_76070 == 32'h0000_0001 ? array_update_76743 : array_update_76733[1];
  assign array_update_76744[2] = add_76070 == 32'h0000_0002 ? array_update_76743 : array_update_76733[2];
  assign array_update_76744[3] = add_76070 == 32'h0000_0003 ? array_update_76743 : array_update_76733[3];
  assign array_update_76744[4] = add_76070 == 32'h0000_0004 ? array_update_76743 : array_update_76733[4];
  assign array_update_76744[5] = add_76070 == 32'h0000_0005 ? array_update_76743 : array_update_76733[5];
  assign array_update_76744[6] = add_76070 == 32'h0000_0006 ? array_update_76743 : array_update_76733[6];
  assign array_update_76744[7] = add_76070 == 32'h0000_0007 ? array_update_76743 : array_update_76733[7];
  assign array_update_76744[8] = add_76070 == 32'h0000_0008 ? array_update_76743 : array_update_76733[8];
  assign array_update_76744[9] = add_76070 == 32'h0000_0009 ? array_update_76743 : array_update_76733[9];
  assign array_index_76746 = array_update_76744[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign add_76748 = add_76613 + 32'h0000_0001;
  assign array_update_76749[0] = add_76748 == 32'h0000_0000 ? 32'h0000_0000 : array_index_76746[0];
  assign array_update_76749[1] = add_76748 == 32'h0000_0001 ? 32'h0000_0000 : array_index_76746[1];
  assign array_update_76749[2] = add_76748 == 32'h0000_0002 ? 32'h0000_0000 : array_index_76746[2];
  assign array_update_76749[3] = add_76748 == 32'h0000_0003 ? 32'h0000_0000 : array_index_76746[3];
  assign array_update_76749[4] = add_76748 == 32'h0000_0004 ? 32'h0000_0000 : array_index_76746[4];
  assign array_update_76749[5] = add_76748 == 32'h0000_0005 ? 32'h0000_0000 : array_index_76746[5];
  assign array_update_76749[6] = add_76748 == 32'h0000_0006 ? 32'h0000_0000 : array_index_76746[6];
  assign array_update_76749[7] = add_76748 == 32'h0000_0007 ? 32'h0000_0000 : array_index_76746[7];
  assign array_update_76749[8] = add_76748 == 32'h0000_0008 ? 32'h0000_0000 : array_index_76746[8];
  assign array_update_76749[9] = add_76748 == 32'h0000_0009 ? 32'h0000_0000 : array_index_76746[9];
  assign literal_76750 = 32'h0000_0000;
  assign array_update_76751[0] = add_76070 == 32'h0000_0000 ? array_update_76749 : array_update_76744[0];
  assign array_update_76751[1] = add_76070 == 32'h0000_0001 ? array_update_76749 : array_update_76744[1];
  assign array_update_76751[2] = add_76070 == 32'h0000_0002 ? array_update_76749 : array_update_76744[2];
  assign array_update_76751[3] = add_76070 == 32'h0000_0003 ? array_update_76749 : array_update_76744[3];
  assign array_update_76751[4] = add_76070 == 32'h0000_0004 ? array_update_76749 : array_update_76744[4];
  assign array_update_76751[5] = add_76070 == 32'h0000_0005 ? array_update_76749 : array_update_76744[5];
  assign array_update_76751[6] = add_76070 == 32'h0000_0006 ? array_update_76749 : array_update_76744[6];
  assign array_update_76751[7] = add_76070 == 32'h0000_0007 ? array_update_76749 : array_update_76744[7];
  assign array_update_76751[8] = add_76070 == 32'h0000_0008 ? array_update_76749 : array_update_76744[8];
  assign array_update_76751[9] = add_76070 == 32'h0000_0009 ? array_update_76749 : array_update_76744[9];
  assign array_index_76753 = array_update_72021[literal_76750 > 32'h0000_0009 ? 4'h9 : literal_76750[3:0]];
  assign array_index_76754 = array_update_76751[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_76758 = smul32b_32b_x_32b(array_index_76077[literal_76750 > 32'h0000_0009 ? 4'h9 : literal_76750[3:0]], array_index_76753[add_76748 > 32'h0000_0009 ? 4'h9 : add_76748[3:0]]);
  assign add_76760 = array_index_76754[add_76748 > 32'h0000_0009 ? 4'h9 : add_76748[3:0]] + smul_76758;
  assign array_update_76762[0] = add_76748 == 32'h0000_0000 ? add_76760 : array_index_76754[0];
  assign array_update_76762[1] = add_76748 == 32'h0000_0001 ? add_76760 : array_index_76754[1];
  assign array_update_76762[2] = add_76748 == 32'h0000_0002 ? add_76760 : array_index_76754[2];
  assign array_update_76762[3] = add_76748 == 32'h0000_0003 ? add_76760 : array_index_76754[3];
  assign array_update_76762[4] = add_76748 == 32'h0000_0004 ? add_76760 : array_index_76754[4];
  assign array_update_76762[5] = add_76748 == 32'h0000_0005 ? add_76760 : array_index_76754[5];
  assign array_update_76762[6] = add_76748 == 32'h0000_0006 ? add_76760 : array_index_76754[6];
  assign array_update_76762[7] = add_76748 == 32'h0000_0007 ? add_76760 : array_index_76754[7];
  assign array_update_76762[8] = add_76748 == 32'h0000_0008 ? add_76760 : array_index_76754[8];
  assign array_update_76762[9] = add_76748 == 32'h0000_0009 ? add_76760 : array_index_76754[9];
  assign add_76763 = literal_76750 + 32'h0000_0001;
  assign array_update_76764[0] = add_76070 == 32'h0000_0000 ? array_update_76762 : array_update_76751[0];
  assign array_update_76764[1] = add_76070 == 32'h0000_0001 ? array_update_76762 : array_update_76751[1];
  assign array_update_76764[2] = add_76070 == 32'h0000_0002 ? array_update_76762 : array_update_76751[2];
  assign array_update_76764[3] = add_76070 == 32'h0000_0003 ? array_update_76762 : array_update_76751[3];
  assign array_update_76764[4] = add_76070 == 32'h0000_0004 ? array_update_76762 : array_update_76751[4];
  assign array_update_76764[5] = add_76070 == 32'h0000_0005 ? array_update_76762 : array_update_76751[5];
  assign array_update_76764[6] = add_76070 == 32'h0000_0006 ? array_update_76762 : array_update_76751[6];
  assign array_update_76764[7] = add_76070 == 32'h0000_0007 ? array_update_76762 : array_update_76751[7];
  assign array_update_76764[8] = add_76070 == 32'h0000_0008 ? array_update_76762 : array_update_76751[8];
  assign array_update_76764[9] = add_76070 == 32'h0000_0009 ? array_update_76762 : array_update_76751[9];
  assign array_index_76766 = array_update_72021[add_76763 > 32'h0000_0009 ? 4'h9 : add_76763[3:0]];
  assign array_index_76767 = array_update_76764[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_76771 = smul32b_32b_x_32b(array_index_76077[add_76763 > 32'h0000_0009 ? 4'h9 : add_76763[3:0]], array_index_76766[add_76748 > 32'h0000_0009 ? 4'h9 : add_76748[3:0]]);
  assign add_76773 = array_index_76767[add_76748 > 32'h0000_0009 ? 4'h9 : add_76748[3:0]] + smul_76771;
  assign array_update_76775[0] = add_76748 == 32'h0000_0000 ? add_76773 : array_index_76767[0];
  assign array_update_76775[1] = add_76748 == 32'h0000_0001 ? add_76773 : array_index_76767[1];
  assign array_update_76775[2] = add_76748 == 32'h0000_0002 ? add_76773 : array_index_76767[2];
  assign array_update_76775[3] = add_76748 == 32'h0000_0003 ? add_76773 : array_index_76767[3];
  assign array_update_76775[4] = add_76748 == 32'h0000_0004 ? add_76773 : array_index_76767[4];
  assign array_update_76775[5] = add_76748 == 32'h0000_0005 ? add_76773 : array_index_76767[5];
  assign array_update_76775[6] = add_76748 == 32'h0000_0006 ? add_76773 : array_index_76767[6];
  assign array_update_76775[7] = add_76748 == 32'h0000_0007 ? add_76773 : array_index_76767[7];
  assign array_update_76775[8] = add_76748 == 32'h0000_0008 ? add_76773 : array_index_76767[8];
  assign array_update_76775[9] = add_76748 == 32'h0000_0009 ? add_76773 : array_index_76767[9];
  assign add_76776 = add_76763 + 32'h0000_0001;
  assign array_update_76777[0] = add_76070 == 32'h0000_0000 ? array_update_76775 : array_update_76764[0];
  assign array_update_76777[1] = add_76070 == 32'h0000_0001 ? array_update_76775 : array_update_76764[1];
  assign array_update_76777[2] = add_76070 == 32'h0000_0002 ? array_update_76775 : array_update_76764[2];
  assign array_update_76777[3] = add_76070 == 32'h0000_0003 ? array_update_76775 : array_update_76764[3];
  assign array_update_76777[4] = add_76070 == 32'h0000_0004 ? array_update_76775 : array_update_76764[4];
  assign array_update_76777[5] = add_76070 == 32'h0000_0005 ? array_update_76775 : array_update_76764[5];
  assign array_update_76777[6] = add_76070 == 32'h0000_0006 ? array_update_76775 : array_update_76764[6];
  assign array_update_76777[7] = add_76070 == 32'h0000_0007 ? array_update_76775 : array_update_76764[7];
  assign array_update_76777[8] = add_76070 == 32'h0000_0008 ? array_update_76775 : array_update_76764[8];
  assign array_update_76777[9] = add_76070 == 32'h0000_0009 ? array_update_76775 : array_update_76764[9];
  assign array_index_76779 = array_update_72021[add_76776 > 32'h0000_0009 ? 4'h9 : add_76776[3:0]];
  assign array_index_76780 = array_update_76777[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_76784 = smul32b_32b_x_32b(array_index_76077[add_76776 > 32'h0000_0009 ? 4'h9 : add_76776[3:0]], array_index_76779[add_76748 > 32'h0000_0009 ? 4'h9 : add_76748[3:0]]);
  assign add_76786 = array_index_76780[add_76748 > 32'h0000_0009 ? 4'h9 : add_76748[3:0]] + smul_76784;
  assign array_update_76788[0] = add_76748 == 32'h0000_0000 ? add_76786 : array_index_76780[0];
  assign array_update_76788[1] = add_76748 == 32'h0000_0001 ? add_76786 : array_index_76780[1];
  assign array_update_76788[2] = add_76748 == 32'h0000_0002 ? add_76786 : array_index_76780[2];
  assign array_update_76788[3] = add_76748 == 32'h0000_0003 ? add_76786 : array_index_76780[3];
  assign array_update_76788[4] = add_76748 == 32'h0000_0004 ? add_76786 : array_index_76780[4];
  assign array_update_76788[5] = add_76748 == 32'h0000_0005 ? add_76786 : array_index_76780[5];
  assign array_update_76788[6] = add_76748 == 32'h0000_0006 ? add_76786 : array_index_76780[6];
  assign array_update_76788[7] = add_76748 == 32'h0000_0007 ? add_76786 : array_index_76780[7];
  assign array_update_76788[8] = add_76748 == 32'h0000_0008 ? add_76786 : array_index_76780[8];
  assign array_update_76788[9] = add_76748 == 32'h0000_0009 ? add_76786 : array_index_76780[9];
  assign add_76789 = add_76776 + 32'h0000_0001;
  assign array_update_76790[0] = add_76070 == 32'h0000_0000 ? array_update_76788 : array_update_76777[0];
  assign array_update_76790[1] = add_76070 == 32'h0000_0001 ? array_update_76788 : array_update_76777[1];
  assign array_update_76790[2] = add_76070 == 32'h0000_0002 ? array_update_76788 : array_update_76777[2];
  assign array_update_76790[3] = add_76070 == 32'h0000_0003 ? array_update_76788 : array_update_76777[3];
  assign array_update_76790[4] = add_76070 == 32'h0000_0004 ? array_update_76788 : array_update_76777[4];
  assign array_update_76790[5] = add_76070 == 32'h0000_0005 ? array_update_76788 : array_update_76777[5];
  assign array_update_76790[6] = add_76070 == 32'h0000_0006 ? array_update_76788 : array_update_76777[6];
  assign array_update_76790[7] = add_76070 == 32'h0000_0007 ? array_update_76788 : array_update_76777[7];
  assign array_update_76790[8] = add_76070 == 32'h0000_0008 ? array_update_76788 : array_update_76777[8];
  assign array_update_76790[9] = add_76070 == 32'h0000_0009 ? array_update_76788 : array_update_76777[9];
  assign array_index_76792 = array_update_72021[add_76789 > 32'h0000_0009 ? 4'h9 : add_76789[3:0]];
  assign array_index_76793 = array_update_76790[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_76797 = smul32b_32b_x_32b(array_index_76077[add_76789 > 32'h0000_0009 ? 4'h9 : add_76789[3:0]], array_index_76792[add_76748 > 32'h0000_0009 ? 4'h9 : add_76748[3:0]]);
  assign add_76799 = array_index_76793[add_76748 > 32'h0000_0009 ? 4'h9 : add_76748[3:0]] + smul_76797;
  assign array_update_76801[0] = add_76748 == 32'h0000_0000 ? add_76799 : array_index_76793[0];
  assign array_update_76801[1] = add_76748 == 32'h0000_0001 ? add_76799 : array_index_76793[1];
  assign array_update_76801[2] = add_76748 == 32'h0000_0002 ? add_76799 : array_index_76793[2];
  assign array_update_76801[3] = add_76748 == 32'h0000_0003 ? add_76799 : array_index_76793[3];
  assign array_update_76801[4] = add_76748 == 32'h0000_0004 ? add_76799 : array_index_76793[4];
  assign array_update_76801[5] = add_76748 == 32'h0000_0005 ? add_76799 : array_index_76793[5];
  assign array_update_76801[6] = add_76748 == 32'h0000_0006 ? add_76799 : array_index_76793[6];
  assign array_update_76801[7] = add_76748 == 32'h0000_0007 ? add_76799 : array_index_76793[7];
  assign array_update_76801[8] = add_76748 == 32'h0000_0008 ? add_76799 : array_index_76793[8];
  assign array_update_76801[9] = add_76748 == 32'h0000_0009 ? add_76799 : array_index_76793[9];
  assign add_76802 = add_76789 + 32'h0000_0001;
  assign array_update_76803[0] = add_76070 == 32'h0000_0000 ? array_update_76801 : array_update_76790[0];
  assign array_update_76803[1] = add_76070 == 32'h0000_0001 ? array_update_76801 : array_update_76790[1];
  assign array_update_76803[2] = add_76070 == 32'h0000_0002 ? array_update_76801 : array_update_76790[2];
  assign array_update_76803[3] = add_76070 == 32'h0000_0003 ? array_update_76801 : array_update_76790[3];
  assign array_update_76803[4] = add_76070 == 32'h0000_0004 ? array_update_76801 : array_update_76790[4];
  assign array_update_76803[5] = add_76070 == 32'h0000_0005 ? array_update_76801 : array_update_76790[5];
  assign array_update_76803[6] = add_76070 == 32'h0000_0006 ? array_update_76801 : array_update_76790[6];
  assign array_update_76803[7] = add_76070 == 32'h0000_0007 ? array_update_76801 : array_update_76790[7];
  assign array_update_76803[8] = add_76070 == 32'h0000_0008 ? array_update_76801 : array_update_76790[8];
  assign array_update_76803[9] = add_76070 == 32'h0000_0009 ? array_update_76801 : array_update_76790[9];
  assign array_index_76805 = array_update_72021[add_76802 > 32'h0000_0009 ? 4'h9 : add_76802[3:0]];
  assign array_index_76806 = array_update_76803[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_76810 = smul32b_32b_x_32b(array_index_76077[add_76802 > 32'h0000_0009 ? 4'h9 : add_76802[3:0]], array_index_76805[add_76748 > 32'h0000_0009 ? 4'h9 : add_76748[3:0]]);
  assign add_76812 = array_index_76806[add_76748 > 32'h0000_0009 ? 4'h9 : add_76748[3:0]] + smul_76810;
  assign array_update_76814[0] = add_76748 == 32'h0000_0000 ? add_76812 : array_index_76806[0];
  assign array_update_76814[1] = add_76748 == 32'h0000_0001 ? add_76812 : array_index_76806[1];
  assign array_update_76814[2] = add_76748 == 32'h0000_0002 ? add_76812 : array_index_76806[2];
  assign array_update_76814[3] = add_76748 == 32'h0000_0003 ? add_76812 : array_index_76806[3];
  assign array_update_76814[4] = add_76748 == 32'h0000_0004 ? add_76812 : array_index_76806[4];
  assign array_update_76814[5] = add_76748 == 32'h0000_0005 ? add_76812 : array_index_76806[5];
  assign array_update_76814[6] = add_76748 == 32'h0000_0006 ? add_76812 : array_index_76806[6];
  assign array_update_76814[7] = add_76748 == 32'h0000_0007 ? add_76812 : array_index_76806[7];
  assign array_update_76814[8] = add_76748 == 32'h0000_0008 ? add_76812 : array_index_76806[8];
  assign array_update_76814[9] = add_76748 == 32'h0000_0009 ? add_76812 : array_index_76806[9];
  assign add_76815 = add_76802 + 32'h0000_0001;
  assign array_update_76816[0] = add_76070 == 32'h0000_0000 ? array_update_76814 : array_update_76803[0];
  assign array_update_76816[1] = add_76070 == 32'h0000_0001 ? array_update_76814 : array_update_76803[1];
  assign array_update_76816[2] = add_76070 == 32'h0000_0002 ? array_update_76814 : array_update_76803[2];
  assign array_update_76816[3] = add_76070 == 32'h0000_0003 ? array_update_76814 : array_update_76803[3];
  assign array_update_76816[4] = add_76070 == 32'h0000_0004 ? array_update_76814 : array_update_76803[4];
  assign array_update_76816[5] = add_76070 == 32'h0000_0005 ? array_update_76814 : array_update_76803[5];
  assign array_update_76816[6] = add_76070 == 32'h0000_0006 ? array_update_76814 : array_update_76803[6];
  assign array_update_76816[7] = add_76070 == 32'h0000_0007 ? array_update_76814 : array_update_76803[7];
  assign array_update_76816[8] = add_76070 == 32'h0000_0008 ? array_update_76814 : array_update_76803[8];
  assign array_update_76816[9] = add_76070 == 32'h0000_0009 ? array_update_76814 : array_update_76803[9];
  assign array_index_76818 = array_update_72021[add_76815 > 32'h0000_0009 ? 4'h9 : add_76815[3:0]];
  assign array_index_76819 = array_update_76816[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_76823 = smul32b_32b_x_32b(array_index_76077[add_76815 > 32'h0000_0009 ? 4'h9 : add_76815[3:0]], array_index_76818[add_76748 > 32'h0000_0009 ? 4'h9 : add_76748[3:0]]);
  assign add_76825 = array_index_76819[add_76748 > 32'h0000_0009 ? 4'h9 : add_76748[3:0]] + smul_76823;
  assign array_update_76827[0] = add_76748 == 32'h0000_0000 ? add_76825 : array_index_76819[0];
  assign array_update_76827[1] = add_76748 == 32'h0000_0001 ? add_76825 : array_index_76819[1];
  assign array_update_76827[2] = add_76748 == 32'h0000_0002 ? add_76825 : array_index_76819[2];
  assign array_update_76827[3] = add_76748 == 32'h0000_0003 ? add_76825 : array_index_76819[3];
  assign array_update_76827[4] = add_76748 == 32'h0000_0004 ? add_76825 : array_index_76819[4];
  assign array_update_76827[5] = add_76748 == 32'h0000_0005 ? add_76825 : array_index_76819[5];
  assign array_update_76827[6] = add_76748 == 32'h0000_0006 ? add_76825 : array_index_76819[6];
  assign array_update_76827[7] = add_76748 == 32'h0000_0007 ? add_76825 : array_index_76819[7];
  assign array_update_76827[8] = add_76748 == 32'h0000_0008 ? add_76825 : array_index_76819[8];
  assign array_update_76827[9] = add_76748 == 32'h0000_0009 ? add_76825 : array_index_76819[9];
  assign add_76828 = add_76815 + 32'h0000_0001;
  assign array_update_76829[0] = add_76070 == 32'h0000_0000 ? array_update_76827 : array_update_76816[0];
  assign array_update_76829[1] = add_76070 == 32'h0000_0001 ? array_update_76827 : array_update_76816[1];
  assign array_update_76829[2] = add_76070 == 32'h0000_0002 ? array_update_76827 : array_update_76816[2];
  assign array_update_76829[3] = add_76070 == 32'h0000_0003 ? array_update_76827 : array_update_76816[3];
  assign array_update_76829[4] = add_76070 == 32'h0000_0004 ? array_update_76827 : array_update_76816[4];
  assign array_update_76829[5] = add_76070 == 32'h0000_0005 ? array_update_76827 : array_update_76816[5];
  assign array_update_76829[6] = add_76070 == 32'h0000_0006 ? array_update_76827 : array_update_76816[6];
  assign array_update_76829[7] = add_76070 == 32'h0000_0007 ? array_update_76827 : array_update_76816[7];
  assign array_update_76829[8] = add_76070 == 32'h0000_0008 ? array_update_76827 : array_update_76816[8];
  assign array_update_76829[9] = add_76070 == 32'h0000_0009 ? array_update_76827 : array_update_76816[9];
  assign array_index_76831 = array_update_72021[add_76828 > 32'h0000_0009 ? 4'h9 : add_76828[3:0]];
  assign array_index_76832 = array_update_76829[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_76836 = smul32b_32b_x_32b(array_index_76077[add_76828 > 32'h0000_0009 ? 4'h9 : add_76828[3:0]], array_index_76831[add_76748 > 32'h0000_0009 ? 4'h9 : add_76748[3:0]]);
  assign add_76838 = array_index_76832[add_76748 > 32'h0000_0009 ? 4'h9 : add_76748[3:0]] + smul_76836;
  assign array_update_76840[0] = add_76748 == 32'h0000_0000 ? add_76838 : array_index_76832[0];
  assign array_update_76840[1] = add_76748 == 32'h0000_0001 ? add_76838 : array_index_76832[1];
  assign array_update_76840[2] = add_76748 == 32'h0000_0002 ? add_76838 : array_index_76832[2];
  assign array_update_76840[3] = add_76748 == 32'h0000_0003 ? add_76838 : array_index_76832[3];
  assign array_update_76840[4] = add_76748 == 32'h0000_0004 ? add_76838 : array_index_76832[4];
  assign array_update_76840[5] = add_76748 == 32'h0000_0005 ? add_76838 : array_index_76832[5];
  assign array_update_76840[6] = add_76748 == 32'h0000_0006 ? add_76838 : array_index_76832[6];
  assign array_update_76840[7] = add_76748 == 32'h0000_0007 ? add_76838 : array_index_76832[7];
  assign array_update_76840[8] = add_76748 == 32'h0000_0008 ? add_76838 : array_index_76832[8];
  assign array_update_76840[9] = add_76748 == 32'h0000_0009 ? add_76838 : array_index_76832[9];
  assign add_76841 = add_76828 + 32'h0000_0001;
  assign array_update_76842[0] = add_76070 == 32'h0000_0000 ? array_update_76840 : array_update_76829[0];
  assign array_update_76842[1] = add_76070 == 32'h0000_0001 ? array_update_76840 : array_update_76829[1];
  assign array_update_76842[2] = add_76070 == 32'h0000_0002 ? array_update_76840 : array_update_76829[2];
  assign array_update_76842[3] = add_76070 == 32'h0000_0003 ? array_update_76840 : array_update_76829[3];
  assign array_update_76842[4] = add_76070 == 32'h0000_0004 ? array_update_76840 : array_update_76829[4];
  assign array_update_76842[5] = add_76070 == 32'h0000_0005 ? array_update_76840 : array_update_76829[5];
  assign array_update_76842[6] = add_76070 == 32'h0000_0006 ? array_update_76840 : array_update_76829[6];
  assign array_update_76842[7] = add_76070 == 32'h0000_0007 ? array_update_76840 : array_update_76829[7];
  assign array_update_76842[8] = add_76070 == 32'h0000_0008 ? array_update_76840 : array_update_76829[8];
  assign array_update_76842[9] = add_76070 == 32'h0000_0009 ? array_update_76840 : array_update_76829[9];
  assign array_index_76844 = array_update_72021[add_76841 > 32'h0000_0009 ? 4'h9 : add_76841[3:0]];
  assign array_index_76845 = array_update_76842[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_76849 = smul32b_32b_x_32b(array_index_76077[add_76841 > 32'h0000_0009 ? 4'h9 : add_76841[3:0]], array_index_76844[add_76748 > 32'h0000_0009 ? 4'h9 : add_76748[3:0]]);
  assign add_76851 = array_index_76845[add_76748 > 32'h0000_0009 ? 4'h9 : add_76748[3:0]] + smul_76849;
  assign array_update_76853[0] = add_76748 == 32'h0000_0000 ? add_76851 : array_index_76845[0];
  assign array_update_76853[1] = add_76748 == 32'h0000_0001 ? add_76851 : array_index_76845[1];
  assign array_update_76853[2] = add_76748 == 32'h0000_0002 ? add_76851 : array_index_76845[2];
  assign array_update_76853[3] = add_76748 == 32'h0000_0003 ? add_76851 : array_index_76845[3];
  assign array_update_76853[4] = add_76748 == 32'h0000_0004 ? add_76851 : array_index_76845[4];
  assign array_update_76853[5] = add_76748 == 32'h0000_0005 ? add_76851 : array_index_76845[5];
  assign array_update_76853[6] = add_76748 == 32'h0000_0006 ? add_76851 : array_index_76845[6];
  assign array_update_76853[7] = add_76748 == 32'h0000_0007 ? add_76851 : array_index_76845[7];
  assign array_update_76853[8] = add_76748 == 32'h0000_0008 ? add_76851 : array_index_76845[8];
  assign array_update_76853[9] = add_76748 == 32'h0000_0009 ? add_76851 : array_index_76845[9];
  assign add_76854 = add_76841 + 32'h0000_0001;
  assign array_update_76855[0] = add_76070 == 32'h0000_0000 ? array_update_76853 : array_update_76842[0];
  assign array_update_76855[1] = add_76070 == 32'h0000_0001 ? array_update_76853 : array_update_76842[1];
  assign array_update_76855[2] = add_76070 == 32'h0000_0002 ? array_update_76853 : array_update_76842[2];
  assign array_update_76855[3] = add_76070 == 32'h0000_0003 ? array_update_76853 : array_update_76842[3];
  assign array_update_76855[4] = add_76070 == 32'h0000_0004 ? array_update_76853 : array_update_76842[4];
  assign array_update_76855[5] = add_76070 == 32'h0000_0005 ? array_update_76853 : array_update_76842[5];
  assign array_update_76855[6] = add_76070 == 32'h0000_0006 ? array_update_76853 : array_update_76842[6];
  assign array_update_76855[7] = add_76070 == 32'h0000_0007 ? array_update_76853 : array_update_76842[7];
  assign array_update_76855[8] = add_76070 == 32'h0000_0008 ? array_update_76853 : array_update_76842[8];
  assign array_update_76855[9] = add_76070 == 32'h0000_0009 ? array_update_76853 : array_update_76842[9];
  assign array_index_76857 = array_update_72021[add_76854 > 32'h0000_0009 ? 4'h9 : add_76854[3:0]];
  assign array_index_76858 = array_update_76855[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_76862 = smul32b_32b_x_32b(array_index_76077[add_76854 > 32'h0000_0009 ? 4'h9 : add_76854[3:0]], array_index_76857[add_76748 > 32'h0000_0009 ? 4'h9 : add_76748[3:0]]);
  assign add_76864 = array_index_76858[add_76748 > 32'h0000_0009 ? 4'h9 : add_76748[3:0]] + smul_76862;
  assign array_update_76866[0] = add_76748 == 32'h0000_0000 ? add_76864 : array_index_76858[0];
  assign array_update_76866[1] = add_76748 == 32'h0000_0001 ? add_76864 : array_index_76858[1];
  assign array_update_76866[2] = add_76748 == 32'h0000_0002 ? add_76864 : array_index_76858[2];
  assign array_update_76866[3] = add_76748 == 32'h0000_0003 ? add_76864 : array_index_76858[3];
  assign array_update_76866[4] = add_76748 == 32'h0000_0004 ? add_76864 : array_index_76858[4];
  assign array_update_76866[5] = add_76748 == 32'h0000_0005 ? add_76864 : array_index_76858[5];
  assign array_update_76866[6] = add_76748 == 32'h0000_0006 ? add_76864 : array_index_76858[6];
  assign array_update_76866[7] = add_76748 == 32'h0000_0007 ? add_76864 : array_index_76858[7];
  assign array_update_76866[8] = add_76748 == 32'h0000_0008 ? add_76864 : array_index_76858[8];
  assign array_update_76866[9] = add_76748 == 32'h0000_0009 ? add_76864 : array_index_76858[9];
  assign add_76867 = add_76854 + 32'h0000_0001;
  assign array_update_76868[0] = add_76070 == 32'h0000_0000 ? array_update_76866 : array_update_76855[0];
  assign array_update_76868[1] = add_76070 == 32'h0000_0001 ? array_update_76866 : array_update_76855[1];
  assign array_update_76868[2] = add_76070 == 32'h0000_0002 ? array_update_76866 : array_update_76855[2];
  assign array_update_76868[3] = add_76070 == 32'h0000_0003 ? array_update_76866 : array_update_76855[3];
  assign array_update_76868[4] = add_76070 == 32'h0000_0004 ? array_update_76866 : array_update_76855[4];
  assign array_update_76868[5] = add_76070 == 32'h0000_0005 ? array_update_76866 : array_update_76855[5];
  assign array_update_76868[6] = add_76070 == 32'h0000_0006 ? array_update_76866 : array_update_76855[6];
  assign array_update_76868[7] = add_76070 == 32'h0000_0007 ? array_update_76866 : array_update_76855[7];
  assign array_update_76868[8] = add_76070 == 32'h0000_0008 ? array_update_76866 : array_update_76855[8];
  assign array_update_76868[9] = add_76070 == 32'h0000_0009 ? array_update_76866 : array_update_76855[9];
  assign array_index_76870 = array_update_72021[add_76867 > 32'h0000_0009 ? 4'h9 : add_76867[3:0]];
  assign array_index_76871 = array_update_76868[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_76875 = smul32b_32b_x_32b(array_index_76077[add_76867 > 32'h0000_0009 ? 4'h9 : add_76867[3:0]], array_index_76870[add_76748 > 32'h0000_0009 ? 4'h9 : add_76748[3:0]]);
  assign add_76877 = array_index_76871[add_76748 > 32'h0000_0009 ? 4'h9 : add_76748[3:0]] + smul_76875;
  assign array_update_76878[0] = add_76748 == 32'h0000_0000 ? add_76877 : array_index_76871[0];
  assign array_update_76878[1] = add_76748 == 32'h0000_0001 ? add_76877 : array_index_76871[1];
  assign array_update_76878[2] = add_76748 == 32'h0000_0002 ? add_76877 : array_index_76871[2];
  assign array_update_76878[3] = add_76748 == 32'h0000_0003 ? add_76877 : array_index_76871[3];
  assign array_update_76878[4] = add_76748 == 32'h0000_0004 ? add_76877 : array_index_76871[4];
  assign array_update_76878[5] = add_76748 == 32'h0000_0005 ? add_76877 : array_index_76871[5];
  assign array_update_76878[6] = add_76748 == 32'h0000_0006 ? add_76877 : array_index_76871[6];
  assign array_update_76878[7] = add_76748 == 32'h0000_0007 ? add_76877 : array_index_76871[7];
  assign array_update_76878[8] = add_76748 == 32'h0000_0008 ? add_76877 : array_index_76871[8];
  assign array_update_76878[9] = add_76748 == 32'h0000_0009 ? add_76877 : array_index_76871[9];
  assign array_update_76879[0] = add_76070 == 32'h0000_0000 ? array_update_76878 : array_update_76868[0];
  assign array_update_76879[1] = add_76070 == 32'h0000_0001 ? array_update_76878 : array_update_76868[1];
  assign array_update_76879[2] = add_76070 == 32'h0000_0002 ? array_update_76878 : array_update_76868[2];
  assign array_update_76879[3] = add_76070 == 32'h0000_0003 ? array_update_76878 : array_update_76868[3];
  assign array_update_76879[4] = add_76070 == 32'h0000_0004 ? array_update_76878 : array_update_76868[4];
  assign array_update_76879[5] = add_76070 == 32'h0000_0005 ? array_update_76878 : array_update_76868[5];
  assign array_update_76879[6] = add_76070 == 32'h0000_0006 ? array_update_76878 : array_update_76868[6];
  assign array_update_76879[7] = add_76070 == 32'h0000_0007 ? array_update_76878 : array_update_76868[7];
  assign array_update_76879[8] = add_76070 == 32'h0000_0008 ? array_update_76878 : array_update_76868[8];
  assign array_update_76879[9] = add_76070 == 32'h0000_0009 ? array_update_76878 : array_update_76868[9];
  assign array_index_76881 = array_update_76879[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign add_76883 = add_76748 + 32'h0000_0001;
  assign array_update_76884[0] = add_76883 == 32'h0000_0000 ? 32'h0000_0000 : array_index_76881[0];
  assign array_update_76884[1] = add_76883 == 32'h0000_0001 ? 32'h0000_0000 : array_index_76881[1];
  assign array_update_76884[2] = add_76883 == 32'h0000_0002 ? 32'h0000_0000 : array_index_76881[2];
  assign array_update_76884[3] = add_76883 == 32'h0000_0003 ? 32'h0000_0000 : array_index_76881[3];
  assign array_update_76884[4] = add_76883 == 32'h0000_0004 ? 32'h0000_0000 : array_index_76881[4];
  assign array_update_76884[5] = add_76883 == 32'h0000_0005 ? 32'h0000_0000 : array_index_76881[5];
  assign array_update_76884[6] = add_76883 == 32'h0000_0006 ? 32'h0000_0000 : array_index_76881[6];
  assign array_update_76884[7] = add_76883 == 32'h0000_0007 ? 32'h0000_0000 : array_index_76881[7];
  assign array_update_76884[8] = add_76883 == 32'h0000_0008 ? 32'h0000_0000 : array_index_76881[8];
  assign array_update_76884[9] = add_76883 == 32'h0000_0009 ? 32'h0000_0000 : array_index_76881[9];
  assign literal_76885 = 32'h0000_0000;
  assign array_update_76886[0] = add_76070 == 32'h0000_0000 ? array_update_76884 : array_update_76879[0];
  assign array_update_76886[1] = add_76070 == 32'h0000_0001 ? array_update_76884 : array_update_76879[1];
  assign array_update_76886[2] = add_76070 == 32'h0000_0002 ? array_update_76884 : array_update_76879[2];
  assign array_update_76886[3] = add_76070 == 32'h0000_0003 ? array_update_76884 : array_update_76879[3];
  assign array_update_76886[4] = add_76070 == 32'h0000_0004 ? array_update_76884 : array_update_76879[4];
  assign array_update_76886[5] = add_76070 == 32'h0000_0005 ? array_update_76884 : array_update_76879[5];
  assign array_update_76886[6] = add_76070 == 32'h0000_0006 ? array_update_76884 : array_update_76879[6];
  assign array_update_76886[7] = add_76070 == 32'h0000_0007 ? array_update_76884 : array_update_76879[7];
  assign array_update_76886[8] = add_76070 == 32'h0000_0008 ? array_update_76884 : array_update_76879[8];
  assign array_update_76886[9] = add_76070 == 32'h0000_0009 ? array_update_76884 : array_update_76879[9];
  assign array_index_76888 = array_update_72021[literal_76885 > 32'h0000_0009 ? 4'h9 : literal_76885[3:0]];
  assign array_index_76889 = array_update_76886[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_76893 = smul32b_32b_x_32b(array_index_76077[literal_76885 > 32'h0000_0009 ? 4'h9 : literal_76885[3:0]], array_index_76888[add_76883 > 32'h0000_0009 ? 4'h9 : add_76883[3:0]]);
  assign add_76895 = array_index_76889[add_76883 > 32'h0000_0009 ? 4'h9 : add_76883[3:0]] + smul_76893;
  assign array_update_76897[0] = add_76883 == 32'h0000_0000 ? add_76895 : array_index_76889[0];
  assign array_update_76897[1] = add_76883 == 32'h0000_0001 ? add_76895 : array_index_76889[1];
  assign array_update_76897[2] = add_76883 == 32'h0000_0002 ? add_76895 : array_index_76889[2];
  assign array_update_76897[3] = add_76883 == 32'h0000_0003 ? add_76895 : array_index_76889[3];
  assign array_update_76897[4] = add_76883 == 32'h0000_0004 ? add_76895 : array_index_76889[4];
  assign array_update_76897[5] = add_76883 == 32'h0000_0005 ? add_76895 : array_index_76889[5];
  assign array_update_76897[6] = add_76883 == 32'h0000_0006 ? add_76895 : array_index_76889[6];
  assign array_update_76897[7] = add_76883 == 32'h0000_0007 ? add_76895 : array_index_76889[7];
  assign array_update_76897[8] = add_76883 == 32'h0000_0008 ? add_76895 : array_index_76889[8];
  assign array_update_76897[9] = add_76883 == 32'h0000_0009 ? add_76895 : array_index_76889[9];
  assign add_76898 = literal_76885 + 32'h0000_0001;
  assign array_update_76899[0] = add_76070 == 32'h0000_0000 ? array_update_76897 : array_update_76886[0];
  assign array_update_76899[1] = add_76070 == 32'h0000_0001 ? array_update_76897 : array_update_76886[1];
  assign array_update_76899[2] = add_76070 == 32'h0000_0002 ? array_update_76897 : array_update_76886[2];
  assign array_update_76899[3] = add_76070 == 32'h0000_0003 ? array_update_76897 : array_update_76886[3];
  assign array_update_76899[4] = add_76070 == 32'h0000_0004 ? array_update_76897 : array_update_76886[4];
  assign array_update_76899[5] = add_76070 == 32'h0000_0005 ? array_update_76897 : array_update_76886[5];
  assign array_update_76899[6] = add_76070 == 32'h0000_0006 ? array_update_76897 : array_update_76886[6];
  assign array_update_76899[7] = add_76070 == 32'h0000_0007 ? array_update_76897 : array_update_76886[7];
  assign array_update_76899[8] = add_76070 == 32'h0000_0008 ? array_update_76897 : array_update_76886[8];
  assign array_update_76899[9] = add_76070 == 32'h0000_0009 ? array_update_76897 : array_update_76886[9];
  assign array_index_76901 = array_update_72021[add_76898 > 32'h0000_0009 ? 4'h9 : add_76898[3:0]];
  assign array_index_76902 = array_update_76899[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_76906 = smul32b_32b_x_32b(array_index_76077[add_76898 > 32'h0000_0009 ? 4'h9 : add_76898[3:0]], array_index_76901[add_76883 > 32'h0000_0009 ? 4'h9 : add_76883[3:0]]);
  assign add_76908 = array_index_76902[add_76883 > 32'h0000_0009 ? 4'h9 : add_76883[3:0]] + smul_76906;
  assign array_update_76910[0] = add_76883 == 32'h0000_0000 ? add_76908 : array_index_76902[0];
  assign array_update_76910[1] = add_76883 == 32'h0000_0001 ? add_76908 : array_index_76902[1];
  assign array_update_76910[2] = add_76883 == 32'h0000_0002 ? add_76908 : array_index_76902[2];
  assign array_update_76910[3] = add_76883 == 32'h0000_0003 ? add_76908 : array_index_76902[3];
  assign array_update_76910[4] = add_76883 == 32'h0000_0004 ? add_76908 : array_index_76902[4];
  assign array_update_76910[5] = add_76883 == 32'h0000_0005 ? add_76908 : array_index_76902[5];
  assign array_update_76910[6] = add_76883 == 32'h0000_0006 ? add_76908 : array_index_76902[6];
  assign array_update_76910[7] = add_76883 == 32'h0000_0007 ? add_76908 : array_index_76902[7];
  assign array_update_76910[8] = add_76883 == 32'h0000_0008 ? add_76908 : array_index_76902[8];
  assign array_update_76910[9] = add_76883 == 32'h0000_0009 ? add_76908 : array_index_76902[9];
  assign add_76911 = add_76898 + 32'h0000_0001;
  assign array_update_76912[0] = add_76070 == 32'h0000_0000 ? array_update_76910 : array_update_76899[0];
  assign array_update_76912[1] = add_76070 == 32'h0000_0001 ? array_update_76910 : array_update_76899[1];
  assign array_update_76912[2] = add_76070 == 32'h0000_0002 ? array_update_76910 : array_update_76899[2];
  assign array_update_76912[3] = add_76070 == 32'h0000_0003 ? array_update_76910 : array_update_76899[3];
  assign array_update_76912[4] = add_76070 == 32'h0000_0004 ? array_update_76910 : array_update_76899[4];
  assign array_update_76912[5] = add_76070 == 32'h0000_0005 ? array_update_76910 : array_update_76899[5];
  assign array_update_76912[6] = add_76070 == 32'h0000_0006 ? array_update_76910 : array_update_76899[6];
  assign array_update_76912[7] = add_76070 == 32'h0000_0007 ? array_update_76910 : array_update_76899[7];
  assign array_update_76912[8] = add_76070 == 32'h0000_0008 ? array_update_76910 : array_update_76899[8];
  assign array_update_76912[9] = add_76070 == 32'h0000_0009 ? array_update_76910 : array_update_76899[9];
  assign array_index_76914 = array_update_72021[add_76911 > 32'h0000_0009 ? 4'h9 : add_76911[3:0]];
  assign array_index_76915 = array_update_76912[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_76919 = smul32b_32b_x_32b(array_index_76077[add_76911 > 32'h0000_0009 ? 4'h9 : add_76911[3:0]], array_index_76914[add_76883 > 32'h0000_0009 ? 4'h9 : add_76883[3:0]]);
  assign add_76921 = array_index_76915[add_76883 > 32'h0000_0009 ? 4'h9 : add_76883[3:0]] + smul_76919;
  assign array_update_76923[0] = add_76883 == 32'h0000_0000 ? add_76921 : array_index_76915[0];
  assign array_update_76923[1] = add_76883 == 32'h0000_0001 ? add_76921 : array_index_76915[1];
  assign array_update_76923[2] = add_76883 == 32'h0000_0002 ? add_76921 : array_index_76915[2];
  assign array_update_76923[3] = add_76883 == 32'h0000_0003 ? add_76921 : array_index_76915[3];
  assign array_update_76923[4] = add_76883 == 32'h0000_0004 ? add_76921 : array_index_76915[4];
  assign array_update_76923[5] = add_76883 == 32'h0000_0005 ? add_76921 : array_index_76915[5];
  assign array_update_76923[6] = add_76883 == 32'h0000_0006 ? add_76921 : array_index_76915[6];
  assign array_update_76923[7] = add_76883 == 32'h0000_0007 ? add_76921 : array_index_76915[7];
  assign array_update_76923[8] = add_76883 == 32'h0000_0008 ? add_76921 : array_index_76915[8];
  assign array_update_76923[9] = add_76883 == 32'h0000_0009 ? add_76921 : array_index_76915[9];
  assign add_76924 = add_76911 + 32'h0000_0001;
  assign array_update_76925[0] = add_76070 == 32'h0000_0000 ? array_update_76923 : array_update_76912[0];
  assign array_update_76925[1] = add_76070 == 32'h0000_0001 ? array_update_76923 : array_update_76912[1];
  assign array_update_76925[2] = add_76070 == 32'h0000_0002 ? array_update_76923 : array_update_76912[2];
  assign array_update_76925[3] = add_76070 == 32'h0000_0003 ? array_update_76923 : array_update_76912[3];
  assign array_update_76925[4] = add_76070 == 32'h0000_0004 ? array_update_76923 : array_update_76912[4];
  assign array_update_76925[5] = add_76070 == 32'h0000_0005 ? array_update_76923 : array_update_76912[5];
  assign array_update_76925[6] = add_76070 == 32'h0000_0006 ? array_update_76923 : array_update_76912[6];
  assign array_update_76925[7] = add_76070 == 32'h0000_0007 ? array_update_76923 : array_update_76912[7];
  assign array_update_76925[8] = add_76070 == 32'h0000_0008 ? array_update_76923 : array_update_76912[8];
  assign array_update_76925[9] = add_76070 == 32'h0000_0009 ? array_update_76923 : array_update_76912[9];
  assign array_index_76927 = array_update_72021[add_76924 > 32'h0000_0009 ? 4'h9 : add_76924[3:0]];
  assign array_index_76928 = array_update_76925[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_76932 = smul32b_32b_x_32b(array_index_76077[add_76924 > 32'h0000_0009 ? 4'h9 : add_76924[3:0]], array_index_76927[add_76883 > 32'h0000_0009 ? 4'h9 : add_76883[3:0]]);
  assign add_76934 = array_index_76928[add_76883 > 32'h0000_0009 ? 4'h9 : add_76883[3:0]] + smul_76932;
  assign array_update_76936[0] = add_76883 == 32'h0000_0000 ? add_76934 : array_index_76928[0];
  assign array_update_76936[1] = add_76883 == 32'h0000_0001 ? add_76934 : array_index_76928[1];
  assign array_update_76936[2] = add_76883 == 32'h0000_0002 ? add_76934 : array_index_76928[2];
  assign array_update_76936[3] = add_76883 == 32'h0000_0003 ? add_76934 : array_index_76928[3];
  assign array_update_76936[4] = add_76883 == 32'h0000_0004 ? add_76934 : array_index_76928[4];
  assign array_update_76936[5] = add_76883 == 32'h0000_0005 ? add_76934 : array_index_76928[5];
  assign array_update_76936[6] = add_76883 == 32'h0000_0006 ? add_76934 : array_index_76928[6];
  assign array_update_76936[7] = add_76883 == 32'h0000_0007 ? add_76934 : array_index_76928[7];
  assign array_update_76936[8] = add_76883 == 32'h0000_0008 ? add_76934 : array_index_76928[8];
  assign array_update_76936[9] = add_76883 == 32'h0000_0009 ? add_76934 : array_index_76928[9];
  assign add_76937 = add_76924 + 32'h0000_0001;
  assign array_update_76938[0] = add_76070 == 32'h0000_0000 ? array_update_76936 : array_update_76925[0];
  assign array_update_76938[1] = add_76070 == 32'h0000_0001 ? array_update_76936 : array_update_76925[1];
  assign array_update_76938[2] = add_76070 == 32'h0000_0002 ? array_update_76936 : array_update_76925[2];
  assign array_update_76938[3] = add_76070 == 32'h0000_0003 ? array_update_76936 : array_update_76925[3];
  assign array_update_76938[4] = add_76070 == 32'h0000_0004 ? array_update_76936 : array_update_76925[4];
  assign array_update_76938[5] = add_76070 == 32'h0000_0005 ? array_update_76936 : array_update_76925[5];
  assign array_update_76938[6] = add_76070 == 32'h0000_0006 ? array_update_76936 : array_update_76925[6];
  assign array_update_76938[7] = add_76070 == 32'h0000_0007 ? array_update_76936 : array_update_76925[7];
  assign array_update_76938[8] = add_76070 == 32'h0000_0008 ? array_update_76936 : array_update_76925[8];
  assign array_update_76938[9] = add_76070 == 32'h0000_0009 ? array_update_76936 : array_update_76925[9];
  assign array_index_76940 = array_update_72021[add_76937 > 32'h0000_0009 ? 4'h9 : add_76937[3:0]];
  assign array_index_76941 = array_update_76938[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_76945 = smul32b_32b_x_32b(array_index_76077[add_76937 > 32'h0000_0009 ? 4'h9 : add_76937[3:0]], array_index_76940[add_76883 > 32'h0000_0009 ? 4'h9 : add_76883[3:0]]);
  assign add_76947 = array_index_76941[add_76883 > 32'h0000_0009 ? 4'h9 : add_76883[3:0]] + smul_76945;
  assign array_update_76949[0] = add_76883 == 32'h0000_0000 ? add_76947 : array_index_76941[0];
  assign array_update_76949[1] = add_76883 == 32'h0000_0001 ? add_76947 : array_index_76941[1];
  assign array_update_76949[2] = add_76883 == 32'h0000_0002 ? add_76947 : array_index_76941[2];
  assign array_update_76949[3] = add_76883 == 32'h0000_0003 ? add_76947 : array_index_76941[3];
  assign array_update_76949[4] = add_76883 == 32'h0000_0004 ? add_76947 : array_index_76941[4];
  assign array_update_76949[5] = add_76883 == 32'h0000_0005 ? add_76947 : array_index_76941[5];
  assign array_update_76949[6] = add_76883 == 32'h0000_0006 ? add_76947 : array_index_76941[6];
  assign array_update_76949[7] = add_76883 == 32'h0000_0007 ? add_76947 : array_index_76941[7];
  assign array_update_76949[8] = add_76883 == 32'h0000_0008 ? add_76947 : array_index_76941[8];
  assign array_update_76949[9] = add_76883 == 32'h0000_0009 ? add_76947 : array_index_76941[9];
  assign add_76950 = add_76937 + 32'h0000_0001;
  assign array_update_76951[0] = add_76070 == 32'h0000_0000 ? array_update_76949 : array_update_76938[0];
  assign array_update_76951[1] = add_76070 == 32'h0000_0001 ? array_update_76949 : array_update_76938[1];
  assign array_update_76951[2] = add_76070 == 32'h0000_0002 ? array_update_76949 : array_update_76938[2];
  assign array_update_76951[3] = add_76070 == 32'h0000_0003 ? array_update_76949 : array_update_76938[3];
  assign array_update_76951[4] = add_76070 == 32'h0000_0004 ? array_update_76949 : array_update_76938[4];
  assign array_update_76951[5] = add_76070 == 32'h0000_0005 ? array_update_76949 : array_update_76938[5];
  assign array_update_76951[6] = add_76070 == 32'h0000_0006 ? array_update_76949 : array_update_76938[6];
  assign array_update_76951[7] = add_76070 == 32'h0000_0007 ? array_update_76949 : array_update_76938[7];
  assign array_update_76951[8] = add_76070 == 32'h0000_0008 ? array_update_76949 : array_update_76938[8];
  assign array_update_76951[9] = add_76070 == 32'h0000_0009 ? array_update_76949 : array_update_76938[9];
  assign array_index_76953 = array_update_72021[add_76950 > 32'h0000_0009 ? 4'h9 : add_76950[3:0]];
  assign array_index_76954 = array_update_76951[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_76958 = smul32b_32b_x_32b(array_index_76077[add_76950 > 32'h0000_0009 ? 4'h9 : add_76950[3:0]], array_index_76953[add_76883 > 32'h0000_0009 ? 4'h9 : add_76883[3:0]]);
  assign add_76960 = array_index_76954[add_76883 > 32'h0000_0009 ? 4'h9 : add_76883[3:0]] + smul_76958;
  assign array_update_76962[0] = add_76883 == 32'h0000_0000 ? add_76960 : array_index_76954[0];
  assign array_update_76962[1] = add_76883 == 32'h0000_0001 ? add_76960 : array_index_76954[1];
  assign array_update_76962[2] = add_76883 == 32'h0000_0002 ? add_76960 : array_index_76954[2];
  assign array_update_76962[3] = add_76883 == 32'h0000_0003 ? add_76960 : array_index_76954[3];
  assign array_update_76962[4] = add_76883 == 32'h0000_0004 ? add_76960 : array_index_76954[4];
  assign array_update_76962[5] = add_76883 == 32'h0000_0005 ? add_76960 : array_index_76954[5];
  assign array_update_76962[6] = add_76883 == 32'h0000_0006 ? add_76960 : array_index_76954[6];
  assign array_update_76962[7] = add_76883 == 32'h0000_0007 ? add_76960 : array_index_76954[7];
  assign array_update_76962[8] = add_76883 == 32'h0000_0008 ? add_76960 : array_index_76954[8];
  assign array_update_76962[9] = add_76883 == 32'h0000_0009 ? add_76960 : array_index_76954[9];
  assign add_76963 = add_76950 + 32'h0000_0001;
  assign array_update_76964[0] = add_76070 == 32'h0000_0000 ? array_update_76962 : array_update_76951[0];
  assign array_update_76964[1] = add_76070 == 32'h0000_0001 ? array_update_76962 : array_update_76951[1];
  assign array_update_76964[2] = add_76070 == 32'h0000_0002 ? array_update_76962 : array_update_76951[2];
  assign array_update_76964[3] = add_76070 == 32'h0000_0003 ? array_update_76962 : array_update_76951[3];
  assign array_update_76964[4] = add_76070 == 32'h0000_0004 ? array_update_76962 : array_update_76951[4];
  assign array_update_76964[5] = add_76070 == 32'h0000_0005 ? array_update_76962 : array_update_76951[5];
  assign array_update_76964[6] = add_76070 == 32'h0000_0006 ? array_update_76962 : array_update_76951[6];
  assign array_update_76964[7] = add_76070 == 32'h0000_0007 ? array_update_76962 : array_update_76951[7];
  assign array_update_76964[8] = add_76070 == 32'h0000_0008 ? array_update_76962 : array_update_76951[8];
  assign array_update_76964[9] = add_76070 == 32'h0000_0009 ? array_update_76962 : array_update_76951[9];
  assign array_index_76966 = array_update_72021[add_76963 > 32'h0000_0009 ? 4'h9 : add_76963[3:0]];
  assign array_index_76967 = array_update_76964[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_76971 = smul32b_32b_x_32b(array_index_76077[add_76963 > 32'h0000_0009 ? 4'h9 : add_76963[3:0]], array_index_76966[add_76883 > 32'h0000_0009 ? 4'h9 : add_76883[3:0]]);
  assign add_76973 = array_index_76967[add_76883 > 32'h0000_0009 ? 4'h9 : add_76883[3:0]] + smul_76971;
  assign array_update_76975[0] = add_76883 == 32'h0000_0000 ? add_76973 : array_index_76967[0];
  assign array_update_76975[1] = add_76883 == 32'h0000_0001 ? add_76973 : array_index_76967[1];
  assign array_update_76975[2] = add_76883 == 32'h0000_0002 ? add_76973 : array_index_76967[2];
  assign array_update_76975[3] = add_76883 == 32'h0000_0003 ? add_76973 : array_index_76967[3];
  assign array_update_76975[4] = add_76883 == 32'h0000_0004 ? add_76973 : array_index_76967[4];
  assign array_update_76975[5] = add_76883 == 32'h0000_0005 ? add_76973 : array_index_76967[5];
  assign array_update_76975[6] = add_76883 == 32'h0000_0006 ? add_76973 : array_index_76967[6];
  assign array_update_76975[7] = add_76883 == 32'h0000_0007 ? add_76973 : array_index_76967[7];
  assign array_update_76975[8] = add_76883 == 32'h0000_0008 ? add_76973 : array_index_76967[8];
  assign array_update_76975[9] = add_76883 == 32'h0000_0009 ? add_76973 : array_index_76967[9];
  assign add_76976 = add_76963 + 32'h0000_0001;
  assign array_update_76977[0] = add_76070 == 32'h0000_0000 ? array_update_76975 : array_update_76964[0];
  assign array_update_76977[1] = add_76070 == 32'h0000_0001 ? array_update_76975 : array_update_76964[1];
  assign array_update_76977[2] = add_76070 == 32'h0000_0002 ? array_update_76975 : array_update_76964[2];
  assign array_update_76977[3] = add_76070 == 32'h0000_0003 ? array_update_76975 : array_update_76964[3];
  assign array_update_76977[4] = add_76070 == 32'h0000_0004 ? array_update_76975 : array_update_76964[4];
  assign array_update_76977[5] = add_76070 == 32'h0000_0005 ? array_update_76975 : array_update_76964[5];
  assign array_update_76977[6] = add_76070 == 32'h0000_0006 ? array_update_76975 : array_update_76964[6];
  assign array_update_76977[7] = add_76070 == 32'h0000_0007 ? array_update_76975 : array_update_76964[7];
  assign array_update_76977[8] = add_76070 == 32'h0000_0008 ? array_update_76975 : array_update_76964[8];
  assign array_update_76977[9] = add_76070 == 32'h0000_0009 ? array_update_76975 : array_update_76964[9];
  assign array_index_76979 = array_update_72021[add_76976 > 32'h0000_0009 ? 4'h9 : add_76976[3:0]];
  assign array_index_76980 = array_update_76977[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_76984 = smul32b_32b_x_32b(array_index_76077[add_76976 > 32'h0000_0009 ? 4'h9 : add_76976[3:0]], array_index_76979[add_76883 > 32'h0000_0009 ? 4'h9 : add_76883[3:0]]);
  assign add_76986 = array_index_76980[add_76883 > 32'h0000_0009 ? 4'h9 : add_76883[3:0]] + smul_76984;
  assign array_update_76988[0] = add_76883 == 32'h0000_0000 ? add_76986 : array_index_76980[0];
  assign array_update_76988[1] = add_76883 == 32'h0000_0001 ? add_76986 : array_index_76980[1];
  assign array_update_76988[2] = add_76883 == 32'h0000_0002 ? add_76986 : array_index_76980[2];
  assign array_update_76988[3] = add_76883 == 32'h0000_0003 ? add_76986 : array_index_76980[3];
  assign array_update_76988[4] = add_76883 == 32'h0000_0004 ? add_76986 : array_index_76980[4];
  assign array_update_76988[5] = add_76883 == 32'h0000_0005 ? add_76986 : array_index_76980[5];
  assign array_update_76988[6] = add_76883 == 32'h0000_0006 ? add_76986 : array_index_76980[6];
  assign array_update_76988[7] = add_76883 == 32'h0000_0007 ? add_76986 : array_index_76980[7];
  assign array_update_76988[8] = add_76883 == 32'h0000_0008 ? add_76986 : array_index_76980[8];
  assign array_update_76988[9] = add_76883 == 32'h0000_0009 ? add_76986 : array_index_76980[9];
  assign add_76989 = add_76976 + 32'h0000_0001;
  assign array_update_76990[0] = add_76070 == 32'h0000_0000 ? array_update_76988 : array_update_76977[0];
  assign array_update_76990[1] = add_76070 == 32'h0000_0001 ? array_update_76988 : array_update_76977[1];
  assign array_update_76990[2] = add_76070 == 32'h0000_0002 ? array_update_76988 : array_update_76977[2];
  assign array_update_76990[3] = add_76070 == 32'h0000_0003 ? array_update_76988 : array_update_76977[3];
  assign array_update_76990[4] = add_76070 == 32'h0000_0004 ? array_update_76988 : array_update_76977[4];
  assign array_update_76990[5] = add_76070 == 32'h0000_0005 ? array_update_76988 : array_update_76977[5];
  assign array_update_76990[6] = add_76070 == 32'h0000_0006 ? array_update_76988 : array_update_76977[6];
  assign array_update_76990[7] = add_76070 == 32'h0000_0007 ? array_update_76988 : array_update_76977[7];
  assign array_update_76990[8] = add_76070 == 32'h0000_0008 ? array_update_76988 : array_update_76977[8];
  assign array_update_76990[9] = add_76070 == 32'h0000_0009 ? array_update_76988 : array_update_76977[9];
  assign array_index_76992 = array_update_72021[add_76989 > 32'h0000_0009 ? 4'h9 : add_76989[3:0]];
  assign array_index_76993 = array_update_76990[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_76997 = smul32b_32b_x_32b(array_index_76077[add_76989 > 32'h0000_0009 ? 4'h9 : add_76989[3:0]], array_index_76992[add_76883 > 32'h0000_0009 ? 4'h9 : add_76883[3:0]]);
  assign add_76999 = array_index_76993[add_76883 > 32'h0000_0009 ? 4'h9 : add_76883[3:0]] + smul_76997;
  assign array_update_77001[0] = add_76883 == 32'h0000_0000 ? add_76999 : array_index_76993[0];
  assign array_update_77001[1] = add_76883 == 32'h0000_0001 ? add_76999 : array_index_76993[1];
  assign array_update_77001[2] = add_76883 == 32'h0000_0002 ? add_76999 : array_index_76993[2];
  assign array_update_77001[3] = add_76883 == 32'h0000_0003 ? add_76999 : array_index_76993[3];
  assign array_update_77001[4] = add_76883 == 32'h0000_0004 ? add_76999 : array_index_76993[4];
  assign array_update_77001[5] = add_76883 == 32'h0000_0005 ? add_76999 : array_index_76993[5];
  assign array_update_77001[6] = add_76883 == 32'h0000_0006 ? add_76999 : array_index_76993[6];
  assign array_update_77001[7] = add_76883 == 32'h0000_0007 ? add_76999 : array_index_76993[7];
  assign array_update_77001[8] = add_76883 == 32'h0000_0008 ? add_76999 : array_index_76993[8];
  assign array_update_77001[9] = add_76883 == 32'h0000_0009 ? add_76999 : array_index_76993[9];
  assign add_77002 = add_76989 + 32'h0000_0001;
  assign array_update_77003[0] = add_76070 == 32'h0000_0000 ? array_update_77001 : array_update_76990[0];
  assign array_update_77003[1] = add_76070 == 32'h0000_0001 ? array_update_77001 : array_update_76990[1];
  assign array_update_77003[2] = add_76070 == 32'h0000_0002 ? array_update_77001 : array_update_76990[2];
  assign array_update_77003[3] = add_76070 == 32'h0000_0003 ? array_update_77001 : array_update_76990[3];
  assign array_update_77003[4] = add_76070 == 32'h0000_0004 ? array_update_77001 : array_update_76990[4];
  assign array_update_77003[5] = add_76070 == 32'h0000_0005 ? array_update_77001 : array_update_76990[5];
  assign array_update_77003[6] = add_76070 == 32'h0000_0006 ? array_update_77001 : array_update_76990[6];
  assign array_update_77003[7] = add_76070 == 32'h0000_0007 ? array_update_77001 : array_update_76990[7];
  assign array_update_77003[8] = add_76070 == 32'h0000_0008 ? array_update_77001 : array_update_76990[8];
  assign array_update_77003[9] = add_76070 == 32'h0000_0009 ? array_update_77001 : array_update_76990[9];
  assign array_index_77005 = array_update_72021[add_77002 > 32'h0000_0009 ? 4'h9 : add_77002[3:0]];
  assign array_index_77006 = array_update_77003[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_77010 = smul32b_32b_x_32b(array_index_76077[add_77002 > 32'h0000_0009 ? 4'h9 : add_77002[3:0]], array_index_77005[add_76883 > 32'h0000_0009 ? 4'h9 : add_76883[3:0]]);
  assign add_77012 = array_index_77006[add_76883 > 32'h0000_0009 ? 4'h9 : add_76883[3:0]] + smul_77010;
  assign array_update_77013[0] = add_76883 == 32'h0000_0000 ? add_77012 : array_index_77006[0];
  assign array_update_77013[1] = add_76883 == 32'h0000_0001 ? add_77012 : array_index_77006[1];
  assign array_update_77013[2] = add_76883 == 32'h0000_0002 ? add_77012 : array_index_77006[2];
  assign array_update_77013[3] = add_76883 == 32'h0000_0003 ? add_77012 : array_index_77006[3];
  assign array_update_77013[4] = add_76883 == 32'h0000_0004 ? add_77012 : array_index_77006[4];
  assign array_update_77013[5] = add_76883 == 32'h0000_0005 ? add_77012 : array_index_77006[5];
  assign array_update_77013[6] = add_76883 == 32'h0000_0006 ? add_77012 : array_index_77006[6];
  assign array_update_77013[7] = add_76883 == 32'h0000_0007 ? add_77012 : array_index_77006[7];
  assign array_update_77013[8] = add_76883 == 32'h0000_0008 ? add_77012 : array_index_77006[8];
  assign array_update_77013[9] = add_76883 == 32'h0000_0009 ? add_77012 : array_index_77006[9];
  assign array_update_77014[0] = add_76070 == 32'h0000_0000 ? array_update_77013 : array_update_77003[0];
  assign array_update_77014[1] = add_76070 == 32'h0000_0001 ? array_update_77013 : array_update_77003[1];
  assign array_update_77014[2] = add_76070 == 32'h0000_0002 ? array_update_77013 : array_update_77003[2];
  assign array_update_77014[3] = add_76070 == 32'h0000_0003 ? array_update_77013 : array_update_77003[3];
  assign array_update_77014[4] = add_76070 == 32'h0000_0004 ? array_update_77013 : array_update_77003[4];
  assign array_update_77014[5] = add_76070 == 32'h0000_0005 ? array_update_77013 : array_update_77003[5];
  assign array_update_77014[6] = add_76070 == 32'h0000_0006 ? array_update_77013 : array_update_77003[6];
  assign array_update_77014[7] = add_76070 == 32'h0000_0007 ? array_update_77013 : array_update_77003[7];
  assign array_update_77014[8] = add_76070 == 32'h0000_0008 ? array_update_77013 : array_update_77003[8];
  assign array_update_77014[9] = add_76070 == 32'h0000_0009 ? array_update_77013 : array_update_77003[9];
  assign array_index_77016 = array_update_77014[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign add_77018 = add_76883 + 32'h0000_0001;
  assign array_update_77019[0] = add_77018 == 32'h0000_0000 ? 32'h0000_0000 : array_index_77016[0];
  assign array_update_77019[1] = add_77018 == 32'h0000_0001 ? 32'h0000_0000 : array_index_77016[1];
  assign array_update_77019[2] = add_77018 == 32'h0000_0002 ? 32'h0000_0000 : array_index_77016[2];
  assign array_update_77019[3] = add_77018 == 32'h0000_0003 ? 32'h0000_0000 : array_index_77016[3];
  assign array_update_77019[4] = add_77018 == 32'h0000_0004 ? 32'h0000_0000 : array_index_77016[4];
  assign array_update_77019[5] = add_77018 == 32'h0000_0005 ? 32'h0000_0000 : array_index_77016[5];
  assign array_update_77019[6] = add_77018 == 32'h0000_0006 ? 32'h0000_0000 : array_index_77016[6];
  assign array_update_77019[7] = add_77018 == 32'h0000_0007 ? 32'h0000_0000 : array_index_77016[7];
  assign array_update_77019[8] = add_77018 == 32'h0000_0008 ? 32'h0000_0000 : array_index_77016[8];
  assign array_update_77019[9] = add_77018 == 32'h0000_0009 ? 32'h0000_0000 : array_index_77016[9];
  assign literal_77020 = 32'h0000_0000;
  assign array_update_77021[0] = add_76070 == 32'h0000_0000 ? array_update_77019 : array_update_77014[0];
  assign array_update_77021[1] = add_76070 == 32'h0000_0001 ? array_update_77019 : array_update_77014[1];
  assign array_update_77021[2] = add_76070 == 32'h0000_0002 ? array_update_77019 : array_update_77014[2];
  assign array_update_77021[3] = add_76070 == 32'h0000_0003 ? array_update_77019 : array_update_77014[3];
  assign array_update_77021[4] = add_76070 == 32'h0000_0004 ? array_update_77019 : array_update_77014[4];
  assign array_update_77021[5] = add_76070 == 32'h0000_0005 ? array_update_77019 : array_update_77014[5];
  assign array_update_77021[6] = add_76070 == 32'h0000_0006 ? array_update_77019 : array_update_77014[6];
  assign array_update_77021[7] = add_76070 == 32'h0000_0007 ? array_update_77019 : array_update_77014[7];
  assign array_update_77021[8] = add_76070 == 32'h0000_0008 ? array_update_77019 : array_update_77014[8];
  assign array_update_77021[9] = add_76070 == 32'h0000_0009 ? array_update_77019 : array_update_77014[9];
  assign array_index_77023 = array_update_72021[literal_77020 > 32'h0000_0009 ? 4'h9 : literal_77020[3:0]];
  assign array_index_77024 = array_update_77021[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_77028 = smul32b_32b_x_32b(array_index_76077[literal_77020 > 32'h0000_0009 ? 4'h9 : literal_77020[3:0]], array_index_77023[add_77018 > 32'h0000_0009 ? 4'h9 : add_77018[3:0]]);
  assign add_77030 = array_index_77024[add_77018 > 32'h0000_0009 ? 4'h9 : add_77018[3:0]] + smul_77028;
  assign array_update_77032[0] = add_77018 == 32'h0000_0000 ? add_77030 : array_index_77024[0];
  assign array_update_77032[1] = add_77018 == 32'h0000_0001 ? add_77030 : array_index_77024[1];
  assign array_update_77032[2] = add_77018 == 32'h0000_0002 ? add_77030 : array_index_77024[2];
  assign array_update_77032[3] = add_77018 == 32'h0000_0003 ? add_77030 : array_index_77024[3];
  assign array_update_77032[4] = add_77018 == 32'h0000_0004 ? add_77030 : array_index_77024[4];
  assign array_update_77032[5] = add_77018 == 32'h0000_0005 ? add_77030 : array_index_77024[5];
  assign array_update_77032[6] = add_77018 == 32'h0000_0006 ? add_77030 : array_index_77024[6];
  assign array_update_77032[7] = add_77018 == 32'h0000_0007 ? add_77030 : array_index_77024[7];
  assign array_update_77032[8] = add_77018 == 32'h0000_0008 ? add_77030 : array_index_77024[8];
  assign array_update_77032[9] = add_77018 == 32'h0000_0009 ? add_77030 : array_index_77024[9];
  assign add_77033 = literal_77020 + 32'h0000_0001;
  assign array_update_77034[0] = add_76070 == 32'h0000_0000 ? array_update_77032 : array_update_77021[0];
  assign array_update_77034[1] = add_76070 == 32'h0000_0001 ? array_update_77032 : array_update_77021[1];
  assign array_update_77034[2] = add_76070 == 32'h0000_0002 ? array_update_77032 : array_update_77021[2];
  assign array_update_77034[3] = add_76070 == 32'h0000_0003 ? array_update_77032 : array_update_77021[3];
  assign array_update_77034[4] = add_76070 == 32'h0000_0004 ? array_update_77032 : array_update_77021[4];
  assign array_update_77034[5] = add_76070 == 32'h0000_0005 ? array_update_77032 : array_update_77021[5];
  assign array_update_77034[6] = add_76070 == 32'h0000_0006 ? array_update_77032 : array_update_77021[6];
  assign array_update_77034[7] = add_76070 == 32'h0000_0007 ? array_update_77032 : array_update_77021[7];
  assign array_update_77034[8] = add_76070 == 32'h0000_0008 ? array_update_77032 : array_update_77021[8];
  assign array_update_77034[9] = add_76070 == 32'h0000_0009 ? array_update_77032 : array_update_77021[9];
  assign array_index_77036 = array_update_72021[add_77033 > 32'h0000_0009 ? 4'h9 : add_77033[3:0]];
  assign array_index_77037 = array_update_77034[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_77041 = smul32b_32b_x_32b(array_index_76077[add_77033 > 32'h0000_0009 ? 4'h9 : add_77033[3:0]], array_index_77036[add_77018 > 32'h0000_0009 ? 4'h9 : add_77018[3:0]]);
  assign add_77043 = array_index_77037[add_77018 > 32'h0000_0009 ? 4'h9 : add_77018[3:0]] + smul_77041;
  assign array_update_77045[0] = add_77018 == 32'h0000_0000 ? add_77043 : array_index_77037[0];
  assign array_update_77045[1] = add_77018 == 32'h0000_0001 ? add_77043 : array_index_77037[1];
  assign array_update_77045[2] = add_77018 == 32'h0000_0002 ? add_77043 : array_index_77037[2];
  assign array_update_77045[3] = add_77018 == 32'h0000_0003 ? add_77043 : array_index_77037[3];
  assign array_update_77045[4] = add_77018 == 32'h0000_0004 ? add_77043 : array_index_77037[4];
  assign array_update_77045[5] = add_77018 == 32'h0000_0005 ? add_77043 : array_index_77037[5];
  assign array_update_77045[6] = add_77018 == 32'h0000_0006 ? add_77043 : array_index_77037[6];
  assign array_update_77045[7] = add_77018 == 32'h0000_0007 ? add_77043 : array_index_77037[7];
  assign array_update_77045[8] = add_77018 == 32'h0000_0008 ? add_77043 : array_index_77037[8];
  assign array_update_77045[9] = add_77018 == 32'h0000_0009 ? add_77043 : array_index_77037[9];
  assign add_77046 = add_77033 + 32'h0000_0001;
  assign array_update_77047[0] = add_76070 == 32'h0000_0000 ? array_update_77045 : array_update_77034[0];
  assign array_update_77047[1] = add_76070 == 32'h0000_0001 ? array_update_77045 : array_update_77034[1];
  assign array_update_77047[2] = add_76070 == 32'h0000_0002 ? array_update_77045 : array_update_77034[2];
  assign array_update_77047[3] = add_76070 == 32'h0000_0003 ? array_update_77045 : array_update_77034[3];
  assign array_update_77047[4] = add_76070 == 32'h0000_0004 ? array_update_77045 : array_update_77034[4];
  assign array_update_77047[5] = add_76070 == 32'h0000_0005 ? array_update_77045 : array_update_77034[5];
  assign array_update_77047[6] = add_76070 == 32'h0000_0006 ? array_update_77045 : array_update_77034[6];
  assign array_update_77047[7] = add_76070 == 32'h0000_0007 ? array_update_77045 : array_update_77034[7];
  assign array_update_77047[8] = add_76070 == 32'h0000_0008 ? array_update_77045 : array_update_77034[8];
  assign array_update_77047[9] = add_76070 == 32'h0000_0009 ? array_update_77045 : array_update_77034[9];
  assign array_index_77049 = array_update_72021[add_77046 > 32'h0000_0009 ? 4'h9 : add_77046[3:0]];
  assign array_index_77050 = array_update_77047[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_77054 = smul32b_32b_x_32b(array_index_76077[add_77046 > 32'h0000_0009 ? 4'h9 : add_77046[3:0]], array_index_77049[add_77018 > 32'h0000_0009 ? 4'h9 : add_77018[3:0]]);
  assign add_77056 = array_index_77050[add_77018 > 32'h0000_0009 ? 4'h9 : add_77018[3:0]] + smul_77054;
  assign array_update_77058[0] = add_77018 == 32'h0000_0000 ? add_77056 : array_index_77050[0];
  assign array_update_77058[1] = add_77018 == 32'h0000_0001 ? add_77056 : array_index_77050[1];
  assign array_update_77058[2] = add_77018 == 32'h0000_0002 ? add_77056 : array_index_77050[2];
  assign array_update_77058[3] = add_77018 == 32'h0000_0003 ? add_77056 : array_index_77050[3];
  assign array_update_77058[4] = add_77018 == 32'h0000_0004 ? add_77056 : array_index_77050[4];
  assign array_update_77058[5] = add_77018 == 32'h0000_0005 ? add_77056 : array_index_77050[5];
  assign array_update_77058[6] = add_77018 == 32'h0000_0006 ? add_77056 : array_index_77050[6];
  assign array_update_77058[7] = add_77018 == 32'h0000_0007 ? add_77056 : array_index_77050[7];
  assign array_update_77058[8] = add_77018 == 32'h0000_0008 ? add_77056 : array_index_77050[8];
  assign array_update_77058[9] = add_77018 == 32'h0000_0009 ? add_77056 : array_index_77050[9];
  assign add_77059 = add_77046 + 32'h0000_0001;
  assign array_update_77060[0] = add_76070 == 32'h0000_0000 ? array_update_77058 : array_update_77047[0];
  assign array_update_77060[1] = add_76070 == 32'h0000_0001 ? array_update_77058 : array_update_77047[1];
  assign array_update_77060[2] = add_76070 == 32'h0000_0002 ? array_update_77058 : array_update_77047[2];
  assign array_update_77060[3] = add_76070 == 32'h0000_0003 ? array_update_77058 : array_update_77047[3];
  assign array_update_77060[4] = add_76070 == 32'h0000_0004 ? array_update_77058 : array_update_77047[4];
  assign array_update_77060[5] = add_76070 == 32'h0000_0005 ? array_update_77058 : array_update_77047[5];
  assign array_update_77060[6] = add_76070 == 32'h0000_0006 ? array_update_77058 : array_update_77047[6];
  assign array_update_77060[7] = add_76070 == 32'h0000_0007 ? array_update_77058 : array_update_77047[7];
  assign array_update_77060[8] = add_76070 == 32'h0000_0008 ? array_update_77058 : array_update_77047[8];
  assign array_update_77060[9] = add_76070 == 32'h0000_0009 ? array_update_77058 : array_update_77047[9];
  assign array_index_77062 = array_update_72021[add_77059 > 32'h0000_0009 ? 4'h9 : add_77059[3:0]];
  assign array_index_77063 = array_update_77060[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_77067 = smul32b_32b_x_32b(array_index_76077[add_77059 > 32'h0000_0009 ? 4'h9 : add_77059[3:0]], array_index_77062[add_77018 > 32'h0000_0009 ? 4'h9 : add_77018[3:0]]);
  assign add_77069 = array_index_77063[add_77018 > 32'h0000_0009 ? 4'h9 : add_77018[3:0]] + smul_77067;
  assign array_update_77071[0] = add_77018 == 32'h0000_0000 ? add_77069 : array_index_77063[0];
  assign array_update_77071[1] = add_77018 == 32'h0000_0001 ? add_77069 : array_index_77063[1];
  assign array_update_77071[2] = add_77018 == 32'h0000_0002 ? add_77069 : array_index_77063[2];
  assign array_update_77071[3] = add_77018 == 32'h0000_0003 ? add_77069 : array_index_77063[3];
  assign array_update_77071[4] = add_77018 == 32'h0000_0004 ? add_77069 : array_index_77063[4];
  assign array_update_77071[5] = add_77018 == 32'h0000_0005 ? add_77069 : array_index_77063[5];
  assign array_update_77071[6] = add_77018 == 32'h0000_0006 ? add_77069 : array_index_77063[6];
  assign array_update_77071[7] = add_77018 == 32'h0000_0007 ? add_77069 : array_index_77063[7];
  assign array_update_77071[8] = add_77018 == 32'h0000_0008 ? add_77069 : array_index_77063[8];
  assign array_update_77071[9] = add_77018 == 32'h0000_0009 ? add_77069 : array_index_77063[9];
  assign add_77072 = add_77059 + 32'h0000_0001;
  assign array_update_77073[0] = add_76070 == 32'h0000_0000 ? array_update_77071 : array_update_77060[0];
  assign array_update_77073[1] = add_76070 == 32'h0000_0001 ? array_update_77071 : array_update_77060[1];
  assign array_update_77073[2] = add_76070 == 32'h0000_0002 ? array_update_77071 : array_update_77060[2];
  assign array_update_77073[3] = add_76070 == 32'h0000_0003 ? array_update_77071 : array_update_77060[3];
  assign array_update_77073[4] = add_76070 == 32'h0000_0004 ? array_update_77071 : array_update_77060[4];
  assign array_update_77073[5] = add_76070 == 32'h0000_0005 ? array_update_77071 : array_update_77060[5];
  assign array_update_77073[6] = add_76070 == 32'h0000_0006 ? array_update_77071 : array_update_77060[6];
  assign array_update_77073[7] = add_76070 == 32'h0000_0007 ? array_update_77071 : array_update_77060[7];
  assign array_update_77073[8] = add_76070 == 32'h0000_0008 ? array_update_77071 : array_update_77060[8];
  assign array_update_77073[9] = add_76070 == 32'h0000_0009 ? array_update_77071 : array_update_77060[9];
  assign array_index_77075 = array_update_72021[add_77072 > 32'h0000_0009 ? 4'h9 : add_77072[3:0]];
  assign array_index_77076 = array_update_77073[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_77080 = smul32b_32b_x_32b(array_index_76077[add_77072 > 32'h0000_0009 ? 4'h9 : add_77072[3:0]], array_index_77075[add_77018 > 32'h0000_0009 ? 4'h9 : add_77018[3:0]]);
  assign add_77082 = array_index_77076[add_77018 > 32'h0000_0009 ? 4'h9 : add_77018[3:0]] + smul_77080;
  assign array_update_77084[0] = add_77018 == 32'h0000_0000 ? add_77082 : array_index_77076[0];
  assign array_update_77084[1] = add_77018 == 32'h0000_0001 ? add_77082 : array_index_77076[1];
  assign array_update_77084[2] = add_77018 == 32'h0000_0002 ? add_77082 : array_index_77076[2];
  assign array_update_77084[3] = add_77018 == 32'h0000_0003 ? add_77082 : array_index_77076[3];
  assign array_update_77084[4] = add_77018 == 32'h0000_0004 ? add_77082 : array_index_77076[4];
  assign array_update_77084[5] = add_77018 == 32'h0000_0005 ? add_77082 : array_index_77076[5];
  assign array_update_77084[6] = add_77018 == 32'h0000_0006 ? add_77082 : array_index_77076[6];
  assign array_update_77084[7] = add_77018 == 32'h0000_0007 ? add_77082 : array_index_77076[7];
  assign array_update_77084[8] = add_77018 == 32'h0000_0008 ? add_77082 : array_index_77076[8];
  assign array_update_77084[9] = add_77018 == 32'h0000_0009 ? add_77082 : array_index_77076[9];
  assign add_77085 = add_77072 + 32'h0000_0001;
  assign array_update_77086[0] = add_76070 == 32'h0000_0000 ? array_update_77084 : array_update_77073[0];
  assign array_update_77086[1] = add_76070 == 32'h0000_0001 ? array_update_77084 : array_update_77073[1];
  assign array_update_77086[2] = add_76070 == 32'h0000_0002 ? array_update_77084 : array_update_77073[2];
  assign array_update_77086[3] = add_76070 == 32'h0000_0003 ? array_update_77084 : array_update_77073[3];
  assign array_update_77086[4] = add_76070 == 32'h0000_0004 ? array_update_77084 : array_update_77073[4];
  assign array_update_77086[5] = add_76070 == 32'h0000_0005 ? array_update_77084 : array_update_77073[5];
  assign array_update_77086[6] = add_76070 == 32'h0000_0006 ? array_update_77084 : array_update_77073[6];
  assign array_update_77086[7] = add_76070 == 32'h0000_0007 ? array_update_77084 : array_update_77073[7];
  assign array_update_77086[8] = add_76070 == 32'h0000_0008 ? array_update_77084 : array_update_77073[8];
  assign array_update_77086[9] = add_76070 == 32'h0000_0009 ? array_update_77084 : array_update_77073[9];
  assign array_index_77088 = array_update_72021[add_77085 > 32'h0000_0009 ? 4'h9 : add_77085[3:0]];
  assign array_index_77089 = array_update_77086[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_77093 = smul32b_32b_x_32b(array_index_76077[add_77085 > 32'h0000_0009 ? 4'h9 : add_77085[3:0]], array_index_77088[add_77018 > 32'h0000_0009 ? 4'h9 : add_77018[3:0]]);
  assign add_77095 = array_index_77089[add_77018 > 32'h0000_0009 ? 4'h9 : add_77018[3:0]] + smul_77093;
  assign array_update_77097[0] = add_77018 == 32'h0000_0000 ? add_77095 : array_index_77089[0];
  assign array_update_77097[1] = add_77018 == 32'h0000_0001 ? add_77095 : array_index_77089[1];
  assign array_update_77097[2] = add_77018 == 32'h0000_0002 ? add_77095 : array_index_77089[2];
  assign array_update_77097[3] = add_77018 == 32'h0000_0003 ? add_77095 : array_index_77089[3];
  assign array_update_77097[4] = add_77018 == 32'h0000_0004 ? add_77095 : array_index_77089[4];
  assign array_update_77097[5] = add_77018 == 32'h0000_0005 ? add_77095 : array_index_77089[5];
  assign array_update_77097[6] = add_77018 == 32'h0000_0006 ? add_77095 : array_index_77089[6];
  assign array_update_77097[7] = add_77018 == 32'h0000_0007 ? add_77095 : array_index_77089[7];
  assign array_update_77097[8] = add_77018 == 32'h0000_0008 ? add_77095 : array_index_77089[8];
  assign array_update_77097[9] = add_77018 == 32'h0000_0009 ? add_77095 : array_index_77089[9];
  assign add_77098 = add_77085 + 32'h0000_0001;
  assign array_update_77099[0] = add_76070 == 32'h0000_0000 ? array_update_77097 : array_update_77086[0];
  assign array_update_77099[1] = add_76070 == 32'h0000_0001 ? array_update_77097 : array_update_77086[1];
  assign array_update_77099[2] = add_76070 == 32'h0000_0002 ? array_update_77097 : array_update_77086[2];
  assign array_update_77099[3] = add_76070 == 32'h0000_0003 ? array_update_77097 : array_update_77086[3];
  assign array_update_77099[4] = add_76070 == 32'h0000_0004 ? array_update_77097 : array_update_77086[4];
  assign array_update_77099[5] = add_76070 == 32'h0000_0005 ? array_update_77097 : array_update_77086[5];
  assign array_update_77099[6] = add_76070 == 32'h0000_0006 ? array_update_77097 : array_update_77086[6];
  assign array_update_77099[7] = add_76070 == 32'h0000_0007 ? array_update_77097 : array_update_77086[7];
  assign array_update_77099[8] = add_76070 == 32'h0000_0008 ? array_update_77097 : array_update_77086[8];
  assign array_update_77099[9] = add_76070 == 32'h0000_0009 ? array_update_77097 : array_update_77086[9];
  assign array_index_77101 = array_update_72021[add_77098 > 32'h0000_0009 ? 4'h9 : add_77098[3:0]];
  assign array_index_77102 = array_update_77099[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_77106 = smul32b_32b_x_32b(array_index_76077[add_77098 > 32'h0000_0009 ? 4'h9 : add_77098[3:0]], array_index_77101[add_77018 > 32'h0000_0009 ? 4'h9 : add_77018[3:0]]);
  assign add_77108 = array_index_77102[add_77018 > 32'h0000_0009 ? 4'h9 : add_77018[3:0]] + smul_77106;
  assign array_update_77110[0] = add_77018 == 32'h0000_0000 ? add_77108 : array_index_77102[0];
  assign array_update_77110[1] = add_77018 == 32'h0000_0001 ? add_77108 : array_index_77102[1];
  assign array_update_77110[2] = add_77018 == 32'h0000_0002 ? add_77108 : array_index_77102[2];
  assign array_update_77110[3] = add_77018 == 32'h0000_0003 ? add_77108 : array_index_77102[3];
  assign array_update_77110[4] = add_77018 == 32'h0000_0004 ? add_77108 : array_index_77102[4];
  assign array_update_77110[5] = add_77018 == 32'h0000_0005 ? add_77108 : array_index_77102[5];
  assign array_update_77110[6] = add_77018 == 32'h0000_0006 ? add_77108 : array_index_77102[6];
  assign array_update_77110[7] = add_77018 == 32'h0000_0007 ? add_77108 : array_index_77102[7];
  assign array_update_77110[8] = add_77018 == 32'h0000_0008 ? add_77108 : array_index_77102[8];
  assign array_update_77110[9] = add_77018 == 32'h0000_0009 ? add_77108 : array_index_77102[9];
  assign add_77111 = add_77098 + 32'h0000_0001;
  assign array_update_77112[0] = add_76070 == 32'h0000_0000 ? array_update_77110 : array_update_77099[0];
  assign array_update_77112[1] = add_76070 == 32'h0000_0001 ? array_update_77110 : array_update_77099[1];
  assign array_update_77112[2] = add_76070 == 32'h0000_0002 ? array_update_77110 : array_update_77099[2];
  assign array_update_77112[3] = add_76070 == 32'h0000_0003 ? array_update_77110 : array_update_77099[3];
  assign array_update_77112[4] = add_76070 == 32'h0000_0004 ? array_update_77110 : array_update_77099[4];
  assign array_update_77112[5] = add_76070 == 32'h0000_0005 ? array_update_77110 : array_update_77099[5];
  assign array_update_77112[6] = add_76070 == 32'h0000_0006 ? array_update_77110 : array_update_77099[6];
  assign array_update_77112[7] = add_76070 == 32'h0000_0007 ? array_update_77110 : array_update_77099[7];
  assign array_update_77112[8] = add_76070 == 32'h0000_0008 ? array_update_77110 : array_update_77099[8];
  assign array_update_77112[9] = add_76070 == 32'h0000_0009 ? array_update_77110 : array_update_77099[9];
  assign array_index_77114 = array_update_72021[add_77111 > 32'h0000_0009 ? 4'h9 : add_77111[3:0]];
  assign array_index_77115 = array_update_77112[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_77119 = smul32b_32b_x_32b(array_index_76077[add_77111 > 32'h0000_0009 ? 4'h9 : add_77111[3:0]], array_index_77114[add_77018 > 32'h0000_0009 ? 4'h9 : add_77018[3:0]]);
  assign add_77121 = array_index_77115[add_77018 > 32'h0000_0009 ? 4'h9 : add_77018[3:0]] + smul_77119;
  assign array_update_77123[0] = add_77018 == 32'h0000_0000 ? add_77121 : array_index_77115[0];
  assign array_update_77123[1] = add_77018 == 32'h0000_0001 ? add_77121 : array_index_77115[1];
  assign array_update_77123[2] = add_77018 == 32'h0000_0002 ? add_77121 : array_index_77115[2];
  assign array_update_77123[3] = add_77018 == 32'h0000_0003 ? add_77121 : array_index_77115[3];
  assign array_update_77123[4] = add_77018 == 32'h0000_0004 ? add_77121 : array_index_77115[4];
  assign array_update_77123[5] = add_77018 == 32'h0000_0005 ? add_77121 : array_index_77115[5];
  assign array_update_77123[6] = add_77018 == 32'h0000_0006 ? add_77121 : array_index_77115[6];
  assign array_update_77123[7] = add_77018 == 32'h0000_0007 ? add_77121 : array_index_77115[7];
  assign array_update_77123[8] = add_77018 == 32'h0000_0008 ? add_77121 : array_index_77115[8];
  assign array_update_77123[9] = add_77018 == 32'h0000_0009 ? add_77121 : array_index_77115[9];
  assign add_77124 = add_77111 + 32'h0000_0001;
  assign array_update_77125[0] = add_76070 == 32'h0000_0000 ? array_update_77123 : array_update_77112[0];
  assign array_update_77125[1] = add_76070 == 32'h0000_0001 ? array_update_77123 : array_update_77112[1];
  assign array_update_77125[2] = add_76070 == 32'h0000_0002 ? array_update_77123 : array_update_77112[2];
  assign array_update_77125[3] = add_76070 == 32'h0000_0003 ? array_update_77123 : array_update_77112[3];
  assign array_update_77125[4] = add_76070 == 32'h0000_0004 ? array_update_77123 : array_update_77112[4];
  assign array_update_77125[5] = add_76070 == 32'h0000_0005 ? array_update_77123 : array_update_77112[5];
  assign array_update_77125[6] = add_76070 == 32'h0000_0006 ? array_update_77123 : array_update_77112[6];
  assign array_update_77125[7] = add_76070 == 32'h0000_0007 ? array_update_77123 : array_update_77112[7];
  assign array_update_77125[8] = add_76070 == 32'h0000_0008 ? array_update_77123 : array_update_77112[8];
  assign array_update_77125[9] = add_76070 == 32'h0000_0009 ? array_update_77123 : array_update_77112[9];
  assign array_index_77127 = array_update_72021[add_77124 > 32'h0000_0009 ? 4'h9 : add_77124[3:0]];
  assign array_index_77128 = array_update_77125[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_77132 = smul32b_32b_x_32b(array_index_76077[add_77124 > 32'h0000_0009 ? 4'h9 : add_77124[3:0]], array_index_77127[add_77018 > 32'h0000_0009 ? 4'h9 : add_77018[3:0]]);
  assign add_77134 = array_index_77128[add_77018 > 32'h0000_0009 ? 4'h9 : add_77018[3:0]] + smul_77132;
  assign array_update_77136[0] = add_77018 == 32'h0000_0000 ? add_77134 : array_index_77128[0];
  assign array_update_77136[1] = add_77018 == 32'h0000_0001 ? add_77134 : array_index_77128[1];
  assign array_update_77136[2] = add_77018 == 32'h0000_0002 ? add_77134 : array_index_77128[2];
  assign array_update_77136[3] = add_77018 == 32'h0000_0003 ? add_77134 : array_index_77128[3];
  assign array_update_77136[4] = add_77018 == 32'h0000_0004 ? add_77134 : array_index_77128[4];
  assign array_update_77136[5] = add_77018 == 32'h0000_0005 ? add_77134 : array_index_77128[5];
  assign array_update_77136[6] = add_77018 == 32'h0000_0006 ? add_77134 : array_index_77128[6];
  assign array_update_77136[7] = add_77018 == 32'h0000_0007 ? add_77134 : array_index_77128[7];
  assign array_update_77136[8] = add_77018 == 32'h0000_0008 ? add_77134 : array_index_77128[8];
  assign array_update_77136[9] = add_77018 == 32'h0000_0009 ? add_77134 : array_index_77128[9];
  assign add_77137 = add_77124 + 32'h0000_0001;
  assign array_update_77138[0] = add_76070 == 32'h0000_0000 ? array_update_77136 : array_update_77125[0];
  assign array_update_77138[1] = add_76070 == 32'h0000_0001 ? array_update_77136 : array_update_77125[1];
  assign array_update_77138[2] = add_76070 == 32'h0000_0002 ? array_update_77136 : array_update_77125[2];
  assign array_update_77138[3] = add_76070 == 32'h0000_0003 ? array_update_77136 : array_update_77125[3];
  assign array_update_77138[4] = add_76070 == 32'h0000_0004 ? array_update_77136 : array_update_77125[4];
  assign array_update_77138[5] = add_76070 == 32'h0000_0005 ? array_update_77136 : array_update_77125[5];
  assign array_update_77138[6] = add_76070 == 32'h0000_0006 ? array_update_77136 : array_update_77125[6];
  assign array_update_77138[7] = add_76070 == 32'h0000_0007 ? array_update_77136 : array_update_77125[7];
  assign array_update_77138[8] = add_76070 == 32'h0000_0008 ? array_update_77136 : array_update_77125[8];
  assign array_update_77138[9] = add_76070 == 32'h0000_0009 ? array_update_77136 : array_update_77125[9];
  assign array_index_77140 = array_update_72021[add_77137 > 32'h0000_0009 ? 4'h9 : add_77137[3:0]];
  assign array_index_77141 = array_update_77138[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_77145 = smul32b_32b_x_32b(array_index_76077[add_77137 > 32'h0000_0009 ? 4'h9 : add_77137[3:0]], array_index_77140[add_77018 > 32'h0000_0009 ? 4'h9 : add_77018[3:0]]);
  assign add_77147 = array_index_77141[add_77018 > 32'h0000_0009 ? 4'h9 : add_77018[3:0]] + smul_77145;
  assign array_update_77148[0] = add_77018 == 32'h0000_0000 ? add_77147 : array_index_77141[0];
  assign array_update_77148[1] = add_77018 == 32'h0000_0001 ? add_77147 : array_index_77141[1];
  assign array_update_77148[2] = add_77018 == 32'h0000_0002 ? add_77147 : array_index_77141[2];
  assign array_update_77148[3] = add_77018 == 32'h0000_0003 ? add_77147 : array_index_77141[3];
  assign array_update_77148[4] = add_77018 == 32'h0000_0004 ? add_77147 : array_index_77141[4];
  assign array_update_77148[5] = add_77018 == 32'h0000_0005 ? add_77147 : array_index_77141[5];
  assign array_update_77148[6] = add_77018 == 32'h0000_0006 ? add_77147 : array_index_77141[6];
  assign array_update_77148[7] = add_77018 == 32'h0000_0007 ? add_77147 : array_index_77141[7];
  assign array_update_77148[8] = add_77018 == 32'h0000_0008 ? add_77147 : array_index_77141[8];
  assign array_update_77148[9] = add_77018 == 32'h0000_0009 ? add_77147 : array_index_77141[9];
  assign array_update_77149[0] = add_76070 == 32'h0000_0000 ? array_update_77148 : array_update_77138[0];
  assign array_update_77149[1] = add_76070 == 32'h0000_0001 ? array_update_77148 : array_update_77138[1];
  assign array_update_77149[2] = add_76070 == 32'h0000_0002 ? array_update_77148 : array_update_77138[2];
  assign array_update_77149[3] = add_76070 == 32'h0000_0003 ? array_update_77148 : array_update_77138[3];
  assign array_update_77149[4] = add_76070 == 32'h0000_0004 ? array_update_77148 : array_update_77138[4];
  assign array_update_77149[5] = add_76070 == 32'h0000_0005 ? array_update_77148 : array_update_77138[5];
  assign array_update_77149[6] = add_76070 == 32'h0000_0006 ? array_update_77148 : array_update_77138[6];
  assign array_update_77149[7] = add_76070 == 32'h0000_0007 ? array_update_77148 : array_update_77138[7];
  assign array_update_77149[8] = add_76070 == 32'h0000_0008 ? array_update_77148 : array_update_77138[8];
  assign array_update_77149[9] = add_76070 == 32'h0000_0009 ? array_update_77148 : array_update_77138[9];
  assign array_index_77151 = array_update_77149[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign add_77153 = add_77018 + 32'h0000_0001;
  assign array_update_77154[0] = add_77153 == 32'h0000_0000 ? 32'h0000_0000 : array_index_77151[0];
  assign array_update_77154[1] = add_77153 == 32'h0000_0001 ? 32'h0000_0000 : array_index_77151[1];
  assign array_update_77154[2] = add_77153 == 32'h0000_0002 ? 32'h0000_0000 : array_index_77151[2];
  assign array_update_77154[3] = add_77153 == 32'h0000_0003 ? 32'h0000_0000 : array_index_77151[3];
  assign array_update_77154[4] = add_77153 == 32'h0000_0004 ? 32'h0000_0000 : array_index_77151[4];
  assign array_update_77154[5] = add_77153 == 32'h0000_0005 ? 32'h0000_0000 : array_index_77151[5];
  assign array_update_77154[6] = add_77153 == 32'h0000_0006 ? 32'h0000_0000 : array_index_77151[6];
  assign array_update_77154[7] = add_77153 == 32'h0000_0007 ? 32'h0000_0000 : array_index_77151[7];
  assign array_update_77154[8] = add_77153 == 32'h0000_0008 ? 32'h0000_0000 : array_index_77151[8];
  assign array_update_77154[9] = add_77153 == 32'h0000_0009 ? 32'h0000_0000 : array_index_77151[9];
  assign literal_77155 = 32'h0000_0000;
  assign array_update_77156[0] = add_76070 == 32'h0000_0000 ? array_update_77154 : array_update_77149[0];
  assign array_update_77156[1] = add_76070 == 32'h0000_0001 ? array_update_77154 : array_update_77149[1];
  assign array_update_77156[2] = add_76070 == 32'h0000_0002 ? array_update_77154 : array_update_77149[2];
  assign array_update_77156[3] = add_76070 == 32'h0000_0003 ? array_update_77154 : array_update_77149[3];
  assign array_update_77156[4] = add_76070 == 32'h0000_0004 ? array_update_77154 : array_update_77149[4];
  assign array_update_77156[5] = add_76070 == 32'h0000_0005 ? array_update_77154 : array_update_77149[5];
  assign array_update_77156[6] = add_76070 == 32'h0000_0006 ? array_update_77154 : array_update_77149[6];
  assign array_update_77156[7] = add_76070 == 32'h0000_0007 ? array_update_77154 : array_update_77149[7];
  assign array_update_77156[8] = add_76070 == 32'h0000_0008 ? array_update_77154 : array_update_77149[8];
  assign array_update_77156[9] = add_76070 == 32'h0000_0009 ? array_update_77154 : array_update_77149[9];
  assign array_index_77158 = array_update_72021[literal_77155 > 32'h0000_0009 ? 4'h9 : literal_77155[3:0]];
  assign array_index_77159 = array_update_77156[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_77163 = smul32b_32b_x_32b(array_index_76077[literal_77155 > 32'h0000_0009 ? 4'h9 : literal_77155[3:0]], array_index_77158[add_77153 > 32'h0000_0009 ? 4'h9 : add_77153[3:0]]);
  assign add_77165 = array_index_77159[add_77153 > 32'h0000_0009 ? 4'h9 : add_77153[3:0]] + smul_77163;
  assign array_update_77167[0] = add_77153 == 32'h0000_0000 ? add_77165 : array_index_77159[0];
  assign array_update_77167[1] = add_77153 == 32'h0000_0001 ? add_77165 : array_index_77159[1];
  assign array_update_77167[2] = add_77153 == 32'h0000_0002 ? add_77165 : array_index_77159[2];
  assign array_update_77167[3] = add_77153 == 32'h0000_0003 ? add_77165 : array_index_77159[3];
  assign array_update_77167[4] = add_77153 == 32'h0000_0004 ? add_77165 : array_index_77159[4];
  assign array_update_77167[5] = add_77153 == 32'h0000_0005 ? add_77165 : array_index_77159[5];
  assign array_update_77167[6] = add_77153 == 32'h0000_0006 ? add_77165 : array_index_77159[6];
  assign array_update_77167[7] = add_77153 == 32'h0000_0007 ? add_77165 : array_index_77159[7];
  assign array_update_77167[8] = add_77153 == 32'h0000_0008 ? add_77165 : array_index_77159[8];
  assign array_update_77167[9] = add_77153 == 32'h0000_0009 ? add_77165 : array_index_77159[9];
  assign add_77168 = literal_77155 + 32'h0000_0001;
  assign array_update_77169[0] = add_76070 == 32'h0000_0000 ? array_update_77167 : array_update_77156[0];
  assign array_update_77169[1] = add_76070 == 32'h0000_0001 ? array_update_77167 : array_update_77156[1];
  assign array_update_77169[2] = add_76070 == 32'h0000_0002 ? array_update_77167 : array_update_77156[2];
  assign array_update_77169[3] = add_76070 == 32'h0000_0003 ? array_update_77167 : array_update_77156[3];
  assign array_update_77169[4] = add_76070 == 32'h0000_0004 ? array_update_77167 : array_update_77156[4];
  assign array_update_77169[5] = add_76070 == 32'h0000_0005 ? array_update_77167 : array_update_77156[5];
  assign array_update_77169[6] = add_76070 == 32'h0000_0006 ? array_update_77167 : array_update_77156[6];
  assign array_update_77169[7] = add_76070 == 32'h0000_0007 ? array_update_77167 : array_update_77156[7];
  assign array_update_77169[8] = add_76070 == 32'h0000_0008 ? array_update_77167 : array_update_77156[8];
  assign array_update_77169[9] = add_76070 == 32'h0000_0009 ? array_update_77167 : array_update_77156[9];
  assign array_index_77171 = array_update_72021[add_77168 > 32'h0000_0009 ? 4'h9 : add_77168[3:0]];
  assign array_index_77172 = array_update_77169[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_77176 = smul32b_32b_x_32b(array_index_76077[add_77168 > 32'h0000_0009 ? 4'h9 : add_77168[3:0]], array_index_77171[add_77153 > 32'h0000_0009 ? 4'h9 : add_77153[3:0]]);
  assign add_77178 = array_index_77172[add_77153 > 32'h0000_0009 ? 4'h9 : add_77153[3:0]] + smul_77176;
  assign array_update_77180[0] = add_77153 == 32'h0000_0000 ? add_77178 : array_index_77172[0];
  assign array_update_77180[1] = add_77153 == 32'h0000_0001 ? add_77178 : array_index_77172[1];
  assign array_update_77180[2] = add_77153 == 32'h0000_0002 ? add_77178 : array_index_77172[2];
  assign array_update_77180[3] = add_77153 == 32'h0000_0003 ? add_77178 : array_index_77172[3];
  assign array_update_77180[4] = add_77153 == 32'h0000_0004 ? add_77178 : array_index_77172[4];
  assign array_update_77180[5] = add_77153 == 32'h0000_0005 ? add_77178 : array_index_77172[5];
  assign array_update_77180[6] = add_77153 == 32'h0000_0006 ? add_77178 : array_index_77172[6];
  assign array_update_77180[7] = add_77153 == 32'h0000_0007 ? add_77178 : array_index_77172[7];
  assign array_update_77180[8] = add_77153 == 32'h0000_0008 ? add_77178 : array_index_77172[8];
  assign array_update_77180[9] = add_77153 == 32'h0000_0009 ? add_77178 : array_index_77172[9];
  assign add_77181 = add_77168 + 32'h0000_0001;
  assign array_update_77182[0] = add_76070 == 32'h0000_0000 ? array_update_77180 : array_update_77169[0];
  assign array_update_77182[1] = add_76070 == 32'h0000_0001 ? array_update_77180 : array_update_77169[1];
  assign array_update_77182[2] = add_76070 == 32'h0000_0002 ? array_update_77180 : array_update_77169[2];
  assign array_update_77182[3] = add_76070 == 32'h0000_0003 ? array_update_77180 : array_update_77169[3];
  assign array_update_77182[4] = add_76070 == 32'h0000_0004 ? array_update_77180 : array_update_77169[4];
  assign array_update_77182[5] = add_76070 == 32'h0000_0005 ? array_update_77180 : array_update_77169[5];
  assign array_update_77182[6] = add_76070 == 32'h0000_0006 ? array_update_77180 : array_update_77169[6];
  assign array_update_77182[7] = add_76070 == 32'h0000_0007 ? array_update_77180 : array_update_77169[7];
  assign array_update_77182[8] = add_76070 == 32'h0000_0008 ? array_update_77180 : array_update_77169[8];
  assign array_update_77182[9] = add_76070 == 32'h0000_0009 ? array_update_77180 : array_update_77169[9];
  assign array_index_77184 = array_update_72021[add_77181 > 32'h0000_0009 ? 4'h9 : add_77181[3:0]];
  assign array_index_77185 = array_update_77182[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_77189 = smul32b_32b_x_32b(array_index_76077[add_77181 > 32'h0000_0009 ? 4'h9 : add_77181[3:0]], array_index_77184[add_77153 > 32'h0000_0009 ? 4'h9 : add_77153[3:0]]);
  assign add_77191 = array_index_77185[add_77153 > 32'h0000_0009 ? 4'h9 : add_77153[3:0]] + smul_77189;
  assign array_update_77193[0] = add_77153 == 32'h0000_0000 ? add_77191 : array_index_77185[0];
  assign array_update_77193[1] = add_77153 == 32'h0000_0001 ? add_77191 : array_index_77185[1];
  assign array_update_77193[2] = add_77153 == 32'h0000_0002 ? add_77191 : array_index_77185[2];
  assign array_update_77193[3] = add_77153 == 32'h0000_0003 ? add_77191 : array_index_77185[3];
  assign array_update_77193[4] = add_77153 == 32'h0000_0004 ? add_77191 : array_index_77185[4];
  assign array_update_77193[5] = add_77153 == 32'h0000_0005 ? add_77191 : array_index_77185[5];
  assign array_update_77193[6] = add_77153 == 32'h0000_0006 ? add_77191 : array_index_77185[6];
  assign array_update_77193[7] = add_77153 == 32'h0000_0007 ? add_77191 : array_index_77185[7];
  assign array_update_77193[8] = add_77153 == 32'h0000_0008 ? add_77191 : array_index_77185[8];
  assign array_update_77193[9] = add_77153 == 32'h0000_0009 ? add_77191 : array_index_77185[9];
  assign add_77194 = add_77181 + 32'h0000_0001;
  assign array_update_77195[0] = add_76070 == 32'h0000_0000 ? array_update_77193 : array_update_77182[0];
  assign array_update_77195[1] = add_76070 == 32'h0000_0001 ? array_update_77193 : array_update_77182[1];
  assign array_update_77195[2] = add_76070 == 32'h0000_0002 ? array_update_77193 : array_update_77182[2];
  assign array_update_77195[3] = add_76070 == 32'h0000_0003 ? array_update_77193 : array_update_77182[3];
  assign array_update_77195[4] = add_76070 == 32'h0000_0004 ? array_update_77193 : array_update_77182[4];
  assign array_update_77195[5] = add_76070 == 32'h0000_0005 ? array_update_77193 : array_update_77182[5];
  assign array_update_77195[6] = add_76070 == 32'h0000_0006 ? array_update_77193 : array_update_77182[6];
  assign array_update_77195[7] = add_76070 == 32'h0000_0007 ? array_update_77193 : array_update_77182[7];
  assign array_update_77195[8] = add_76070 == 32'h0000_0008 ? array_update_77193 : array_update_77182[8];
  assign array_update_77195[9] = add_76070 == 32'h0000_0009 ? array_update_77193 : array_update_77182[9];
  assign array_index_77197 = array_update_72021[add_77194 > 32'h0000_0009 ? 4'h9 : add_77194[3:0]];
  assign array_index_77198 = array_update_77195[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_77202 = smul32b_32b_x_32b(array_index_76077[add_77194 > 32'h0000_0009 ? 4'h9 : add_77194[3:0]], array_index_77197[add_77153 > 32'h0000_0009 ? 4'h9 : add_77153[3:0]]);
  assign add_77204 = array_index_77198[add_77153 > 32'h0000_0009 ? 4'h9 : add_77153[3:0]] + smul_77202;
  assign array_update_77206[0] = add_77153 == 32'h0000_0000 ? add_77204 : array_index_77198[0];
  assign array_update_77206[1] = add_77153 == 32'h0000_0001 ? add_77204 : array_index_77198[1];
  assign array_update_77206[2] = add_77153 == 32'h0000_0002 ? add_77204 : array_index_77198[2];
  assign array_update_77206[3] = add_77153 == 32'h0000_0003 ? add_77204 : array_index_77198[3];
  assign array_update_77206[4] = add_77153 == 32'h0000_0004 ? add_77204 : array_index_77198[4];
  assign array_update_77206[5] = add_77153 == 32'h0000_0005 ? add_77204 : array_index_77198[5];
  assign array_update_77206[6] = add_77153 == 32'h0000_0006 ? add_77204 : array_index_77198[6];
  assign array_update_77206[7] = add_77153 == 32'h0000_0007 ? add_77204 : array_index_77198[7];
  assign array_update_77206[8] = add_77153 == 32'h0000_0008 ? add_77204 : array_index_77198[8];
  assign array_update_77206[9] = add_77153 == 32'h0000_0009 ? add_77204 : array_index_77198[9];
  assign add_77207 = add_77194 + 32'h0000_0001;
  assign array_update_77208[0] = add_76070 == 32'h0000_0000 ? array_update_77206 : array_update_77195[0];
  assign array_update_77208[1] = add_76070 == 32'h0000_0001 ? array_update_77206 : array_update_77195[1];
  assign array_update_77208[2] = add_76070 == 32'h0000_0002 ? array_update_77206 : array_update_77195[2];
  assign array_update_77208[3] = add_76070 == 32'h0000_0003 ? array_update_77206 : array_update_77195[3];
  assign array_update_77208[4] = add_76070 == 32'h0000_0004 ? array_update_77206 : array_update_77195[4];
  assign array_update_77208[5] = add_76070 == 32'h0000_0005 ? array_update_77206 : array_update_77195[5];
  assign array_update_77208[6] = add_76070 == 32'h0000_0006 ? array_update_77206 : array_update_77195[6];
  assign array_update_77208[7] = add_76070 == 32'h0000_0007 ? array_update_77206 : array_update_77195[7];
  assign array_update_77208[8] = add_76070 == 32'h0000_0008 ? array_update_77206 : array_update_77195[8];
  assign array_update_77208[9] = add_76070 == 32'h0000_0009 ? array_update_77206 : array_update_77195[9];
  assign array_index_77210 = array_update_72021[add_77207 > 32'h0000_0009 ? 4'h9 : add_77207[3:0]];
  assign array_index_77211 = array_update_77208[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_77215 = smul32b_32b_x_32b(array_index_76077[add_77207 > 32'h0000_0009 ? 4'h9 : add_77207[3:0]], array_index_77210[add_77153 > 32'h0000_0009 ? 4'h9 : add_77153[3:0]]);
  assign add_77217 = array_index_77211[add_77153 > 32'h0000_0009 ? 4'h9 : add_77153[3:0]] + smul_77215;
  assign array_update_77219[0] = add_77153 == 32'h0000_0000 ? add_77217 : array_index_77211[0];
  assign array_update_77219[1] = add_77153 == 32'h0000_0001 ? add_77217 : array_index_77211[1];
  assign array_update_77219[2] = add_77153 == 32'h0000_0002 ? add_77217 : array_index_77211[2];
  assign array_update_77219[3] = add_77153 == 32'h0000_0003 ? add_77217 : array_index_77211[3];
  assign array_update_77219[4] = add_77153 == 32'h0000_0004 ? add_77217 : array_index_77211[4];
  assign array_update_77219[5] = add_77153 == 32'h0000_0005 ? add_77217 : array_index_77211[5];
  assign array_update_77219[6] = add_77153 == 32'h0000_0006 ? add_77217 : array_index_77211[6];
  assign array_update_77219[7] = add_77153 == 32'h0000_0007 ? add_77217 : array_index_77211[7];
  assign array_update_77219[8] = add_77153 == 32'h0000_0008 ? add_77217 : array_index_77211[8];
  assign array_update_77219[9] = add_77153 == 32'h0000_0009 ? add_77217 : array_index_77211[9];
  assign add_77220 = add_77207 + 32'h0000_0001;
  assign array_update_77221[0] = add_76070 == 32'h0000_0000 ? array_update_77219 : array_update_77208[0];
  assign array_update_77221[1] = add_76070 == 32'h0000_0001 ? array_update_77219 : array_update_77208[1];
  assign array_update_77221[2] = add_76070 == 32'h0000_0002 ? array_update_77219 : array_update_77208[2];
  assign array_update_77221[3] = add_76070 == 32'h0000_0003 ? array_update_77219 : array_update_77208[3];
  assign array_update_77221[4] = add_76070 == 32'h0000_0004 ? array_update_77219 : array_update_77208[4];
  assign array_update_77221[5] = add_76070 == 32'h0000_0005 ? array_update_77219 : array_update_77208[5];
  assign array_update_77221[6] = add_76070 == 32'h0000_0006 ? array_update_77219 : array_update_77208[6];
  assign array_update_77221[7] = add_76070 == 32'h0000_0007 ? array_update_77219 : array_update_77208[7];
  assign array_update_77221[8] = add_76070 == 32'h0000_0008 ? array_update_77219 : array_update_77208[8];
  assign array_update_77221[9] = add_76070 == 32'h0000_0009 ? array_update_77219 : array_update_77208[9];
  assign array_index_77223 = array_update_72021[add_77220 > 32'h0000_0009 ? 4'h9 : add_77220[3:0]];
  assign array_index_77224 = array_update_77221[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_77228 = smul32b_32b_x_32b(array_index_76077[add_77220 > 32'h0000_0009 ? 4'h9 : add_77220[3:0]], array_index_77223[add_77153 > 32'h0000_0009 ? 4'h9 : add_77153[3:0]]);
  assign add_77230 = array_index_77224[add_77153 > 32'h0000_0009 ? 4'h9 : add_77153[3:0]] + smul_77228;
  assign array_update_77232[0] = add_77153 == 32'h0000_0000 ? add_77230 : array_index_77224[0];
  assign array_update_77232[1] = add_77153 == 32'h0000_0001 ? add_77230 : array_index_77224[1];
  assign array_update_77232[2] = add_77153 == 32'h0000_0002 ? add_77230 : array_index_77224[2];
  assign array_update_77232[3] = add_77153 == 32'h0000_0003 ? add_77230 : array_index_77224[3];
  assign array_update_77232[4] = add_77153 == 32'h0000_0004 ? add_77230 : array_index_77224[4];
  assign array_update_77232[5] = add_77153 == 32'h0000_0005 ? add_77230 : array_index_77224[5];
  assign array_update_77232[6] = add_77153 == 32'h0000_0006 ? add_77230 : array_index_77224[6];
  assign array_update_77232[7] = add_77153 == 32'h0000_0007 ? add_77230 : array_index_77224[7];
  assign array_update_77232[8] = add_77153 == 32'h0000_0008 ? add_77230 : array_index_77224[8];
  assign array_update_77232[9] = add_77153 == 32'h0000_0009 ? add_77230 : array_index_77224[9];
  assign add_77233 = add_77220 + 32'h0000_0001;
  assign array_update_77234[0] = add_76070 == 32'h0000_0000 ? array_update_77232 : array_update_77221[0];
  assign array_update_77234[1] = add_76070 == 32'h0000_0001 ? array_update_77232 : array_update_77221[1];
  assign array_update_77234[2] = add_76070 == 32'h0000_0002 ? array_update_77232 : array_update_77221[2];
  assign array_update_77234[3] = add_76070 == 32'h0000_0003 ? array_update_77232 : array_update_77221[3];
  assign array_update_77234[4] = add_76070 == 32'h0000_0004 ? array_update_77232 : array_update_77221[4];
  assign array_update_77234[5] = add_76070 == 32'h0000_0005 ? array_update_77232 : array_update_77221[5];
  assign array_update_77234[6] = add_76070 == 32'h0000_0006 ? array_update_77232 : array_update_77221[6];
  assign array_update_77234[7] = add_76070 == 32'h0000_0007 ? array_update_77232 : array_update_77221[7];
  assign array_update_77234[8] = add_76070 == 32'h0000_0008 ? array_update_77232 : array_update_77221[8];
  assign array_update_77234[9] = add_76070 == 32'h0000_0009 ? array_update_77232 : array_update_77221[9];
  assign array_index_77236 = array_update_72021[add_77233 > 32'h0000_0009 ? 4'h9 : add_77233[3:0]];
  assign array_index_77237 = array_update_77234[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_77241 = smul32b_32b_x_32b(array_index_76077[add_77233 > 32'h0000_0009 ? 4'h9 : add_77233[3:0]], array_index_77236[add_77153 > 32'h0000_0009 ? 4'h9 : add_77153[3:0]]);
  assign add_77243 = array_index_77237[add_77153 > 32'h0000_0009 ? 4'h9 : add_77153[3:0]] + smul_77241;
  assign array_update_77245[0] = add_77153 == 32'h0000_0000 ? add_77243 : array_index_77237[0];
  assign array_update_77245[1] = add_77153 == 32'h0000_0001 ? add_77243 : array_index_77237[1];
  assign array_update_77245[2] = add_77153 == 32'h0000_0002 ? add_77243 : array_index_77237[2];
  assign array_update_77245[3] = add_77153 == 32'h0000_0003 ? add_77243 : array_index_77237[3];
  assign array_update_77245[4] = add_77153 == 32'h0000_0004 ? add_77243 : array_index_77237[4];
  assign array_update_77245[5] = add_77153 == 32'h0000_0005 ? add_77243 : array_index_77237[5];
  assign array_update_77245[6] = add_77153 == 32'h0000_0006 ? add_77243 : array_index_77237[6];
  assign array_update_77245[7] = add_77153 == 32'h0000_0007 ? add_77243 : array_index_77237[7];
  assign array_update_77245[8] = add_77153 == 32'h0000_0008 ? add_77243 : array_index_77237[8];
  assign array_update_77245[9] = add_77153 == 32'h0000_0009 ? add_77243 : array_index_77237[9];
  assign add_77246 = add_77233 + 32'h0000_0001;
  assign array_update_77247[0] = add_76070 == 32'h0000_0000 ? array_update_77245 : array_update_77234[0];
  assign array_update_77247[1] = add_76070 == 32'h0000_0001 ? array_update_77245 : array_update_77234[1];
  assign array_update_77247[2] = add_76070 == 32'h0000_0002 ? array_update_77245 : array_update_77234[2];
  assign array_update_77247[3] = add_76070 == 32'h0000_0003 ? array_update_77245 : array_update_77234[3];
  assign array_update_77247[4] = add_76070 == 32'h0000_0004 ? array_update_77245 : array_update_77234[4];
  assign array_update_77247[5] = add_76070 == 32'h0000_0005 ? array_update_77245 : array_update_77234[5];
  assign array_update_77247[6] = add_76070 == 32'h0000_0006 ? array_update_77245 : array_update_77234[6];
  assign array_update_77247[7] = add_76070 == 32'h0000_0007 ? array_update_77245 : array_update_77234[7];
  assign array_update_77247[8] = add_76070 == 32'h0000_0008 ? array_update_77245 : array_update_77234[8];
  assign array_update_77247[9] = add_76070 == 32'h0000_0009 ? array_update_77245 : array_update_77234[9];
  assign array_index_77249 = array_update_72021[add_77246 > 32'h0000_0009 ? 4'h9 : add_77246[3:0]];
  assign array_index_77250 = array_update_77247[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_77254 = smul32b_32b_x_32b(array_index_76077[add_77246 > 32'h0000_0009 ? 4'h9 : add_77246[3:0]], array_index_77249[add_77153 > 32'h0000_0009 ? 4'h9 : add_77153[3:0]]);
  assign add_77256 = array_index_77250[add_77153 > 32'h0000_0009 ? 4'h9 : add_77153[3:0]] + smul_77254;
  assign array_update_77258[0] = add_77153 == 32'h0000_0000 ? add_77256 : array_index_77250[0];
  assign array_update_77258[1] = add_77153 == 32'h0000_0001 ? add_77256 : array_index_77250[1];
  assign array_update_77258[2] = add_77153 == 32'h0000_0002 ? add_77256 : array_index_77250[2];
  assign array_update_77258[3] = add_77153 == 32'h0000_0003 ? add_77256 : array_index_77250[3];
  assign array_update_77258[4] = add_77153 == 32'h0000_0004 ? add_77256 : array_index_77250[4];
  assign array_update_77258[5] = add_77153 == 32'h0000_0005 ? add_77256 : array_index_77250[5];
  assign array_update_77258[6] = add_77153 == 32'h0000_0006 ? add_77256 : array_index_77250[6];
  assign array_update_77258[7] = add_77153 == 32'h0000_0007 ? add_77256 : array_index_77250[7];
  assign array_update_77258[8] = add_77153 == 32'h0000_0008 ? add_77256 : array_index_77250[8];
  assign array_update_77258[9] = add_77153 == 32'h0000_0009 ? add_77256 : array_index_77250[9];
  assign add_77259 = add_77246 + 32'h0000_0001;
  assign array_update_77260[0] = add_76070 == 32'h0000_0000 ? array_update_77258 : array_update_77247[0];
  assign array_update_77260[1] = add_76070 == 32'h0000_0001 ? array_update_77258 : array_update_77247[1];
  assign array_update_77260[2] = add_76070 == 32'h0000_0002 ? array_update_77258 : array_update_77247[2];
  assign array_update_77260[3] = add_76070 == 32'h0000_0003 ? array_update_77258 : array_update_77247[3];
  assign array_update_77260[4] = add_76070 == 32'h0000_0004 ? array_update_77258 : array_update_77247[4];
  assign array_update_77260[5] = add_76070 == 32'h0000_0005 ? array_update_77258 : array_update_77247[5];
  assign array_update_77260[6] = add_76070 == 32'h0000_0006 ? array_update_77258 : array_update_77247[6];
  assign array_update_77260[7] = add_76070 == 32'h0000_0007 ? array_update_77258 : array_update_77247[7];
  assign array_update_77260[8] = add_76070 == 32'h0000_0008 ? array_update_77258 : array_update_77247[8];
  assign array_update_77260[9] = add_76070 == 32'h0000_0009 ? array_update_77258 : array_update_77247[9];
  assign array_index_77262 = array_update_72021[add_77259 > 32'h0000_0009 ? 4'h9 : add_77259[3:0]];
  assign array_index_77263 = array_update_77260[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_77267 = smul32b_32b_x_32b(array_index_76077[add_77259 > 32'h0000_0009 ? 4'h9 : add_77259[3:0]], array_index_77262[add_77153 > 32'h0000_0009 ? 4'h9 : add_77153[3:0]]);
  assign add_77269 = array_index_77263[add_77153 > 32'h0000_0009 ? 4'h9 : add_77153[3:0]] + smul_77267;
  assign array_update_77271[0] = add_77153 == 32'h0000_0000 ? add_77269 : array_index_77263[0];
  assign array_update_77271[1] = add_77153 == 32'h0000_0001 ? add_77269 : array_index_77263[1];
  assign array_update_77271[2] = add_77153 == 32'h0000_0002 ? add_77269 : array_index_77263[2];
  assign array_update_77271[3] = add_77153 == 32'h0000_0003 ? add_77269 : array_index_77263[3];
  assign array_update_77271[4] = add_77153 == 32'h0000_0004 ? add_77269 : array_index_77263[4];
  assign array_update_77271[5] = add_77153 == 32'h0000_0005 ? add_77269 : array_index_77263[5];
  assign array_update_77271[6] = add_77153 == 32'h0000_0006 ? add_77269 : array_index_77263[6];
  assign array_update_77271[7] = add_77153 == 32'h0000_0007 ? add_77269 : array_index_77263[7];
  assign array_update_77271[8] = add_77153 == 32'h0000_0008 ? add_77269 : array_index_77263[8];
  assign array_update_77271[9] = add_77153 == 32'h0000_0009 ? add_77269 : array_index_77263[9];
  assign add_77272 = add_77259 + 32'h0000_0001;
  assign array_update_77273[0] = add_76070 == 32'h0000_0000 ? array_update_77271 : array_update_77260[0];
  assign array_update_77273[1] = add_76070 == 32'h0000_0001 ? array_update_77271 : array_update_77260[1];
  assign array_update_77273[2] = add_76070 == 32'h0000_0002 ? array_update_77271 : array_update_77260[2];
  assign array_update_77273[3] = add_76070 == 32'h0000_0003 ? array_update_77271 : array_update_77260[3];
  assign array_update_77273[4] = add_76070 == 32'h0000_0004 ? array_update_77271 : array_update_77260[4];
  assign array_update_77273[5] = add_76070 == 32'h0000_0005 ? array_update_77271 : array_update_77260[5];
  assign array_update_77273[6] = add_76070 == 32'h0000_0006 ? array_update_77271 : array_update_77260[6];
  assign array_update_77273[7] = add_76070 == 32'h0000_0007 ? array_update_77271 : array_update_77260[7];
  assign array_update_77273[8] = add_76070 == 32'h0000_0008 ? array_update_77271 : array_update_77260[8];
  assign array_update_77273[9] = add_76070 == 32'h0000_0009 ? array_update_77271 : array_update_77260[9];
  assign array_index_77275 = array_update_72021[add_77272 > 32'h0000_0009 ? 4'h9 : add_77272[3:0]];
  assign array_index_77276 = array_update_77273[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_77280 = smul32b_32b_x_32b(array_index_76077[add_77272 > 32'h0000_0009 ? 4'h9 : add_77272[3:0]], array_index_77275[add_77153 > 32'h0000_0009 ? 4'h9 : add_77153[3:0]]);
  assign add_77282 = array_index_77276[add_77153 > 32'h0000_0009 ? 4'h9 : add_77153[3:0]] + smul_77280;
  assign array_update_77283[0] = add_77153 == 32'h0000_0000 ? add_77282 : array_index_77276[0];
  assign array_update_77283[1] = add_77153 == 32'h0000_0001 ? add_77282 : array_index_77276[1];
  assign array_update_77283[2] = add_77153 == 32'h0000_0002 ? add_77282 : array_index_77276[2];
  assign array_update_77283[3] = add_77153 == 32'h0000_0003 ? add_77282 : array_index_77276[3];
  assign array_update_77283[4] = add_77153 == 32'h0000_0004 ? add_77282 : array_index_77276[4];
  assign array_update_77283[5] = add_77153 == 32'h0000_0005 ? add_77282 : array_index_77276[5];
  assign array_update_77283[6] = add_77153 == 32'h0000_0006 ? add_77282 : array_index_77276[6];
  assign array_update_77283[7] = add_77153 == 32'h0000_0007 ? add_77282 : array_index_77276[7];
  assign array_update_77283[8] = add_77153 == 32'h0000_0008 ? add_77282 : array_index_77276[8];
  assign array_update_77283[9] = add_77153 == 32'h0000_0009 ? add_77282 : array_index_77276[9];
  assign array_update_77284[0] = add_76070 == 32'h0000_0000 ? array_update_77283 : array_update_77273[0];
  assign array_update_77284[1] = add_76070 == 32'h0000_0001 ? array_update_77283 : array_update_77273[1];
  assign array_update_77284[2] = add_76070 == 32'h0000_0002 ? array_update_77283 : array_update_77273[2];
  assign array_update_77284[3] = add_76070 == 32'h0000_0003 ? array_update_77283 : array_update_77273[3];
  assign array_update_77284[4] = add_76070 == 32'h0000_0004 ? array_update_77283 : array_update_77273[4];
  assign array_update_77284[5] = add_76070 == 32'h0000_0005 ? array_update_77283 : array_update_77273[5];
  assign array_update_77284[6] = add_76070 == 32'h0000_0006 ? array_update_77283 : array_update_77273[6];
  assign array_update_77284[7] = add_76070 == 32'h0000_0007 ? array_update_77283 : array_update_77273[7];
  assign array_update_77284[8] = add_76070 == 32'h0000_0008 ? array_update_77283 : array_update_77273[8];
  assign array_update_77284[9] = add_76070 == 32'h0000_0009 ? array_update_77283 : array_update_77273[9];
  assign array_index_77286 = array_update_77284[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign add_77288 = add_77153 + 32'h0000_0001;
  assign array_update_77289[0] = add_77288 == 32'h0000_0000 ? 32'h0000_0000 : array_index_77286[0];
  assign array_update_77289[1] = add_77288 == 32'h0000_0001 ? 32'h0000_0000 : array_index_77286[1];
  assign array_update_77289[2] = add_77288 == 32'h0000_0002 ? 32'h0000_0000 : array_index_77286[2];
  assign array_update_77289[3] = add_77288 == 32'h0000_0003 ? 32'h0000_0000 : array_index_77286[3];
  assign array_update_77289[4] = add_77288 == 32'h0000_0004 ? 32'h0000_0000 : array_index_77286[4];
  assign array_update_77289[5] = add_77288 == 32'h0000_0005 ? 32'h0000_0000 : array_index_77286[5];
  assign array_update_77289[6] = add_77288 == 32'h0000_0006 ? 32'h0000_0000 : array_index_77286[6];
  assign array_update_77289[7] = add_77288 == 32'h0000_0007 ? 32'h0000_0000 : array_index_77286[7];
  assign array_update_77289[8] = add_77288 == 32'h0000_0008 ? 32'h0000_0000 : array_index_77286[8];
  assign array_update_77289[9] = add_77288 == 32'h0000_0009 ? 32'h0000_0000 : array_index_77286[9];
  assign literal_77290 = 32'h0000_0000;
  assign array_update_77291[0] = add_76070 == 32'h0000_0000 ? array_update_77289 : array_update_77284[0];
  assign array_update_77291[1] = add_76070 == 32'h0000_0001 ? array_update_77289 : array_update_77284[1];
  assign array_update_77291[2] = add_76070 == 32'h0000_0002 ? array_update_77289 : array_update_77284[2];
  assign array_update_77291[3] = add_76070 == 32'h0000_0003 ? array_update_77289 : array_update_77284[3];
  assign array_update_77291[4] = add_76070 == 32'h0000_0004 ? array_update_77289 : array_update_77284[4];
  assign array_update_77291[5] = add_76070 == 32'h0000_0005 ? array_update_77289 : array_update_77284[5];
  assign array_update_77291[6] = add_76070 == 32'h0000_0006 ? array_update_77289 : array_update_77284[6];
  assign array_update_77291[7] = add_76070 == 32'h0000_0007 ? array_update_77289 : array_update_77284[7];
  assign array_update_77291[8] = add_76070 == 32'h0000_0008 ? array_update_77289 : array_update_77284[8];
  assign array_update_77291[9] = add_76070 == 32'h0000_0009 ? array_update_77289 : array_update_77284[9];
  assign array_index_77293 = array_update_72021[literal_77290 > 32'h0000_0009 ? 4'h9 : literal_77290[3:0]];
  assign array_index_77294 = array_update_77291[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_77298 = smul32b_32b_x_32b(array_index_76077[literal_77290 > 32'h0000_0009 ? 4'h9 : literal_77290[3:0]], array_index_77293[add_77288 > 32'h0000_0009 ? 4'h9 : add_77288[3:0]]);
  assign add_77300 = array_index_77294[add_77288 > 32'h0000_0009 ? 4'h9 : add_77288[3:0]] + smul_77298;
  assign array_update_77302[0] = add_77288 == 32'h0000_0000 ? add_77300 : array_index_77294[0];
  assign array_update_77302[1] = add_77288 == 32'h0000_0001 ? add_77300 : array_index_77294[1];
  assign array_update_77302[2] = add_77288 == 32'h0000_0002 ? add_77300 : array_index_77294[2];
  assign array_update_77302[3] = add_77288 == 32'h0000_0003 ? add_77300 : array_index_77294[3];
  assign array_update_77302[4] = add_77288 == 32'h0000_0004 ? add_77300 : array_index_77294[4];
  assign array_update_77302[5] = add_77288 == 32'h0000_0005 ? add_77300 : array_index_77294[5];
  assign array_update_77302[6] = add_77288 == 32'h0000_0006 ? add_77300 : array_index_77294[6];
  assign array_update_77302[7] = add_77288 == 32'h0000_0007 ? add_77300 : array_index_77294[7];
  assign array_update_77302[8] = add_77288 == 32'h0000_0008 ? add_77300 : array_index_77294[8];
  assign array_update_77302[9] = add_77288 == 32'h0000_0009 ? add_77300 : array_index_77294[9];
  assign add_77303 = literal_77290 + 32'h0000_0001;
  assign array_update_77304[0] = add_76070 == 32'h0000_0000 ? array_update_77302 : array_update_77291[0];
  assign array_update_77304[1] = add_76070 == 32'h0000_0001 ? array_update_77302 : array_update_77291[1];
  assign array_update_77304[2] = add_76070 == 32'h0000_0002 ? array_update_77302 : array_update_77291[2];
  assign array_update_77304[3] = add_76070 == 32'h0000_0003 ? array_update_77302 : array_update_77291[3];
  assign array_update_77304[4] = add_76070 == 32'h0000_0004 ? array_update_77302 : array_update_77291[4];
  assign array_update_77304[5] = add_76070 == 32'h0000_0005 ? array_update_77302 : array_update_77291[5];
  assign array_update_77304[6] = add_76070 == 32'h0000_0006 ? array_update_77302 : array_update_77291[6];
  assign array_update_77304[7] = add_76070 == 32'h0000_0007 ? array_update_77302 : array_update_77291[7];
  assign array_update_77304[8] = add_76070 == 32'h0000_0008 ? array_update_77302 : array_update_77291[8];
  assign array_update_77304[9] = add_76070 == 32'h0000_0009 ? array_update_77302 : array_update_77291[9];
  assign array_index_77306 = array_update_72021[add_77303 > 32'h0000_0009 ? 4'h9 : add_77303[3:0]];
  assign array_index_77307 = array_update_77304[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_77311 = smul32b_32b_x_32b(array_index_76077[add_77303 > 32'h0000_0009 ? 4'h9 : add_77303[3:0]], array_index_77306[add_77288 > 32'h0000_0009 ? 4'h9 : add_77288[3:0]]);
  assign add_77313 = array_index_77307[add_77288 > 32'h0000_0009 ? 4'h9 : add_77288[3:0]] + smul_77311;
  assign array_update_77315[0] = add_77288 == 32'h0000_0000 ? add_77313 : array_index_77307[0];
  assign array_update_77315[1] = add_77288 == 32'h0000_0001 ? add_77313 : array_index_77307[1];
  assign array_update_77315[2] = add_77288 == 32'h0000_0002 ? add_77313 : array_index_77307[2];
  assign array_update_77315[3] = add_77288 == 32'h0000_0003 ? add_77313 : array_index_77307[3];
  assign array_update_77315[4] = add_77288 == 32'h0000_0004 ? add_77313 : array_index_77307[4];
  assign array_update_77315[5] = add_77288 == 32'h0000_0005 ? add_77313 : array_index_77307[5];
  assign array_update_77315[6] = add_77288 == 32'h0000_0006 ? add_77313 : array_index_77307[6];
  assign array_update_77315[7] = add_77288 == 32'h0000_0007 ? add_77313 : array_index_77307[7];
  assign array_update_77315[8] = add_77288 == 32'h0000_0008 ? add_77313 : array_index_77307[8];
  assign array_update_77315[9] = add_77288 == 32'h0000_0009 ? add_77313 : array_index_77307[9];
  assign add_77316 = add_77303 + 32'h0000_0001;
  assign array_update_77317[0] = add_76070 == 32'h0000_0000 ? array_update_77315 : array_update_77304[0];
  assign array_update_77317[1] = add_76070 == 32'h0000_0001 ? array_update_77315 : array_update_77304[1];
  assign array_update_77317[2] = add_76070 == 32'h0000_0002 ? array_update_77315 : array_update_77304[2];
  assign array_update_77317[3] = add_76070 == 32'h0000_0003 ? array_update_77315 : array_update_77304[3];
  assign array_update_77317[4] = add_76070 == 32'h0000_0004 ? array_update_77315 : array_update_77304[4];
  assign array_update_77317[5] = add_76070 == 32'h0000_0005 ? array_update_77315 : array_update_77304[5];
  assign array_update_77317[6] = add_76070 == 32'h0000_0006 ? array_update_77315 : array_update_77304[6];
  assign array_update_77317[7] = add_76070 == 32'h0000_0007 ? array_update_77315 : array_update_77304[7];
  assign array_update_77317[8] = add_76070 == 32'h0000_0008 ? array_update_77315 : array_update_77304[8];
  assign array_update_77317[9] = add_76070 == 32'h0000_0009 ? array_update_77315 : array_update_77304[9];
  assign array_index_77319 = array_update_72021[add_77316 > 32'h0000_0009 ? 4'h9 : add_77316[3:0]];
  assign array_index_77320 = array_update_77317[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_77324 = smul32b_32b_x_32b(array_index_76077[add_77316 > 32'h0000_0009 ? 4'h9 : add_77316[3:0]], array_index_77319[add_77288 > 32'h0000_0009 ? 4'h9 : add_77288[3:0]]);
  assign add_77326 = array_index_77320[add_77288 > 32'h0000_0009 ? 4'h9 : add_77288[3:0]] + smul_77324;
  assign array_update_77328[0] = add_77288 == 32'h0000_0000 ? add_77326 : array_index_77320[0];
  assign array_update_77328[1] = add_77288 == 32'h0000_0001 ? add_77326 : array_index_77320[1];
  assign array_update_77328[2] = add_77288 == 32'h0000_0002 ? add_77326 : array_index_77320[2];
  assign array_update_77328[3] = add_77288 == 32'h0000_0003 ? add_77326 : array_index_77320[3];
  assign array_update_77328[4] = add_77288 == 32'h0000_0004 ? add_77326 : array_index_77320[4];
  assign array_update_77328[5] = add_77288 == 32'h0000_0005 ? add_77326 : array_index_77320[5];
  assign array_update_77328[6] = add_77288 == 32'h0000_0006 ? add_77326 : array_index_77320[6];
  assign array_update_77328[7] = add_77288 == 32'h0000_0007 ? add_77326 : array_index_77320[7];
  assign array_update_77328[8] = add_77288 == 32'h0000_0008 ? add_77326 : array_index_77320[8];
  assign array_update_77328[9] = add_77288 == 32'h0000_0009 ? add_77326 : array_index_77320[9];
  assign add_77329 = add_77316 + 32'h0000_0001;
  assign array_update_77330[0] = add_76070 == 32'h0000_0000 ? array_update_77328 : array_update_77317[0];
  assign array_update_77330[1] = add_76070 == 32'h0000_0001 ? array_update_77328 : array_update_77317[1];
  assign array_update_77330[2] = add_76070 == 32'h0000_0002 ? array_update_77328 : array_update_77317[2];
  assign array_update_77330[3] = add_76070 == 32'h0000_0003 ? array_update_77328 : array_update_77317[3];
  assign array_update_77330[4] = add_76070 == 32'h0000_0004 ? array_update_77328 : array_update_77317[4];
  assign array_update_77330[5] = add_76070 == 32'h0000_0005 ? array_update_77328 : array_update_77317[5];
  assign array_update_77330[6] = add_76070 == 32'h0000_0006 ? array_update_77328 : array_update_77317[6];
  assign array_update_77330[7] = add_76070 == 32'h0000_0007 ? array_update_77328 : array_update_77317[7];
  assign array_update_77330[8] = add_76070 == 32'h0000_0008 ? array_update_77328 : array_update_77317[8];
  assign array_update_77330[9] = add_76070 == 32'h0000_0009 ? array_update_77328 : array_update_77317[9];
  assign array_index_77332 = array_update_72021[add_77329 > 32'h0000_0009 ? 4'h9 : add_77329[3:0]];
  assign array_index_77333 = array_update_77330[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_77337 = smul32b_32b_x_32b(array_index_76077[add_77329 > 32'h0000_0009 ? 4'h9 : add_77329[3:0]], array_index_77332[add_77288 > 32'h0000_0009 ? 4'h9 : add_77288[3:0]]);
  assign add_77339 = array_index_77333[add_77288 > 32'h0000_0009 ? 4'h9 : add_77288[3:0]] + smul_77337;
  assign array_update_77341[0] = add_77288 == 32'h0000_0000 ? add_77339 : array_index_77333[0];
  assign array_update_77341[1] = add_77288 == 32'h0000_0001 ? add_77339 : array_index_77333[1];
  assign array_update_77341[2] = add_77288 == 32'h0000_0002 ? add_77339 : array_index_77333[2];
  assign array_update_77341[3] = add_77288 == 32'h0000_0003 ? add_77339 : array_index_77333[3];
  assign array_update_77341[4] = add_77288 == 32'h0000_0004 ? add_77339 : array_index_77333[4];
  assign array_update_77341[5] = add_77288 == 32'h0000_0005 ? add_77339 : array_index_77333[5];
  assign array_update_77341[6] = add_77288 == 32'h0000_0006 ? add_77339 : array_index_77333[6];
  assign array_update_77341[7] = add_77288 == 32'h0000_0007 ? add_77339 : array_index_77333[7];
  assign array_update_77341[8] = add_77288 == 32'h0000_0008 ? add_77339 : array_index_77333[8];
  assign array_update_77341[9] = add_77288 == 32'h0000_0009 ? add_77339 : array_index_77333[9];
  assign add_77342 = add_77329 + 32'h0000_0001;
  assign array_update_77343[0] = add_76070 == 32'h0000_0000 ? array_update_77341 : array_update_77330[0];
  assign array_update_77343[1] = add_76070 == 32'h0000_0001 ? array_update_77341 : array_update_77330[1];
  assign array_update_77343[2] = add_76070 == 32'h0000_0002 ? array_update_77341 : array_update_77330[2];
  assign array_update_77343[3] = add_76070 == 32'h0000_0003 ? array_update_77341 : array_update_77330[3];
  assign array_update_77343[4] = add_76070 == 32'h0000_0004 ? array_update_77341 : array_update_77330[4];
  assign array_update_77343[5] = add_76070 == 32'h0000_0005 ? array_update_77341 : array_update_77330[5];
  assign array_update_77343[6] = add_76070 == 32'h0000_0006 ? array_update_77341 : array_update_77330[6];
  assign array_update_77343[7] = add_76070 == 32'h0000_0007 ? array_update_77341 : array_update_77330[7];
  assign array_update_77343[8] = add_76070 == 32'h0000_0008 ? array_update_77341 : array_update_77330[8];
  assign array_update_77343[9] = add_76070 == 32'h0000_0009 ? array_update_77341 : array_update_77330[9];
  assign array_index_77345 = array_update_72021[add_77342 > 32'h0000_0009 ? 4'h9 : add_77342[3:0]];
  assign array_index_77346 = array_update_77343[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_77350 = smul32b_32b_x_32b(array_index_76077[add_77342 > 32'h0000_0009 ? 4'h9 : add_77342[3:0]], array_index_77345[add_77288 > 32'h0000_0009 ? 4'h9 : add_77288[3:0]]);
  assign add_77352 = array_index_77346[add_77288 > 32'h0000_0009 ? 4'h9 : add_77288[3:0]] + smul_77350;
  assign array_update_77354[0] = add_77288 == 32'h0000_0000 ? add_77352 : array_index_77346[0];
  assign array_update_77354[1] = add_77288 == 32'h0000_0001 ? add_77352 : array_index_77346[1];
  assign array_update_77354[2] = add_77288 == 32'h0000_0002 ? add_77352 : array_index_77346[2];
  assign array_update_77354[3] = add_77288 == 32'h0000_0003 ? add_77352 : array_index_77346[3];
  assign array_update_77354[4] = add_77288 == 32'h0000_0004 ? add_77352 : array_index_77346[4];
  assign array_update_77354[5] = add_77288 == 32'h0000_0005 ? add_77352 : array_index_77346[5];
  assign array_update_77354[6] = add_77288 == 32'h0000_0006 ? add_77352 : array_index_77346[6];
  assign array_update_77354[7] = add_77288 == 32'h0000_0007 ? add_77352 : array_index_77346[7];
  assign array_update_77354[8] = add_77288 == 32'h0000_0008 ? add_77352 : array_index_77346[8];
  assign array_update_77354[9] = add_77288 == 32'h0000_0009 ? add_77352 : array_index_77346[9];
  assign add_77355 = add_77342 + 32'h0000_0001;
  assign array_update_77356[0] = add_76070 == 32'h0000_0000 ? array_update_77354 : array_update_77343[0];
  assign array_update_77356[1] = add_76070 == 32'h0000_0001 ? array_update_77354 : array_update_77343[1];
  assign array_update_77356[2] = add_76070 == 32'h0000_0002 ? array_update_77354 : array_update_77343[2];
  assign array_update_77356[3] = add_76070 == 32'h0000_0003 ? array_update_77354 : array_update_77343[3];
  assign array_update_77356[4] = add_76070 == 32'h0000_0004 ? array_update_77354 : array_update_77343[4];
  assign array_update_77356[5] = add_76070 == 32'h0000_0005 ? array_update_77354 : array_update_77343[5];
  assign array_update_77356[6] = add_76070 == 32'h0000_0006 ? array_update_77354 : array_update_77343[6];
  assign array_update_77356[7] = add_76070 == 32'h0000_0007 ? array_update_77354 : array_update_77343[7];
  assign array_update_77356[8] = add_76070 == 32'h0000_0008 ? array_update_77354 : array_update_77343[8];
  assign array_update_77356[9] = add_76070 == 32'h0000_0009 ? array_update_77354 : array_update_77343[9];
  assign array_index_77358 = array_update_72021[add_77355 > 32'h0000_0009 ? 4'h9 : add_77355[3:0]];
  assign array_index_77359 = array_update_77356[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_77363 = smul32b_32b_x_32b(array_index_76077[add_77355 > 32'h0000_0009 ? 4'h9 : add_77355[3:0]], array_index_77358[add_77288 > 32'h0000_0009 ? 4'h9 : add_77288[3:0]]);
  assign add_77365 = array_index_77359[add_77288 > 32'h0000_0009 ? 4'h9 : add_77288[3:0]] + smul_77363;
  assign array_update_77367[0] = add_77288 == 32'h0000_0000 ? add_77365 : array_index_77359[0];
  assign array_update_77367[1] = add_77288 == 32'h0000_0001 ? add_77365 : array_index_77359[1];
  assign array_update_77367[2] = add_77288 == 32'h0000_0002 ? add_77365 : array_index_77359[2];
  assign array_update_77367[3] = add_77288 == 32'h0000_0003 ? add_77365 : array_index_77359[3];
  assign array_update_77367[4] = add_77288 == 32'h0000_0004 ? add_77365 : array_index_77359[4];
  assign array_update_77367[5] = add_77288 == 32'h0000_0005 ? add_77365 : array_index_77359[5];
  assign array_update_77367[6] = add_77288 == 32'h0000_0006 ? add_77365 : array_index_77359[6];
  assign array_update_77367[7] = add_77288 == 32'h0000_0007 ? add_77365 : array_index_77359[7];
  assign array_update_77367[8] = add_77288 == 32'h0000_0008 ? add_77365 : array_index_77359[8];
  assign array_update_77367[9] = add_77288 == 32'h0000_0009 ? add_77365 : array_index_77359[9];
  assign add_77368 = add_77355 + 32'h0000_0001;
  assign array_update_77369[0] = add_76070 == 32'h0000_0000 ? array_update_77367 : array_update_77356[0];
  assign array_update_77369[1] = add_76070 == 32'h0000_0001 ? array_update_77367 : array_update_77356[1];
  assign array_update_77369[2] = add_76070 == 32'h0000_0002 ? array_update_77367 : array_update_77356[2];
  assign array_update_77369[3] = add_76070 == 32'h0000_0003 ? array_update_77367 : array_update_77356[3];
  assign array_update_77369[4] = add_76070 == 32'h0000_0004 ? array_update_77367 : array_update_77356[4];
  assign array_update_77369[5] = add_76070 == 32'h0000_0005 ? array_update_77367 : array_update_77356[5];
  assign array_update_77369[6] = add_76070 == 32'h0000_0006 ? array_update_77367 : array_update_77356[6];
  assign array_update_77369[7] = add_76070 == 32'h0000_0007 ? array_update_77367 : array_update_77356[7];
  assign array_update_77369[8] = add_76070 == 32'h0000_0008 ? array_update_77367 : array_update_77356[8];
  assign array_update_77369[9] = add_76070 == 32'h0000_0009 ? array_update_77367 : array_update_77356[9];
  assign array_index_77371 = array_update_72021[add_77368 > 32'h0000_0009 ? 4'h9 : add_77368[3:0]];
  assign array_index_77372 = array_update_77369[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_77376 = smul32b_32b_x_32b(array_index_76077[add_77368 > 32'h0000_0009 ? 4'h9 : add_77368[3:0]], array_index_77371[add_77288 > 32'h0000_0009 ? 4'h9 : add_77288[3:0]]);
  assign add_77378 = array_index_77372[add_77288 > 32'h0000_0009 ? 4'h9 : add_77288[3:0]] + smul_77376;
  assign array_update_77380[0] = add_77288 == 32'h0000_0000 ? add_77378 : array_index_77372[0];
  assign array_update_77380[1] = add_77288 == 32'h0000_0001 ? add_77378 : array_index_77372[1];
  assign array_update_77380[2] = add_77288 == 32'h0000_0002 ? add_77378 : array_index_77372[2];
  assign array_update_77380[3] = add_77288 == 32'h0000_0003 ? add_77378 : array_index_77372[3];
  assign array_update_77380[4] = add_77288 == 32'h0000_0004 ? add_77378 : array_index_77372[4];
  assign array_update_77380[5] = add_77288 == 32'h0000_0005 ? add_77378 : array_index_77372[5];
  assign array_update_77380[6] = add_77288 == 32'h0000_0006 ? add_77378 : array_index_77372[6];
  assign array_update_77380[7] = add_77288 == 32'h0000_0007 ? add_77378 : array_index_77372[7];
  assign array_update_77380[8] = add_77288 == 32'h0000_0008 ? add_77378 : array_index_77372[8];
  assign array_update_77380[9] = add_77288 == 32'h0000_0009 ? add_77378 : array_index_77372[9];
  assign add_77381 = add_77368 + 32'h0000_0001;
  assign array_update_77382[0] = add_76070 == 32'h0000_0000 ? array_update_77380 : array_update_77369[0];
  assign array_update_77382[1] = add_76070 == 32'h0000_0001 ? array_update_77380 : array_update_77369[1];
  assign array_update_77382[2] = add_76070 == 32'h0000_0002 ? array_update_77380 : array_update_77369[2];
  assign array_update_77382[3] = add_76070 == 32'h0000_0003 ? array_update_77380 : array_update_77369[3];
  assign array_update_77382[4] = add_76070 == 32'h0000_0004 ? array_update_77380 : array_update_77369[4];
  assign array_update_77382[5] = add_76070 == 32'h0000_0005 ? array_update_77380 : array_update_77369[5];
  assign array_update_77382[6] = add_76070 == 32'h0000_0006 ? array_update_77380 : array_update_77369[6];
  assign array_update_77382[7] = add_76070 == 32'h0000_0007 ? array_update_77380 : array_update_77369[7];
  assign array_update_77382[8] = add_76070 == 32'h0000_0008 ? array_update_77380 : array_update_77369[8];
  assign array_update_77382[9] = add_76070 == 32'h0000_0009 ? array_update_77380 : array_update_77369[9];
  assign array_index_77384 = array_update_72021[add_77381 > 32'h0000_0009 ? 4'h9 : add_77381[3:0]];
  assign array_index_77385 = array_update_77382[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_77389 = smul32b_32b_x_32b(array_index_76077[add_77381 > 32'h0000_0009 ? 4'h9 : add_77381[3:0]], array_index_77384[add_77288 > 32'h0000_0009 ? 4'h9 : add_77288[3:0]]);
  assign add_77391 = array_index_77385[add_77288 > 32'h0000_0009 ? 4'h9 : add_77288[3:0]] + smul_77389;
  assign array_update_77393[0] = add_77288 == 32'h0000_0000 ? add_77391 : array_index_77385[0];
  assign array_update_77393[1] = add_77288 == 32'h0000_0001 ? add_77391 : array_index_77385[1];
  assign array_update_77393[2] = add_77288 == 32'h0000_0002 ? add_77391 : array_index_77385[2];
  assign array_update_77393[3] = add_77288 == 32'h0000_0003 ? add_77391 : array_index_77385[3];
  assign array_update_77393[4] = add_77288 == 32'h0000_0004 ? add_77391 : array_index_77385[4];
  assign array_update_77393[5] = add_77288 == 32'h0000_0005 ? add_77391 : array_index_77385[5];
  assign array_update_77393[6] = add_77288 == 32'h0000_0006 ? add_77391 : array_index_77385[6];
  assign array_update_77393[7] = add_77288 == 32'h0000_0007 ? add_77391 : array_index_77385[7];
  assign array_update_77393[8] = add_77288 == 32'h0000_0008 ? add_77391 : array_index_77385[8];
  assign array_update_77393[9] = add_77288 == 32'h0000_0009 ? add_77391 : array_index_77385[9];
  assign add_77394 = add_77381 + 32'h0000_0001;
  assign array_update_77395[0] = add_76070 == 32'h0000_0000 ? array_update_77393 : array_update_77382[0];
  assign array_update_77395[1] = add_76070 == 32'h0000_0001 ? array_update_77393 : array_update_77382[1];
  assign array_update_77395[2] = add_76070 == 32'h0000_0002 ? array_update_77393 : array_update_77382[2];
  assign array_update_77395[3] = add_76070 == 32'h0000_0003 ? array_update_77393 : array_update_77382[3];
  assign array_update_77395[4] = add_76070 == 32'h0000_0004 ? array_update_77393 : array_update_77382[4];
  assign array_update_77395[5] = add_76070 == 32'h0000_0005 ? array_update_77393 : array_update_77382[5];
  assign array_update_77395[6] = add_76070 == 32'h0000_0006 ? array_update_77393 : array_update_77382[6];
  assign array_update_77395[7] = add_76070 == 32'h0000_0007 ? array_update_77393 : array_update_77382[7];
  assign array_update_77395[8] = add_76070 == 32'h0000_0008 ? array_update_77393 : array_update_77382[8];
  assign array_update_77395[9] = add_76070 == 32'h0000_0009 ? array_update_77393 : array_update_77382[9];
  assign array_index_77397 = array_update_72021[add_77394 > 32'h0000_0009 ? 4'h9 : add_77394[3:0]];
  assign array_index_77398 = array_update_77395[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_77402 = smul32b_32b_x_32b(array_index_76077[add_77394 > 32'h0000_0009 ? 4'h9 : add_77394[3:0]], array_index_77397[add_77288 > 32'h0000_0009 ? 4'h9 : add_77288[3:0]]);
  assign add_77404 = array_index_77398[add_77288 > 32'h0000_0009 ? 4'h9 : add_77288[3:0]] + smul_77402;
  assign array_update_77406[0] = add_77288 == 32'h0000_0000 ? add_77404 : array_index_77398[0];
  assign array_update_77406[1] = add_77288 == 32'h0000_0001 ? add_77404 : array_index_77398[1];
  assign array_update_77406[2] = add_77288 == 32'h0000_0002 ? add_77404 : array_index_77398[2];
  assign array_update_77406[3] = add_77288 == 32'h0000_0003 ? add_77404 : array_index_77398[3];
  assign array_update_77406[4] = add_77288 == 32'h0000_0004 ? add_77404 : array_index_77398[4];
  assign array_update_77406[5] = add_77288 == 32'h0000_0005 ? add_77404 : array_index_77398[5];
  assign array_update_77406[6] = add_77288 == 32'h0000_0006 ? add_77404 : array_index_77398[6];
  assign array_update_77406[7] = add_77288 == 32'h0000_0007 ? add_77404 : array_index_77398[7];
  assign array_update_77406[8] = add_77288 == 32'h0000_0008 ? add_77404 : array_index_77398[8];
  assign array_update_77406[9] = add_77288 == 32'h0000_0009 ? add_77404 : array_index_77398[9];
  assign add_77407 = add_77394 + 32'h0000_0001;
  assign array_update_77408[0] = add_76070 == 32'h0000_0000 ? array_update_77406 : array_update_77395[0];
  assign array_update_77408[1] = add_76070 == 32'h0000_0001 ? array_update_77406 : array_update_77395[1];
  assign array_update_77408[2] = add_76070 == 32'h0000_0002 ? array_update_77406 : array_update_77395[2];
  assign array_update_77408[3] = add_76070 == 32'h0000_0003 ? array_update_77406 : array_update_77395[3];
  assign array_update_77408[4] = add_76070 == 32'h0000_0004 ? array_update_77406 : array_update_77395[4];
  assign array_update_77408[5] = add_76070 == 32'h0000_0005 ? array_update_77406 : array_update_77395[5];
  assign array_update_77408[6] = add_76070 == 32'h0000_0006 ? array_update_77406 : array_update_77395[6];
  assign array_update_77408[7] = add_76070 == 32'h0000_0007 ? array_update_77406 : array_update_77395[7];
  assign array_update_77408[8] = add_76070 == 32'h0000_0008 ? array_update_77406 : array_update_77395[8];
  assign array_update_77408[9] = add_76070 == 32'h0000_0009 ? array_update_77406 : array_update_77395[9];
  assign array_index_77410 = array_update_72021[add_77407 > 32'h0000_0009 ? 4'h9 : add_77407[3:0]];
  assign array_index_77411 = array_update_77408[add_76070 > 32'h0000_0009 ? 4'h9 : add_76070[3:0]];
  assign smul_77415 = smul32b_32b_x_32b(array_index_76077[add_77407 > 32'h0000_0009 ? 4'h9 : add_77407[3:0]], array_index_77410[add_77288 > 32'h0000_0009 ? 4'h9 : add_77288[3:0]]);
  assign add_77417 = array_index_77411[add_77288 > 32'h0000_0009 ? 4'h9 : add_77288[3:0]] + smul_77415;
  assign array_update_77418[0] = add_77288 == 32'h0000_0000 ? add_77417 : array_index_77411[0];
  assign array_update_77418[1] = add_77288 == 32'h0000_0001 ? add_77417 : array_index_77411[1];
  assign array_update_77418[2] = add_77288 == 32'h0000_0002 ? add_77417 : array_index_77411[2];
  assign array_update_77418[3] = add_77288 == 32'h0000_0003 ? add_77417 : array_index_77411[3];
  assign array_update_77418[4] = add_77288 == 32'h0000_0004 ? add_77417 : array_index_77411[4];
  assign array_update_77418[5] = add_77288 == 32'h0000_0005 ? add_77417 : array_index_77411[5];
  assign array_update_77418[6] = add_77288 == 32'h0000_0006 ? add_77417 : array_index_77411[6];
  assign array_update_77418[7] = add_77288 == 32'h0000_0007 ? add_77417 : array_index_77411[7];
  assign array_update_77418[8] = add_77288 == 32'h0000_0008 ? add_77417 : array_index_77411[8];
  assign array_update_77418[9] = add_77288 == 32'h0000_0009 ? add_77417 : array_index_77411[9];
  assign array_update_77420[0] = add_76070 == 32'h0000_0000 ? array_update_77418 : array_update_77408[0];
  assign array_update_77420[1] = add_76070 == 32'h0000_0001 ? array_update_77418 : array_update_77408[1];
  assign array_update_77420[2] = add_76070 == 32'h0000_0002 ? array_update_77418 : array_update_77408[2];
  assign array_update_77420[3] = add_76070 == 32'h0000_0003 ? array_update_77418 : array_update_77408[3];
  assign array_update_77420[4] = add_76070 == 32'h0000_0004 ? array_update_77418 : array_update_77408[4];
  assign array_update_77420[5] = add_76070 == 32'h0000_0005 ? array_update_77418 : array_update_77408[5];
  assign array_update_77420[6] = add_76070 == 32'h0000_0006 ? array_update_77418 : array_update_77408[6];
  assign array_update_77420[7] = add_76070 == 32'h0000_0007 ? array_update_77418 : array_update_77408[7];
  assign array_update_77420[8] = add_76070 == 32'h0000_0008 ? array_update_77418 : array_update_77408[8];
  assign array_update_77420[9] = add_76070 == 32'h0000_0009 ? array_update_77418 : array_update_77408[9];
  assign add_77421 = add_76070 + 32'h0000_0001;
  assign array_index_77422 = array_update_77420[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign literal_77424 = 32'h0000_0000;
  assign array_update_77425[0] = literal_77424 == 32'h0000_0000 ? 32'h0000_0000 : array_index_77422[0];
  assign array_update_77425[1] = literal_77424 == 32'h0000_0001 ? 32'h0000_0000 : array_index_77422[1];
  assign array_update_77425[2] = literal_77424 == 32'h0000_0002 ? 32'h0000_0000 : array_index_77422[2];
  assign array_update_77425[3] = literal_77424 == 32'h0000_0003 ? 32'h0000_0000 : array_index_77422[3];
  assign array_update_77425[4] = literal_77424 == 32'h0000_0004 ? 32'h0000_0000 : array_index_77422[4];
  assign array_update_77425[5] = literal_77424 == 32'h0000_0005 ? 32'h0000_0000 : array_index_77422[5];
  assign array_update_77425[6] = literal_77424 == 32'h0000_0006 ? 32'h0000_0000 : array_index_77422[6];
  assign array_update_77425[7] = literal_77424 == 32'h0000_0007 ? 32'h0000_0000 : array_index_77422[7];
  assign array_update_77425[8] = literal_77424 == 32'h0000_0008 ? 32'h0000_0000 : array_index_77422[8];
  assign array_update_77425[9] = literal_77424 == 32'h0000_0009 ? 32'h0000_0000 : array_index_77422[9];
  assign literal_77426 = 32'h0000_0000;
  assign array_update_77427[0] = add_77421 == 32'h0000_0000 ? array_update_77425 : array_update_77420[0];
  assign array_update_77427[1] = add_77421 == 32'h0000_0001 ? array_update_77425 : array_update_77420[1];
  assign array_update_77427[2] = add_77421 == 32'h0000_0002 ? array_update_77425 : array_update_77420[2];
  assign array_update_77427[3] = add_77421 == 32'h0000_0003 ? array_update_77425 : array_update_77420[3];
  assign array_update_77427[4] = add_77421 == 32'h0000_0004 ? array_update_77425 : array_update_77420[4];
  assign array_update_77427[5] = add_77421 == 32'h0000_0005 ? array_update_77425 : array_update_77420[5];
  assign array_update_77427[6] = add_77421 == 32'h0000_0006 ? array_update_77425 : array_update_77420[6];
  assign array_update_77427[7] = add_77421 == 32'h0000_0007 ? array_update_77425 : array_update_77420[7];
  assign array_update_77427[8] = add_77421 == 32'h0000_0008 ? array_update_77425 : array_update_77420[8];
  assign array_update_77427[9] = add_77421 == 32'h0000_0009 ? array_update_77425 : array_update_77420[9];
  assign array_index_77428 = array_update_72020[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign array_index_77429 = array_update_72021[literal_77426 > 32'h0000_0009 ? 4'h9 : literal_77426[3:0]];
  assign array_index_77430 = array_update_77427[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_77434 = smul32b_32b_x_32b(array_index_77428[literal_77426 > 32'h0000_0009 ? 4'h9 : literal_77426[3:0]], array_index_77429[literal_77424 > 32'h0000_0009 ? 4'h9 : literal_77424[3:0]]);
  assign add_77436 = array_index_77430[literal_77424 > 32'h0000_0009 ? 4'h9 : literal_77424[3:0]] + smul_77434;
  assign array_update_77438[0] = literal_77424 == 32'h0000_0000 ? add_77436 : array_index_77430[0];
  assign array_update_77438[1] = literal_77424 == 32'h0000_0001 ? add_77436 : array_index_77430[1];
  assign array_update_77438[2] = literal_77424 == 32'h0000_0002 ? add_77436 : array_index_77430[2];
  assign array_update_77438[3] = literal_77424 == 32'h0000_0003 ? add_77436 : array_index_77430[3];
  assign array_update_77438[4] = literal_77424 == 32'h0000_0004 ? add_77436 : array_index_77430[4];
  assign array_update_77438[5] = literal_77424 == 32'h0000_0005 ? add_77436 : array_index_77430[5];
  assign array_update_77438[6] = literal_77424 == 32'h0000_0006 ? add_77436 : array_index_77430[6];
  assign array_update_77438[7] = literal_77424 == 32'h0000_0007 ? add_77436 : array_index_77430[7];
  assign array_update_77438[8] = literal_77424 == 32'h0000_0008 ? add_77436 : array_index_77430[8];
  assign array_update_77438[9] = literal_77424 == 32'h0000_0009 ? add_77436 : array_index_77430[9];
  assign add_77439 = literal_77426 + 32'h0000_0001;
  assign array_update_77440[0] = add_77421 == 32'h0000_0000 ? array_update_77438 : array_update_77427[0];
  assign array_update_77440[1] = add_77421 == 32'h0000_0001 ? array_update_77438 : array_update_77427[1];
  assign array_update_77440[2] = add_77421 == 32'h0000_0002 ? array_update_77438 : array_update_77427[2];
  assign array_update_77440[3] = add_77421 == 32'h0000_0003 ? array_update_77438 : array_update_77427[3];
  assign array_update_77440[4] = add_77421 == 32'h0000_0004 ? array_update_77438 : array_update_77427[4];
  assign array_update_77440[5] = add_77421 == 32'h0000_0005 ? array_update_77438 : array_update_77427[5];
  assign array_update_77440[6] = add_77421 == 32'h0000_0006 ? array_update_77438 : array_update_77427[6];
  assign array_update_77440[7] = add_77421 == 32'h0000_0007 ? array_update_77438 : array_update_77427[7];
  assign array_update_77440[8] = add_77421 == 32'h0000_0008 ? array_update_77438 : array_update_77427[8];
  assign array_update_77440[9] = add_77421 == 32'h0000_0009 ? array_update_77438 : array_update_77427[9];
  assign array_index_77442 = array_update_72021[add_77439 > 32'h0000_0009 ? 4'h9 : add_77439[3:0]];
  assign array_index_77443 = array_update_77440[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_77447 = smul32b_32b_x_32b(array_index_77428[add_77439 > 32'h0000_0009 ? 4'h9 : add_77439[3:0]], array_index_77442[literal_77424 > 32'h0000_0009 ? 4'h9 : literal_77424[3:0]]);
  assign add_77449 = array_index_77443[literal_77424 > 32'h0000_0009 ? 4'h9 : literal_77424[3:0]] + smul_77447;
  assign array_update_77451[0] = literal_77424 == 32'h0000_0000 ? add_77449 : array_index_77443[0];
  assign array_update_77451[1] = literal_77424 == 32'h0000_0001 ? add_77449 : array_index_77443[1];
  assign array_update_77451[2] = literal_77424 == 32'h0000_0002 ? add_77449 : array_index_77443[2];
  assign array_update_77451[3] = literal_77424 == 32'h0000_0003 ? add_77449 : array_index_77443[3];
  assign array_update_77451[4] = literal_77424 == 32'h0000_0004 ? add_77449 : array_index_77443[4];
  assign array_update_77451[5] = literal_77424 == 32'h0000_0005 ? add_77449 : array_index_77443[5];
  assign array_update_77451[6] = literal_77424 == 32'h0000_0006 ? add_77449 : array_index_77443[6];
  assign array_update_77451[7] = literal_77424 == 32'h0000_0007 ? add_77449 : array_index_77443[7];
  assign array_update_77451[8] = literal_77424 == 32'h0000_0008 ? add_77449 : array_index_77443[8];
  assign array_update_77451[9] = literal_77424 == 32'h0000_0009 ? add_77449 : array_index_77443[9];
  assign add_77452 = add_77439 + 32'h0000_0001;
  assign array_update_77453[0] = add_77421 == 32'h0000_0000 ? array_update_77451 : array_update_77440[0];
  assign array_update_77453[1] = add_77421 == 32'h0000_0001 ? array_update_77451 : array_update_77440[1];
  assign array_update_77453[2] = add_77421 == 32'h0000_0002 ? array_update_77451 : array_update_77440[2];
  assign array_update_77453[3] = add_77421 == 32'h0000_0003 ? array_update_77451 : array_update_77440[3];
  assign array_update_77453[4] = add_77421 == 32'h0000_0004 ? array_update_77451 : array_update_77440[4];
  assign array_update_77453[5] = add_77421 == 32'h0000_0005 ? array_update_77451 : array_update_77440[5];
  assign array_update_77453[6] = add_77421 == 32'h0000_0006 ? array_update_77451 : array_update_77440[6];
  assign array_update_77453[7] = add_77421 == 32'h0000_0007 ? array_update_77451 : array_update_77440[7];
  assign array_update_77453[8] = add_77421 == 32'h0000_0008 ? array_update_77451 : array_update_77440[8];
  assign array_update_77453[9] = add_77421 == 32'h0000_0009 ? array_update_77451 : array_update_77440[9];
  assign array_index_77455 = array_update_72021[add_77452 > 32'h0000_0009 ? 4'h9 : add_77452[3:0]];
  assign array_index_77456 = array_update_77453[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_77460 = smul32b_32b_x_32b(array_index_77428[add_77452 > 32'h0000_0009 ? 4'h9 : add_77452[3:0]], array_index_77455[literal_77424 > 32'h0000_0009 ? 4'h9 : literal_77424[3:0]]);
  assign add_77462 = array_index_77456[literal_77424 > 32'h0000_0009 ? 4'h9 : literal_77424[3:0]] + smul_77460;
  assign array_update_77464[0] = literal_77424 == 32'h0000_0000 ? add_77462 : array_index_77456[0];
  assign array_update_77464[1] = literal_77424 == 32'h0000_0001 ? add_77462 : array_index_77456[1];
  assign array_update_77464[2] = literal_77424 == 32'h0000_0002 ? add_77462 : array_index_77456[2];
  assign array_update_77464[3] = literal_77424 == 32'h0000_0003 ? add_77462 : array_index_77456[3];
  assign array_update_77464[4] = literal_77424 == 32'h0000_0004 ? add_77462 : array_index_77456[4];
  assign array_update_77464[5] = literal_77424 == 32'h0000_0005 ? add_77462 : array_index_77456[5];
  assign array_update_77464[6] = literal_77424 == 32'h0000_0006 ? add_77462 : array_index_77456[6];
  assign array_update_77464[7] = literal_77424 == 32'h0000_0007 ? add_77462 : array_index_77456[7];
  assign array_update_77464[8] = literal_77424 == 32'h0000_0008 ? add_77462 : array_index_77456[8];
  assign array_update_77464[9] = literal_77424 == 32'h0000_0009 ? add_77462 : array_index_77456[9];
  assign add_77465 = add_77452 + 32'h0000_0001;
  assign array_update_77466[0] = add_77421 == 32'h0000_0000 ? array_update_77464 : array_update_77453[0];
  assign array_update_77466[1] = add_77421 == 32'h0000_0001 ? array_update_77464 : array_update_77453[1];
  assign array_update_77466[2] = add_77421 == 32'h0000_0002 ? array_update_77464 : array_update_77453[2];
  assign array_update_77466[3] = add_77421 == 32'h0000_0003 ? array_update_77464 : array_update_77453[3];
  assign array_update_77466[4] = add_77421 == 32'h0000_0004 ? array_update_77464 : array_update_77453[4];
  assign array_update_77466[5] = add_77421 == 32'h0000_0005 ? array_update_77464 : array_update_77453[5];
  assign array_update_77466[6] = add_77421 == 32'h0000_0006 ? array_update_77464 : array_update_77453[6];
  assign array_update_77466[7] = add_77421 == 32'h0000_0007 ? array_update_77464 : array_update_77453[7];
  assign array_update_77466[8] = add_77421 == 32'h0000_0008 ? array_update_77464 : array_update_77453[8];
  assign array_update_77466[9] = add_77421 == 32'h0000_0009 ? array_update_77464 : array_update_77453[9];
  assign array_index_77468 = array_update_72021[add_77465 > 32'h0000_0009 ? 4'h9 : add_77465[3:0]];
  assign array_index_77469 = array_update_77466[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_77473 = smul32b_32b_x_32b(array_index_77428[add_77465 > 32'h0000_0009 ? 4'h9 : add_77465[3:0]], array_index_77468[literal_77424 > 32'h0000_0009 ? 4'h9 : literal_77424[3:0]]);
  assign add_77475 = array_index_77469[literal_77424 > 32'h0000_0009 ? 4'h9 : literal_77424[3:0]] + smul_77473;
  assign array_update_77477[0] = literal_77424 == 32'h0000_0000 ? add_77475 : array_index_77469[0];
  assign array_update_77477[1] = literal_77424 == 32'h0000_0001 ? add_77475 : array_index_77469[1];
  assign array_update_77477[2] = literal_77424 == 32'h0000_0002 ? add_77475 : array_index_77469[2];
  assign array_update_77477[3] = literal_77424 == 32'h0000_0003 ? add_77475 : array_index_77469[3];
  assign array_update_77477[4] = literal_77424 == 32'h0000_0004 ? add_77475 : array_index_77469[4];
  assign array_update_77477[5] = literal_77424 == 32'h0000_0005 ? add_77475 : array_index_77469[5];
  assign array_update_77477[6] = literal_77424 == 32'h0000_0006 ? add_77475 : array_index_77469[6];
  assign array_update_77477[7] = literal_77424 == 32'h0000_0007 ? add_77475 : array_index_77469[7];
  assign array_update_77477[8] = literal_77424 == 32'h0000_0008 ? add_77475 : array_index_77469[8];
  assign array_update_77477[9] = literal_77424 == 32'h0000_0009 ? add_77475 : array_index_77469[9];
  assign add_77478 = add_77465 + 32'h0000_0001;
  assign array_update_77479[0] = add_77421 == 32'h0000_0000 ? array_update_77477 : array_update_77466[0];
  assign array_update_77479[1] = add_77421 == 32'h0000_0001 ? array_update_77477 : array_update_77466[1];
  assign array_update_77479[2] = add_77421 == 32'h0000_0002 ? array_update_77477 : array_update_77466[2];
  assign array_update_77479[3] = add_77421 == 32'h0000_0003 ? array_update_77477 : array_update_77466[3];
  assign array_update_77479[4] = add_77421 == 32'h0000_0004 ? array_update_77477 : array_update_77466[4];
  assign array_update_77479[5] = add_77421 == 32'h0000_0005 ? array_update_77477 : array_update_77466[5];
  assign array_update_77479[6] = add_77421 == 32'h0000_0006 ? array_update_77477 : array_update_77466[6];
  assign array_update_77479[7] = add_77421 == 32'h0000_0007 ? array_update_77477 : array_update_77466[7];
  assign array_update_77479[8] = add_77421 == 32'h0000_0008 ? array_update_77477 : array_update_77466[8];
  assign array_update_77479[9] = add_77421 == 32'h0000_0009 ? array_update_77477 : array_update_77466[9];
  assign array_index_77481 = array_update_72021[add_77478 > 32'h0000_0009 ? 4'h9 : add_77478[3:0]];
  assign array_index_77482 = array_update_77479[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_77486 = smul32b_32b_x_32b(array_index_77428[add_77478 > 32'h0000_0009 ? 4'h9 : add_77478[3:0]], array_index_77481[literal_77424 > 32'h0000_0009 ? 4'h9 : literal_77424[3:0]]);
  assign add_77488 = array_index_77482[literal_77424 > 32'h0000_0009 ? 4'h9 : literal_77424[3:0]] + smul_77486;
  assign array_update_77490[0] = literal_77424 == 32'h0000_0000 ? add_77488 : array_index_77482[0];
  assign array_update_77490[1] = literal_77424 == 32'h0000_0001 ? add_77488 : array_index_77482[1];
  assign array_update_77490[2] = literal_77424 == 32'h0000_0002 ? add_77488 : array_index_77482[2];
  assign array_update_77490[3] = literal_77424 == 32'h0000_0003 ? add_77488 : array_index_77482[3];
  assign array_update_77490[4] = literal_77424 == 32'h0000_0004 ? add_77488 : array_index_77482[4];
  assign array_update_77490[5] = literal_77424 == 32'h0000_0005 ? add_77488 : array_index_77482[5];
  assign array_update_77490[6] = literal_77424 == 32'h0000_0006 ? add_77488 : array_index_77482[6];
  assign array_update_77490[7] = literal_77424 == 32'h0000_0007 ? add_77488 : array_index_77482[7];
  assign array_update_77490[8] = literal_77424 == 32'h0000_0008 ? add_77488 : array_index_77482[8];
  assign array_update_77490[9] = literal_77424 == 32'h0000_0009 ? add_77488 : array_index_77482[9];
  assign add_77491 = add_77478 + 32'h0000_0001;
  assign array_update_77492[0] = add_77421 == 32'h0000_0000 ? array_update_77490 : array_update_77479[0];
  assign array_update_77492[1] = add_77421 == 32'h0000_0001 ? array_update_77490 : array_update_77479[1];
  assign array_update_77492[2] = add_77421 == 32'h0000_0002 ? array_update_77490 : array_update_77479[2];
  assign array_update_77492[3] = add_77421 == 32'h0000_0003 ? array_update_77490 : array_update_77479[3];
  assign array_update_77492[4] = add_77421 == 32'h0000_0004 ? array_update_77490 : array_update_77479[4];
  assign array_update_77492[5] = add_77421 == 32'h0000_0005 ? array_update_77490 : array_update_77479[5];
  assign array_update_77492[6] = add_77421 == 32'h0000_0006 ? array_update_77490 : array_update_77479[6];
  assign array_update_77492[7] = add_77421 == 32'h0000_0007 ? array_update_77490 : array_update_77479[7];
  assign array_update_77492[8] = add_77421 == 32'h0000_0008 ? array_update_77490 : array_update_77479[8];
  assign array_update_77492[9] = add_77421 == 32'h0000_0009 ? array_update_77490 : array_update_77479[9];
  assign array_index_77494 = array_update_72021[add_77491 > 32'h0000_0009 ? 4'h9 : add_77491[3:0]];
  assign array_index_77495 = array_update_77492[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_77499 = smul32b_32b_x_32b(array_index_77428[add_77491 > 32'h0000_0009 ? 4'h9 : add_77491[3:0]], array_index_77494[literal_77424 > 32'h0000_0009 ? 4'h9 : literal_77424[3:0]]);
  assign add_77501 = array_index_77495[literal_77424 > 32'h0000_0009 ? 4'h9 : literal_77424[3:0]] + smul_77499;
  assign array_update_77503[0] = literal_77424 == 32'h0000_0000 ? add_77501 : array_index_77495[0];
  assign array_update_77503[1] = literal_77424 == 32'h0000_0001 ? add_77501 : array_index_77495[1];
  assign array_update_77503[2] = literal_77424 == 32'h0000_0002 ? add_77501 : array_index_77495[2];
  assign array_update_77503[3] = literal_77424 == 32'h0000_0003 ? add_77501 : array_index_77495[3];
  assign array_update_77503[4] = literal_77424 == 32'h0000_0004 ? add_77501 : array_index_77495[4];
  assign array_update_77503[5] = literal_77424 == 32'h0000_0005 ? add_77501 : array_index_77495[5];
  assign array_update_77503[6] = literal_77424 == 32'h0000_0006 ? add_77501 : array_index_77495[6];
  assign array_update_77503[7] = literal_77424 == 32'h0000_0007 ? add_77501 : array_index_77495[7];
  assign array_update_77503[8] = literal_77424 == 32'h0000_0008 ? add_77501 : array_index_77495[8];
  assign array_update_77503[9] = literal_77424 == 32'h0000_0009 ? add_77501 : array_index_77495[9];
  assign add_77504 = add_77491 + 32'h0000_0001;
  assign array_update_77505[0] = add_77421 == 32'h0000_0000 ? array_update_77503 : array_update_77492[0];
  assign array_update_77505[1] = add_77421 == 32'h0000_0001 ? array_update_77503 : array_update_77492[1];
  assign array_update_77505[2] = add_77421 == 32'h0000_0002 ? array_update_77503 : array_update_77492[2];
  assign array_update_77505[3] = add_77421 == 32'h0000_0003 ? array_update_77503 : array_update_77492[3];
  assign array_update_77505[4] = add_77421 == 32'h0000_0004 ? array_update_77503 : array_update_77492[4];
  assign array_update_77505[5] = add_77421 == 32'h0000_0005 ? array_update_77503 : array_update_77492[5];
  assign array_update_77505[6] = add_77421 == 32'h0000_0006 ? array_update_77503 : array_update_77492[6];
  assign array_update_77505[7] = add_77421 == 32'h0000_0007 ? array_update_77503 : array_update_77492[7];
  assign array_update_77505[8] = add_77421 == 32'h0000_0008 ? array_update_77503 : array_update_77492[8];
  assign array_update_77505[9] = add_77421 == 32'h0000_0009 ? array_update_77503 : array_update_77492[9];
  assign array_index_77507 = array_update_72021[add_77504 > 32'h0000_0009 ? 4'h9 : add_77504[3:0]];
  assign array_index_77508 = array_update_77505[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_77512 = smul32b_32b_x_32b(array_index_77428[add_77504 > 32'h0000_0009 ? 4'h9 : add_77504[3:0]], array_index_77507[literal_77424 > 32'h0000_0009 ? 4'h9 : literal_77424[3:0]]);
  assign add_77514 = array_index_77508[literal_77424 > 32'h0000_0009 ? 4'h9 : literal_77424[3:0]] + smul_77512;
  assign array_update_77516[0] = literal_77424 == 32'h0000_0000 ? add_77514 : array_index_77508[0];
  assign array_update_77516[1] = literal_77424 == 32'h0000_0001 ? add_77514 : array_index_77508[1];
  assign array_update_77516[2] = literal_77424 == 32'h0000_0002 ? add_77514 : array_index_77508[2];
  assign array_update_77516[3] = literal_77424 == 32'h0000_0003 ? add_77514 : array_index_77508[3];
  assign array_update_77516[4] = literal_77424 == 32'h0000_0004 ? add_77514 : array_index_77508[4];
  assign array_update_77516[5] = literal_77424 == 32'h0000_0005 ? add_77514 : array_index_77508[5];
  assign array_update_77516[6] = literal_77424 == 32'h0000_0006 ? add_77514 : array_index_77508[6];
  assign array_update_77516[7] = literal_77424 == 32'h0000_0007 ? add_77514 : array_index_77508[7];
  assign array_update_77516[8] = literal_77424 == 32'h0000_0008 ? add_77514 : array_index_77508[8];
  assign array_update_77516[9] = literal_77424 == 32'h0000_0009 ? add_77514 : array_index_77508[9];
  assign add_77517 = add_77504 + 32'h0000_0001;
  assign array_update_77518[0] = add_77421 == 32'h0000_0000 ? array_update_77516 : array_update_77505[0];
  assign array_update_77518[1] = add_77421 == 32'h0000_0001 ? array_update_77516 : array_update_77505[1];
  assign array_update_77518[2] = add_77421 == 32'h0000_0002 ? array_update_77516 : array_update_77505[2];
  assign array_update_77518[3] = add_77421 == 32'h0000_0003 ? array_update_77516 : array_update_77505[3];
  assign array_update_77518[4] = add_77421 == 32'h0000_0004 ? array_update_77516 : array_update_77505[4];
  assign array_update_77518[5] = add_77421 == 32'h0000_0005 ? array_update_77516 : array_update_77505[5];
  assign array_update_77518[6] = add_77421 == 32'h0000_0006 ? array_update_77516 : array_update_77505[6];
  assign array_update_77518[7] = add_77421 == 32'h0000_0007 ? array_update_77516 : array_update_77505[7];
  assign array_update_77518[8] = add_77421 == 32'h0000_0008 ? array_update_77516 : array_update_77505[8];
  assign array_update_77518[9] = add_77421 == 32'h0000_0009 ? array_update_77516 : array_update_77505[9];
  assign array_index_77520 = array_update_72021[add_77517 > 32'h0000_0009 ? 4'h9 : add_77517[3:0]];
  assign array_index_77521 = array_update_77518[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_77525 = smul32b_32b_x_32b(array_index_77428[add_77517 > 32'h0000_0009 ? 4'h9 : add_77517[3:0]], array_index_77520[literal_77424 > 32'h0000_0009 ? 4'h9 : literal_77424[3:0]]);
  assign add_77527 = array_index_77521[literal_77424 > 32'h0000_0009 ? 4'h9 : literal_77424[3:0]] + smul_77525;
  assign array_update_77529[0] = literal_77424 == 32'h0000_0000 ? add_77527 : array_index_77521[0];
  assign array_update_77529[1] = literal_77424 == 32'h0000_0001 ? add_77527 : array_index_77521[1];
  assign array_update_77529[2] = literal_77424 == 32'h0000_0002 ? add_77527 : array_index_77521[2];
  assign array_update_77529[3] = literal_77424 == 32'h0000_0003 ? add_77527 : array_index_77521[3];
  assign array_update_77529[4] = literal_77424 == 32'h0000_0004 ? add_77527 : array_index_77521[4];
  assign array_update_77529[5] = literal_77424 == 32'h0000_0005 ? add_77527 : array_index_77521[5];
  assign array_update_77529[6] = literal_77424 == 32'h0000_0006 ? add_77527 : array_index_77521[6];
  assign array_update_77529[7] = literal_77424 == 32'h0000_0007 ? add_77527 : array_index_77521[7];
  assign array_update_77529[8] = literal_77424 == 32'h0000_0008 ? add_77527 : array_index_77521[8];
  assign array_update_77529[9] = literal_77424 == 32'h0000_0009 ? add_77527 : array_index_77521[9];
  assign add_77530 = add_77517 + 32'h0000_0001;
  assign array_update_77531[0] = add_77421 == 32'h0000_0000 ? array_update_77529 : array_update_77518[0];
  assign array_update_77531[1] = add_77421 == 32'h0000_0001 ? array_update_77529 : array_update_77518[1];
  assign array_update_77531[2] = add_77421 == 32'h0000_0002 ? array_update_77529 : array_update_77518[2];
  assign array_update_77531[3] = add_77421 == 32'h0000_0003 ? array_update_77529 : array_update_77518[3];
  assign array_update_77531[4] = add_77421 == 32'h0000_0004 ? array_update_77529 : array_update_77518[4];
  assign array_update_77531[5] = add_77421 == 32'h0000_0005 ? array_update_77529 : array_update_77518[5];
  assign array_update_77531[6] = add_77421 == 32'h0000_0006 ? array_update_77529 : array_update_77518[6];
  assign array_update_77531[7] = add_77421 == 32'h0000_0007 ? array_update_77529 : array_update_77518[7];
  assign array_update_77531[8] = add_77421 == 32'h0000_0008 ? array_update_77529 : array_update_77518[8];
  assign array_update_77531[9] = add_77421 == 32'h0000_0009 ? array_update_77529 : array_update_77518[9];
  assign array_index_77533 = array_update_72021[add_77530 > 32'h0000_0009 ? 4'h9 : add_77530[3:0]];
  assign array_index_77534 = array_update_77531[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_77538 = smul32b_32b_x_32b(array_index_77428[add_77530 > 32'h0000_0009 ? 4'h9 : add_77530[3:0]], array_index_77533[literal_77424 > 32'h0000_0009 ? 4'h9 : literal_77424[3:0]]);
  assign add_77540 = array_index_77534[literal_77424 > 32'h0000_0009 ? 4'h9 : literal_77424[3:0]] + smul_77538;
  assign array_update_77542[0] = literal_77424 == 32'h0000_0000 ? add_77540 : array_index_77534[0];
  assign array_update_77542[1] = literal_77424 == 32'h0000_0001 ? add_77540 : array_index_77534[1];
  assign array_update_77542[2] = literal_77424 == 32'h0000_0002 ? add_77540 : array_index_77534[2];
  assign array_update_77542[3] = literal_77424 == 32'h0000_0003 ? add_77540 : array_index_77534[3];
  assign array_update_77542[4] = literal_77424 == 32'h0000_0004 ? add_77540 : array_index_77534[4];
  assign array_update_77542[5] = literal_77424 == 32'h0000_0005 ? add_77540 : array_index_77534[5];
  assign array_update_77542[6] = literal_77424 == 32'h0000_0006 ? add_77540 : array_index_77534[6];
  assign array_update_77542[7] = literal_77424 == 32'h0000_0007 ? add_77540 : array_index_77534[7];
  assign array_update_77542[8] = literal_77424 == 32'h0000_0008 ? add_77540 : array_index_77534[8];
  assign array_update_77542[9] = literal_77424 == 32'h0000_0009 ? add_77540 : array_index_77534[9];
  assign add_77543 = add_77530 + 32'h0000_0001;
  assign array_update_77544[0] = add_77421 == 32'h0000_0000 ? array_update_77542 : array_update_77531[0];
  assign array_update_77544[1] = add_77421 == 32'h0000_0001 ? array_update_77542 : array_update_77531[1];
  assign array_update_77544[2] = add_77421 == 32'h0000_0002 ? array_update_77542 : array_update_77531[2];
  assign array_update_77544[3] = add_77421 == 32'h0000_0003 ? array_update_77542 : array_update_77531[3];
  assign array_update_77544[4] = add_77421 == 32'h0000_0004 ? array_update_77542 : array_update_77531[4];
  assign array_update_77544[5] = add_77421 == 32'h0000_0005 ? array_update_77542 : array_update_77531[5];
  assign array_update_77544[6] = add_77421 == 32'h0000_0006 ? array_update_77542 : array_update_77531[6];
  assign array_update_77544[7] = add_77421 == 32'h0000_0007 ? array_update_77542 : array_update_77531[7];
  assign array_update_77544[8] = add_77421 == 32'h0000_0008 ? array_update_77542 : array_update_77531[8];
  assign array_update_77544[9] = add_77421 == 32'h0000_0009 ? array_update_77542 : array_update_77531[9];
  assign array_index_77546 = array_update_72021[add_77543 > 32'h0000_0009 ? 4'h9 : add_77543[3:0]];
  assign array_index_77547 = array_update_77544[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_77551 = smul32b_32b_x_32b(array_index_77428[add_77543 > 32'h0000_0009 ? 4'h9 : add_77543[3:0]], array_index_77546[literal_77424 > 32'h0000_0009 ? 4'h9 : literal_77424[3:0]]);
  assign add_77553 = array_index_77547[literal_77424 > 32'h0000_0009 ? 4'h9 : literal_77424[3:0]] + smul_77551;
  assign array_update_77554[0] = literal_77424 == 32'h0000_0000 ? add_77553 : array_index_77547[0];
  assign array_update_77554[1] = literal_77424 == 32'h0000_0001 ? add_77553 : array_index_77547[1];
  assign array_update_77554[2] = literal_77424 == 32'h0000_0002 ? add_77553 : array_index_77547[2];
  assign array_update_77554[3] = literal_77424 == 32'h0000_0003 ? add_77553 : array_index_77547[3];
  assign array_update_77554[4] = literal_77424 == 32'h0000_0004 ? add_77553 : array_index_77547[4];
  assign array_update_77554[5] = literal_77424 == 32'h0000_0005 ? add_77553 : array_index_77547[5];
  assign array_update_77554[6] = literal_77424 == 32'h0000_0006 ? add_77553 : array_index_77547[6];
  assign array_update_77554[7] = literal_77424 == 32'h0000_0007 ? add_77553 : array_index_77547[7];
  assign array_update_77554[8] = literal_77424 == 32'h0000_0008 ? add_77553 : array_index_77547[8];
  assign array_update_77554[9] = literal_77424 == 32'h0000_0009 ? add_77553 : array_index_77547[9];
  assign array_update_77555[0] = add_77421 == 32'h0000_0000 ? array_update_77554 : array_update_77544[0];
  assign array_update_77555[1] = add_77421 == 32'h0000_0001 ? array_update_77554 : array_update_77544[1];
  assign array_update_77555[2] = add_77421 == 32'h0000_0002 ? array_update_77554 : array_update_77544[2];
  assign array_update_77555[3] = add_77421 == 32'h0000_0003 ? array_update_77554 : array_update_77544[3];
  assign array_update_77555[4] = add_77421 == 32'h0000_0004 ? array_update_77554 : array_update_77544[4];
  assign array_update_77555[5] = add_77421 == 32'h0000_0005 ? array_update_77554 : array_update_77544[5];
  assign array_update_77555[6] = add_77421 == 32'h0000_0006 ? array_update_77554 : array_update_77544[6];
  assign array_update_77555[7] = add_77421 == 32'h0000_0007 ? array_update_77554 : array_update_77544[7];
  assign array_update_77555[8] = add_77421 == 32'h0000_0008 ? array_update_77554 : array_update_77544[8];
  assign array_update_77555[9] = add_77421 == 32'h0000_0009 ? array_update_77554 : array_update_77544[9];
  assign array_index_77557 = array_update_77555[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign add_77559 = literal_77424 + 32'h0000_0001;
  assign array_update_77560[0] = add_77559 == 32'h0000_0000 ? 32'h0000_0000 : array_index_77557[0];
  assign array_update_77560[1] = add_77559 == 32'h0000_0001 ? 32'h0000_0000 : array_index_77557[1];
  assign array_update_77560[2] = add_77559 == 32'h0000_0002 ? 32'h0000_0000 : array_index_77557[2];
  assign array_update_77560[3] = add_77559 == 32'h0000_0003 ? 32'h0000_0000 : array_index_77557[3];
  assign array_update_77560[4] = add_77559 == 32'h0000_0004 ? 32'h0000_0000 : array_index_77557[4];
  assign array_update_77560[5] = add_77559 == 32'h0000_0005 ? 32'h0000_0000 : array_index_77557[5];
  assign array_update_77560[6] = add_77559 == 32'h0000_0006 ? 32'h0000_0000 : array_index_77557[6];
  assign array_update_77560[7] = add_77559 == 32'h0000_0007 ? 32'h0000_0000 : array_index_77557[7];
  assign array_update_77560[8] = add_77559 == 32'h0000_0008 ? 32'h0000_0000 : array_index_77557[8];
  assign array_update_77560[9] = add_77559 == 32'h0000_0009 ? 32'h0000_0000 : array_index_77557[9];
  assign literal_77561 = 32'h0000_0000;
  assign array_update_77562[0] = add_77421 == 32'h0000_0000 ? array_update_77560 : array_update_77555[0];
  assign array_update_77562[1] = add_77421 == 32'h0000_0001 ? array_update_77560 : array_update_77555[1];
  assign array_update_77562[2] = add_77421 == 32'h0000_0002 ? array_update_77560 : array_update_77555[2];
  assign array_update_77562[3] = add_77421 == 32'h0000_0003 ? array_update_77560 : array_update_77555[3];
  assign array_update_77562[4] = add_77421 == 32'h0000_0004 ? array_update_77560 : array_update_77555[4];
  assign array_update_77562[5] = add_77421 == 32'h0000_0005 ? array_update_77560 : array_update_77555[5];
  assign array_update_77562[6] = add_77421 == 32'h0000_0006 ? array_update_77560 : array_update_77555[6];
  assign array_update_77562[7] = add_77421 == 32'h0000_0007 ? array_update_77560 : array_update_77555[7];
  assign array_update_77562[8] = add_77421 == 32'h0000_0008 ? array_update_77560 : array_update_77555[8];
  assign array_update_77562[9] = add_77421 == 32'h0000_0009 ? array_update_77560 : array_update_77555[9];
  assign array_index_77564 = array_update_72021[literal_77561 > 32'h0000_0009 ? 4'h9 : literal_77561[3:0]];
  assign array_index_77565 = array_update_77562[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_77569 = smul32b_32b_x_32b(array_index_77428[literal_77561 > 32'h0000_0009 ? 4'h9 : literal_77561[3:0]], array_index_77564[add_77559 > 32'h0000_0009 ? 4'h9 : add_77559[3:0]]);
  assign add_77571 = array_index_77565[add_77559 > 32'h0000_0009 ? 4'h9 : add_77559[3:0]] + smul_77569;
  assign array_update_77573[0] = add_77559 == 32'h0000_0000 ? add_77571 : array_index_77565[0];
  assign array_update_77573[1] = add_77559 == 32'h0000_0001 ? add_77571 : array_index_77565[1];
  assign array_update_77573[2] = add_77559 == 32'h0000_0002 ? add_77571 : array_index_77565[2];
  assign array_update_77573[3] = add_77559 == 32'h0000_0003 ? add_77571 : array_index_77565[3];
  assign array_update_77573[4] = add_77559 == 32'h0000_0004 ? add_77571 : array_index_77565[4];
  assign array_update_77573[5] = add_77559 == 32'h0000_0005 ? add_77571 : array_index_77565[5];
  assign array_update_77573[6] = add_77559 == 32'h0000_0006 ? add_77571 : array_index_77565[6];
  assign array_update_77573[7] = add_77559 == 32'h0000_0007 ? add_77571 : array_index_77565[7];
  assign array_update_77573[8] = add_77559 == 32'h0000_0008 ? add_77571 : array_index_77565[8];
  assign array_update_77573[9] = add_77559 == 32'h0000_0009 ? add_77571 : array_index_77565[9];
  assign add_77574 = literal_77561 + 32'h0000_0001;
  assign array_update_77575[0] = add_77421 == 32'h0000_0000 ? array_update_77573 : array_update_77562[0];
  assign array_update_77575[1] = add_77421 == 32'h0000_0001 ? array_update_77573 : array_update_77562[1];
  assign array_update_77575[2] = add_77421 == 32'h0000_0002 ? array_update_77573 : array_update_77562[2];
  assign array_update_77575[3] = add_77421 == 32'h0000_0003 ? array_update_77573 : array_update_77562[3];
  assign array_update_77575[4] = add_77421 == 32'h0000_0004 ? array_update_77573 : array_update_77562[4];
  assign array_update_77575[5] = add_77421 == 32'h0000_0005 ? array_update_77573 : array_update_77562[5];
  assign array_update_77575[6] = add_77421 == 32'h0000_0006 ? array_update_77573 : array_update_77562[6];
  assign array_update_77575[7] = add_77421 == 32'h0000_0007 ? array_update_77573 : array_update_77562[7];
  assign array_update_77575[8] = add_77421 == 32'h0000_0008 ? array_update_77573 : array_update_77562[8];
  assign array_update_77575[9] = add_77421 == 32'h0000_0009 ? array_update_77573 : array_update_77562[9];
  assign array_index_77577 = array_update_72021[add_77574 > 32'h0000_0009 ? 4'h9 : add_77574[3:0]];
  assign array_index_77578 = array_update_77575[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_77582 = smul32b_32b_x_32b(array_index_77428[add_77574 > 32'h0000_0009 ? 4'h9 : add_77574[3:0]], array_index_77577[add_77559 > 32'h0000_0009 ? 4'h9 : add_77559[3:0]]);
  assign add_77584 = array_index_77578[add_77559 > 32'h0000_0009 ? 4'h9 : add_77559[3:0]] + smul_77582;
  assign array_update_77586[0] = add_77559 == 32'h0000_0000 ? add_77584 : array_index_77578[0];
  assign array_update_77586[1] = add_77559 == 32'h0000_0001 ? add_77584 : array_index_77578[1];
  assign array_update_77586[2] = add_77559 == 32'h0000_0002 ? add_77584 : array_index_77578[2];
  assign array_update_77586[3] = add_77559 == 32'h0000_0003 ? add_77584 : array_index_77578[3];
  assign array_update_77586[4] = add_77559 == 32'h0000_0004 ? add_77584 : array_index_77578[4];
  assign array_update_77586[5] = add_77559 == 32'h0000_0005 ? add_77584 : array_index_77578[5];
  assign array_update_77586[6] = add_77559 == 32'h0000_0006 ? add_77584 : array_index_77578[6];
  assign array_update_77586[7] = add_77559 == 32'h0000_0007 ? add_77584 : array_index_77578[7];
  assign array_update_77586[8] = add_77559 == 32'h0000_0008 ? add_77584 : array_index_77578[8];
  assign array_update_77586[9] = add_77559 == 32'h0000_0009 ? add_77584 : array_index_77578[9];
  assign add_77587 = add_77574 + 32'h0000_0001;
  assign array_update_77588[0] = add_77421 == 32'h0000_0000 ? array_update_77586 : array_update_77575[0];
  assign array_update_77588[1] = add_77421 == 32'h0000_0001 ? array_update_77586 : array_update_77575[1];
  assign array_update_77588[2] = add_77421 == 32'h0000_0002 ? array_update_77586 : array_update_77575[2];
  assign array_update_77588[3] = add_77421 == 32'h0000_0003 ? array_update_77586 : array_update_77575[3];
  assign array_update_77588[4] = add_77421 == 32'h0000_0004 ? array_update_77586 : array_update_77575[4];
  assign array_update_77588[5] = add_77421 == 32'h0000_0005 ? array_update_77586 : array_update_77575[5];
  assign array_update_77588[6] = add_77421 == 32'h0000_0006 ? array_update_77586 : array_update_77575[6];
  assign array_update_77588[7] = add_77421 == 32'h0000_0007 ? array_update_77586 : array_update_77575[7];
  assign array_update_77588[8] = add_77421 == 32'h0000_0008 ? array_update_77586 : array_update_77575[8];
  assign array_update_77588[9] = add_77421 == 32'h0000_0009 ? array_update_77586 : array_update_77575[9];
  assign array_index_77590 = array_update_72021[add_77587 > 32'h0000_0009 ? 4'h9 : add_77587[3:0]];
  assign array_index_77591 = array_update_77588[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_77595 = smul32b_32b_x_32b(array_index_77428[add_77587 > 32'h0000_0009 ? 4'h9 : add_77587[3:0]], array_index_77590[add_77559 > 32'h0000_0009 ? 4'h9 : add_77559[3:0]]);
  assign add_77597 = array_index_77591[add_77559 > 32'h0000_0009 ? 4'h9 : add_77559[3:0]] + smul_77595;
  assign array_update_77599[0] = add_77559 == 32'h0000_0000 ? add_77597 : array_index_77591[0];
  assign array_update_77599[1] = add_77559 == 32'h0000_0001 ? add_77597 : array_index_77591[1];
  assign array_update_77599[2] = add_77559 == 32'h0000_0002 ? add_77597 : array_index_77591[2];
  assign array_update_77599[3] = add_77559 == 32'h0000_0003 ? add_77597 : array_index_77591[3];
  assign array_update_77599[4] = add_77559 == 32'h0000_0004 ? add_77597 : array_index_77591[4];
  assign array_update_77599[5] = add_77559 == 32'h0000_0005 ? add_77597 : array_index_77591[5];
  assign array_update_77599[6] = add_77559 == 32'h0000_0006 ? add_77597 : array_index_77591[6];
  assign array_update_77599[7] = add_77559 == 32'h0000_0007 ? add_77597 : array_index_77591[7];
  assign array_update_77599[8] = add_77559 == 32'h0000_0008 ? add_77597 : array_index_77591[8];
  assign array_update_77599[9] = add_77559 == 32'h0000_0009 ? add_77597 : array_index_77591[9];
  assign add_77600 = add_77587 + 32'h0000_0001;
  assign array_update_77601[0] = add_77421 == 32'h0000_0000 ? array_update_77599 : array_update_77588[0];
  assign array_update_77601[1] = add_77421 == 32'h0000_0001 ? array_update_77599 : array_update_77588[1];
  assign array_update_77601[2] = add_77421 == 32'h0000_0002 ? array_update_77599 : array_update_77588[2];
  assign array_update_77601[3] = add_77421 == 32'h0000_0003 ? array_update_77599 : array_update_77588[3];
  assign array_update_77601[4] = add_77421 == 32'h0000_0004 ? array_update_77599 : array_update_77588[4];
  assign array_update_77601[5] = add_77421 == 32'h0000_0005 ? array_update_77599 : array_update_77588[5];
  assign array_update_77601[6] = add_77421 == 32'h0000_0006 ? array_update_77599 : array_update_77588[6];
  assign array_update_77601[7] = add_77421 == 32'h0000_0007 ? array_update_77599 : array_update_77588[7];
  assign array_update_77601[8] = add_77421 == 32'h0000_0008 ? array_update_77599 : array_update_77588[8];
  assign array_update_77601[9] = add_77421 == 32'h0000_0009 ? array_update_77599 : array_update_77588[9];
  assign array_index_77603 = array_update_72021[add_77600 > 32'h0000_0009 ? 4'h9 : add_77600[3:0]];
  assign array_index_77604 = array_update_77601[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_77608 = smul32b_32b_x_32b(array_index_77428[add_77600 > 32'h0000_0009 ? 4'h9 : add_77600[3:0]], array_index_77603[add_77559 > 32'h0000_0009 ? 4'h9 : add_77559[3:0]]);
  assign add_77610 = array_index_77604[add_77559 > 32'h0000_0009 ? 4'h9 : add_77559[3:0]] + smul_77608;
  assign array_update_77612[0] = add_77559 == 32'h0000_0000 ? add_77610 : array_index_77604[0];
  assign array_update_77612[1] = add_77559 == 32'h0000_0001 ? add_77610 : array_index_77604[1];
  assign array_update_77612[2] = add_77559 == 32'h0000_0002 ? add_77610 : array_index_77604[2];
  assign array_update_77612[3] = add_77559 == 32'h0000_0003 ? add_77610 : array_index_77604[3];
  assign array_update_77612[4] = add_77559 == 32'h0000_0004 ? add_77610 : array_index_77604[4];
  assign array_update_77612[5] = add_77559 == 32'h0000_0005 ? add_77610 : array_index_77604[5];
  assign array_update_77612[6] = add_77559 == 32'h0000_0006 ? add_77610 : array_index_77604[6];
  assign array_update_77612[7] = add_77559 == 32'h0000_0007 ? add_77610 : array_index_77604[7];
  assign array_update_77612[8] = add_77559 == 32'h0000_0008 ? add_77610 : array_index_77604[8];
  assign array_update_77612[9] = add_77559 == 32'h0000_0009 ? add_77610 : array_index_77604[9];
  assign add_77613 = add_77600 + 32'h0000_0001;
  assign array_update_77614[0] = add_77421 == 32'h0000_0000 ? array_update_77612 : array_update_77601[0];
  assign array_update_77614[1] = add_77421 == 32'h0000_0001 ? array_update_77612 : array_update_77601[1];
  assign array_update_77614[2] = add_77421 == 32'h0000_0002 ? array_update_77612 : array_update_77601[2];
  assign array_update_77614[3] = add_77421 == 32'h0000_0003 ? array_update_77612 : array_update_77601[3];
  assign array_update_77614[4] = add_77421 == 32'h0000_0004 ? array_update_77612 : array_update_77601[4];
  assign array_update_77614[5] = add_77421 == 32'h0000_0005 ? array_update_77612 : array_update_77601[5];
  assign array_update_77614[6] = add_77421 == 32'h0000_0006 ? array_update_77612 : array_update_77601[6];
  assign array_update_77614[7] = add_77421 == 32'h0000_0007 ? array_update_77612 : array_update_77601[7];
  assign array_update_77614[8] = add_77421 == 32'h0000_0008 ? array_update_77612 : array_update_77601[8];
  assign array_update_77614[9] = add_77421 == 32'h0000_0009 ? array_update_77612 : array_update_77601[9];
  assign array_index_77616 = array_update_72021[add_77613 > 32'h0000_0009 ? 4'h9 : add_77613[3:0]];
  assign array_index_77617 = array_update_77614[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_77621 = smul32b_32b_x_32b(array_index_77428[add_77613 > 32'h0000_0009 ? 4'h9 : add_77613[3:0]], array_index_77616[add_77559 > 32'h0000_0009 ? 4'h9 : add_77559[3:0]]);
  assign add_77623 = array_index_77617[add_77559 > 32'h0000_0009 ? 4'h9 : add_77559[3:0]] + smul_77621;
  assign array_update_77625[0] = add_77559 == 32'h0000_0000 ? add_77623 : array_index_77617[0];
  assign array_update_77625[1] = add_77559 == 32'h0000_0001 ? add_77623 : array_index_77617[1];
  assign array_update_77625[2] = add_77559 == 32'h0000_0002 ? add_77623 : array_index_77617[2];
  assign array_update_77625[3] = add_77559 == 32'h0000_0003 ? add_77623 : array_index_77617[3];
  assign array_update_77625[4] = add_77559 == 32'h0000_0004 ? add_77623 : array_index_77617[4];
  assign array_update_77625[5] = add_77559 == 32'h0000_0005 ? add_77623 : array_index_77617[5];
  assign array_update_77625[6] = add_77559 == 32'h0000_0006 ? add_77623 : array_index_77617[6];
  assign array_update_77625[7] = add_77559 == 32'h0000_0007 ? add_77623 : array_index_77617[7];
  assign array_update_77625[8] = add_77559 == 32'h0000_0008 ? add_77623 : array_index_77617[8];
  assign array_update_77625[9] = add_77559 == 32'h0000_0009 ? add_77623 : array_index_77617[9];
  assign add_77626 = add_77613 + 32'h0000_0001;
  assign array_update_77627[0] = add_77421 == 32'h0000_0000 ? array_update_77625 : array_update_77614[0];
  assign array_update_77627[1] = add_77421 == 32'h0000_0001 ? array_update_77625 : array_update_77614[1];
  assign array_update_77627[2] = add_77421 == 32'h0000_0002 ? array_update_77625 : array_update_77614[2];
  assign array_update_77627[3] = add_77421 == 32'h0000_0003 ? array_update_77625 : array_update_77614[3];
  assign array_update_77627[4] = add_77421 == 32'h0000_0004 ? array_update_77625 : array_update_77614[4];
  assign array_update_77627[5] = add_77421 == 32'h0000_0005 ? array_update_77625 : array_update_77614[5];
  assign array_update_77627[6] = add_77421 == 32'h0000_0006 ? array_update_77625 : array_update_77614[6];
  assign array_update_77627[7] = add_77421 == 32'h0000_0007 ? array_update_77625 : array_update_77614[7];
  assign array_update_77627[8] = add_77421 == 32'h0000_0008 ? array_update_77625 : array_update_77614[8];
  assign array_update_77627[9] = add_77421 == 32'h0000_0009 ? array_update_77625 : array_update_77614[9];
  assign array_index_77629 = array_update_72021[add_77626 > 32'h0000_0009 ? 4'h9 : add_77626[3:0]];
  assign array_index_77630 = array_update_77627[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_77634 = smul32b_32b_x_32b(array_index_77428[add_77626 > 32'h0000_0009 ? 4'h9 : add_77626[3:0]], array_index_77629[add_77559 > 32'h0000_0009 ? 4'h9 : add_77559[3:0]]);
  assign add_77636 = array_index_77630[add_77559 > 32'h0000_0009 ? 4'h9 : add_77559[3:0]] + smul_77634;
  assign array_update_77638[0] = add_77559 == 32'h0000_0000 ? add_77636 : array_index_77630[0];
  assign array_update_77638[1] = add_77559 == 32'h0000_0001 ? add_77636 : array_index_77630[1];
  assign array_update_77638[2] = add_77559 == 32'h0000_0002 ? add_77636 : array_index_77630[2];
  assign array_update_77638[3] = add_77559 == 32'h0000_0003 ? add_77636 : array_index_77630[3];
  assign array_update_77638[4] = add_77559 == 32'h0000_0004 ? add_77636 : array_index_77630[4];
  assign array_update_77638[5] = add_77559 == 32'h0000_0005 ? add_77636 : array_index_77630[5];
  assign array_update_77638[6] = add_77559 == 32'h0000_0006 ? add_77636 : array_index_77630[6];
  assign array_update_77638[7] = add_77559 == 32'h0000_0007 ? add_77636 : array_index_77630[7];
  assign array_update_77638[8] = add_77559 == 32'h0000_0008 ? add_77636 : array_index_77630[8];
  assign array_update_77638[9] = add_77559 == 32'h0000_0009 ? add_77636 : array_index_77630[9];
  assign add_77639 = add_77626 + 32'h0000_0001;
  assign array_update_77640[0] = add_77421 == 32'h0000_0000 ? array_update_77638 : array_update_77627[0];
  assign array_update_77640[1] = add_77421 == 32'h0000_0001 ? array_update_77638 : array_update_77627[1];
  assign array_update_77640[2] = add_77421 == 32'h0000_0002 ? array_update_77638 : array_update_77627[2];
  assign array_update_77640[3] = add_77421 == 32'h0000_0003 ? array_update_77638 : array_update_77627[3];
  assign array_update_77640[4] = add_77421 == 32'h0000_0004 ? array_update_77638 : array_update_77627[4];
  assign array_update_77640[5] = add_77421 == 32'h0000_0005 ? array_update_77638 : array_update_77627[5];
  assign array_update_77640[6] = add_77421 == 32'h0000_0006 ? array_update_77638 : array_update_77627[6];
  assign array_update_77640[7] = add_77421 == 32'h0000_0007 ? array_update_77638 : array_update_77627[7];
  assign array_update_77640[8] = add_77421 == 32'h0000_0008 ? array_update_77638 : array_update_77627[8];
  assign array_update_77640[9] = add_77421 == 32'h0000_0009 ? array_update_77638 : array_update_77627[9];
  assign array_index_77642 = array_update_72021[add_77639 > 32'h0000_0009 ? 4'h9 : add_77639[3:0]];
  assign array_index_77643 = array_update_77640[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_77647 = smul32b_32b_x_32b(array_index_77428[add_77639 > 32'h0000_0009 ? 4'h9 : add_77639[3:0]], array_index_77642[add_77559 > 32'h0000_0009 ? 4'h9 : add_77559[3:0]]);
  assign add_77649 = array_index_77643[add_77559 > 32'h0000_0009 ? 4'h9 : add_77559[3:0]] + smul_77647;
  assign array_update_77651[0] = add_77559 == 32'h0000_0000 ? add_77649 : array_index_77643[0];
  assign array_update_77651[1] = add_77559 == 32'h0000_0001 ? add_77649 : array_index_77643[1];
  assign array_update_77651[2] = add_77559 == 32'h0000_0002 ? add_77649 : array_index_77643[2];
  assign array_update_77651[3] = add_77559 == 32'h0000_0003 ? add_77649 : array_index_77643[3];
  assign array_update_77651[4] = add_77559 == 32'h0000_0004 ? add_77649 : array_index_77643[4];
  assign array_update_77651[5] = add_77559 == 32'h0000_0005 ? add_77649 : array_index_77643[5];
  assign array_update_77651[6] = add_77559 == 32'h0000_0006 ? add_77649 : array_index_77643[6];
  assign array_update_77651[7] = add_77559 == 32'h0000_0007 ? add_77649 : array_index_77643[7];
  assign array_update_77651[8] = add_77559 == 32'h0000_0008 ? add_77649 : array_index_77643[8];
  assign array_update_77651[9] = add_77559 == 32'h0000_0009 ? add_77649 : array_index_77643[9];
  assign add_77652 = add_77639 + 32'h0000_0001;
  assign array_update_77653[0] = add_77421 == 32'h0000_0000 ? array_update_77651 : array_update_77640[0];
  assign array_update_77653[1] = add_77421 == 32'h0000_0001 ? array_update_77651 : array_update_77640[1];
  assign array_update_77653[2] = add_77421 == 32'h0000_0002 ? array_update_77651 : array_update_77640[2];
  assign array_update_77653[3] = add_77421 == 32'h0000_0003 ? array_update_77651 : array_update_77640[3];
  assign array_update_77653[4] = add_77421 == 32'h0000_0004 ? array_update_77651 : array_update_77640[4];
  assign array_update_77653[5] = add_77421 == 32'h0000_0005 ? array_update_77651 : array_update_77640[5];
  assign array_update_77653[6] = add_77421 == 32'h0000_0006 ? array_update_77651 : array_update_77640[6];
  assign array_update_77653[7] = add_77421 == 32'h0000_0007 ? array_update_77651 : array_update_77640[7];
  assign array_update_77653[8] = add_77421 == 32'h0000_0008 ? array_update_77651 : array_update_77640[8];
  assign array_update_77653[9] = add_77421 == 32'h0000_0009 ? array_update_77651 : array_update_77640[9];
  assign array_index_77655 = array_update_72021[add_77652 > 32'h0000_0009 ? 4'h9 : add_77652[3:0]];
  assign array_index_77656 = array_update_77653[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_77660 = smul32b_32b_x_32b(array_index_77428[add_77652 > 32'h0000_0009 ? 4'h9 : add_77652[3:0]], array_index_77655[add_77559 > 32'h0000_0009 ? 4'h9 : add_77559[3:0]]);
  assign add_77662 = array_index_77656[add_77559 > 32'h0000_0009 ? 4'h9 : add_77559[3:0]] + smul_77660;
  assign array_update_77664[0] = add_77559 == 32'h0000_0000 ? add_77662 : array_index_77656[0];
  assign array_update_77664[1] = add_77559 == 32'h0000_0001 ? add_77662 : array_index_77656[1];
  assign array_update_77664[2] = add_77559 == 32'h0000_0002 ? add_77662 : array_index_77656[2];
  assign array_update_77664[3] = add_77559 == 32'h0000_0003 ? add_77662 : array_index_77656[3];
  assign array_update_77664[4] = add_77559 == 32'h0000_0004 ? add_77662 : array_index_77656[4];
  assign array_update_77664[5] = add_77559 == 32'h0000_0005 ? add_77662 : array_index_77656[5];
  assign array_update_77664[6] = add_77559 == 32'h0000_0006 ? add_77662 : array_index_77656[6];
  assign array_update_77664[7] = add_77559 == 32'h0000_0007 ? add_77662 : array_index_77656[7];
  assign array_update_77664[8] = add_77559 == 32'h0000_0008 ? add_77662 : array_index_77656[8];
  assign array_update_77664[9] = add_77559 == 32'h0000_0009 ? add_77662 : array_index_77656[9];
  assign add_77665 = add_77652 + 32'h0000_0001;
  assign array_update_77666[0] = add_77421 == 32'h0000_0000 ? array_update_77664 : array_update_77653[0];
  assign array_update_77666[1] = add_77421 == 32'h0000_0001 ? array_update_77664 : array_update_77653[1];
  assign array_update_77666[2] = add_77421 == 32'h0000_0002 ? array_update_77664 : array_update_77653[2];
  assign array_update_77666[3] = add_77421 == 32'h0000_0003 ? array_update_77664 : array_update_77653[3];
  assign array_update_77666[4] = add_77421 == 32'h0000_0004 ? array_update_77664 : array_update_77653[4];
  assign array_update_77666[5] = add_77421 == 32'h0000_0005 ? array_update_77664 : array_update_77653[5];
  assign array_update_77666[6] = add_77421 == 32'h0000_0006 ? array_update_77664 : array_update_77653[6];
  assign array_update_77666[7] = add_77421 == 32'h0000_0007 ? array_update_77664 : array_update_77653[7];
  assign array_update_77666[8] = add_77421 == 32'h0000_0008 ? array_update_77664 : array_update_77653[8];
  assign array_update_77666[9] = add_77421 == 32'h0000_0009 ? array_update_77664 : array_update_77653[9];
  assign array_index_77668 = array_update_72021[add_77665 > 32'h0000_0009 ? 4'h9 : add_77665[3:0]];
  assign array_index_77669 = array_update_77666[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_77673 = smul32b_32b_x_32b(array_index_77428[add_77665 > 32'h0000_0009 ? 4'h9 : add_77665[3:0]], array_index_77668[add_77559 > 32'h0000_0009 ? 4'h9 : add_77559[3:0]]);
  assign add_77675 = array_index_77669[add_77559 > 32'h0000_0009 ? 4'h9 : add_77559[3:0]] + smul_77673;
  assign array_update_77677[0] = add_77559 == 32'h0000_0000 ? add_77675 : array_index_77669[0];
  assign array_update_77677[1] = add_77559 == 32'h0000_0001 ? add_77675 : array_index_77669[1];
  assign array_update_77677[2] = add_77559 == 32'h0000_0002 ? add_77675 : array_index_77669[2];
  assign array_update_77677[3] = add_77559 == 32'h0000_0003 ? add_77675 : array_index_77669[3];
  assign array_update_77677[4] = add_77559 == 32'h0000_0004 ? add_77675 : array_index_77669[4];
  assign array_update_77677[5] = add_77559 == 32'h0000_0005 ? add_77675 : array_index_77669[5];
  assign array_update_77677[6] = add_77559 == 32'h0000_0006 ? add_77675 : array_index_77669[6];
  assign array_update_77677[7] = add_77559 == 32'h0000_0007 ? add_77675 : array_index_77669[7];
  assign array_update_77677[8] = add_77559 == 32'h0000_0008 ? add_77675 : array_index_77669[8];
  assign array_update_77677[9] = add_77559 == 32'h0000_0009 ? add_77675 : array_index_77669[9];
  assign add_77678 = add_77665 + 32'h0000_0001;
  assign array_update_77679[0] = add_77421 == 32'h0000_0000 ? array_update_77677 : array_update_77666[0];
  assign array_update_77679[1] = add_77421 == 32'h0000_0001 ? array_update_77677 : array_update_77666[1];
  assign array_update_77679[2] = add_77421 == 32'h0000_0002 ? array_update_77677 : array_update_77666[2];
  assign array_update_77679[3] = add_77421 == 32'h0000_0003 ? array_update_77677 : array_update_77666[3];
  assign array_update_77679[4] = add_77421 == 32'h0000_0004 ? array_update_77677 : array_update_77666[4];
  assign array_update_77679[5] = add_77421 == 32'h0000_0005 ? array_update_77677 : array_update_77666[5];
  assign array_update_77679[6] = add_77421 == 32'h0000_0006 ? array_update_77677 : array_update_77666[6];
  assign array_update_77679[7] = add_77421 == 32'h0000_0007 ? array_update_77677 : array_update_77666[7];
  assign array_update_77679[8] = add_77421 == 32'h0000_0008 ? array_update_77677 : array_update_77666[8];
  assign array_update_77679[9] = add_77421 == 32'h0000_0009 ? array_update_77677 : array_update_77666[9];
  assign array_index_77681 = array_update_72021[add_77678 > 32'h0000_0009 ? 4'h9 : add_77678[3:0]];
  assign array_index_77682 = array_update_77679[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_77686 = smul32b_32b_x_32b(array_index_77428[add_77678 > 32'h0000_0009 ? 4'h9 : add_77678[3:0]], array_index_77681[add_77559 > 32'h0000_0009 ? 4'h9 : add_77559[3:0]]);
  assign add_77688 = array_index_77682[add_77559 > 32'h0000_0009 ? 4'h9 : add_77559[3:0]] + smul_77686;
  assign array_update_77689[0] = add_77559 == 32'h0000_0000 ? add_77688 : array_index_77682[0];
  assign array_update_77689[1] = add_77559 == 32'h0000_0001 ? add_77688 : array_index_77682[1];
  assign array_update_77689[2] = add_77559 == 32'h0000_0002 ? add_77688 : array_index_77682[2];
  assign array_update_77689[3] = add_77559 == 32'h0000_0003 ? add_77688 : array_index_77682[3];
  assign array_update_77689[4] = add_77559 == 32'h0000_0004 ? add_77688 : array_index_77682[4];
  assign array_update_77689[5] = add_77559 == 32'h0000_0005 ? add_77688 : array_index_77682[5];
  assign array_update_77689[6] = add_77559 == 32'h0000_0006 ? add_77688 : array_index_77682[6];
  assign array_update_77689[7] = add_77559 == 32'h0000_0007 ? add_77688 : array_index_77682[7];
  assign array_update_77689[8] = add_77559 == 32'h0000_0008 ? add_77688 : array_index_77682[8];
  assign array_update_77689[9] = add_77559 == 32'h0000_0009 ? add_77688 : array_index_77682[9];
  assign array_update_77690[0] = add_77421 == 32'h0000_0000 ? array_update_77689 : array_update_77679[0];
  assign array_update_77690[1] = add_77421 == 32'h0000_0001 ? array_update_77689 : array_update_77679[1];
  assign array_update_77690[2] = add_77421 == 32'h0000_0002 ? array_update_77689 : array_update_77679[2];
  assign array_update_77690[3] = add_77421 == 32'h0000_0003 ? array_update_77689 : array_update_77679[3];
  assign array_update_77690[4] = add_77421 == 32'h0000_0004 ? array_update_77689 : array_update_77679[4];
  assign array_update_77690[5] = add_77421 == 32'h0000_0005 ? array_update_77689 : array_update_77679[5];
  assign array_update_77690[6] = add_77421 == 32'h0000_0006 ? array_update_77689 : array_update_77679[6];
  assign array_update_77690[7] = add_77421 == 32'h0000_0007 ? array_update_77689 : array_update_77679[7];
  assign array_update_77690[8] = add_77421 == 32'h0000_0008 ? array_update_77689 : array_update_77679[8];
  assign array_update_77690[9] = add_77421 == 32'h0000_0009 ? array_update_77689 : array_update_77679[9];
  assign array_index_77692 = array_update_77690[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign add_77694 = add_77559 + 32'h0000_0001;
  assign array_update_77695[0] = add_77694 == 32'h0000_0000 ? 32'h0000_0000 : array_index_77692[0];
  assign array_update_77695[1] = add_77694 == 32'h0000_0001 ? 32'h0000_0000 : array_index_77692[1];
  assign array_update_77695[2] = add_77694 == 32'h0000_0002 ? 32'h0000_0000 : array_index_77692[2];
  assign array_update_77695[3] = add_77694 == 32'h0000_0003 ? 32'h0000_0000 : array_index_77692[3];
  assign array_update_77695[4] = add_77694 == 32'h0000_0004 ? 32'h0000_0000 : array_index_77692[4];
  assign array_update_77695[5] = add_77694 == 32'h0000_0005 ? 32'h0000_0000 : array_index_77692[5];
  assign array_update_77695[6] = add_77694 == 32'h0000_0006 ? 32'h0000_0000 : array_index_77692[6];
  assign array_update_77695[7] = add_77694 == 32'h0000_0007 ? 32'h0000_0000 : array_index_77692[7];
  assign array_update_77695[8] = add_77694 == 32'h0000_0008 ? 32'h0000_0000 : array_index_77692[8];
  assign array_update_77695[9] = add_77694 == 32'h0000_0009 ? 32'h0000_0000 : array_index_77692[9];
  assign literal_77696 = 32'h0000_0000;
  assign array_update_77697[0] = add_77421 == 32'h0000_0000 ? array_update_77695 : array_update_77690[0];
  assign array_update_77697[1] = add_77421 == 32'h0000_0001 ? array_update_77695 : array_update_77690[1];
  assign array_update_77697[2] = add_77421 == 32'h0000_0002 ? array_update_77695 : array_update_77690[2];
  assign array_update_77697[3] = add_77421 == 32'h0000_0003 ? array_update_77695 : array_update_77690[3];
  assign array_update_77697[4] = add_77421 == 32'h0000_0004 ? array_update_77695 : array_update_77690[4];
  assign array_update_77697[5] = add_77421 == 32'h0000_0005 ? array_update_77695 : array_update_77690[5];
  assign array_update_77697[6] = add_77421 == 32'h0000_0006 ? array_update_77695 : array_update_77690[6];
  assign array_update_77697[7] = add_77421 == 32'h0000_0007 ? array_update_77695 : array_update_77690[7];
  assign array_update_77697[8] = add_77421 == 32'h0000_0008 ? array_update_77695 : array_update_77690[8];
  assign array_update_77697[9] = add_77421 == 32'h0000_0009 ? array_update_77695 : array_update_77690[9];
  assign array_index_77699 = array_update_72021[literal_77696 > 32'h0000_0009 ? 4'h9 : literal_77696[3:0]];
  assign array_index_77700 = array_update_77697[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_77704 = smul32b_32b_x_32b(array_index_77428[literal_77696 > 32'h0000_0009 ? 4'h9 : literal_77696[3:0]], array_index_77699[add_77694 > 32'h0000_0009 ? 4'h9 : add_77694[3:0]]);
  assign add_77706 = array_index_77700[add_77694 > 32'h0000_0009 ? 4'h9 : add_77694[3:0]] + smul_77704;
  assign array_update_77708[0] = add_77694 == 32'h0000_0000 ? add_77706 : array_index_77700[0];
  assign array_update_77708[1] = add_77694 == 32'h0000_0001 ? add_77706 : array_index_77700[1];
  assign array_update_77708[2] = add_77694 == 32'h0000_0002 ? add_77706 : array_index_77700[2];
  assign array_update_77708[3] = add_77694 == 32'h0000_0003 ? add_77706 : array_index_77700[3];
  assign array_update_77708[4] = add_77694 == 32'h0000_0004 ? add_77706 : array_index_77700[4];
  assign array_update_77708[5] = add_77694 == 32'h0000_0005 ? add_77706 : array_index_77700[5];
  assign array_update_77708[6] = add_77694 == 32'h0000_0006 ? add_77706 : array_index_77700[6];
  assign array_update_77708[7] = add_77694 == 32'h0000_0007 ? add_77706 : array_index_77700[7];
  assign array_update_77708[8] = add_77694 == 32'h0000_0008 ? add_77706 : array_index_77700[8];
  assign array_update_77708[9] = add_77694 == 32'h0000_0009 ? add_77706 : array_index_77700[9];
  assign add_77709 = literal_77696 + 32'h0000_0001;
  assign array_update_77710[0] = add_77421 == 32'h0000_0000 ? array_update_77708 : array_update_77697[0];
  assign array_update_77710[1] = add_77421 == 32'h0000_0001 ? array_update_77708 : array_update_77697[1];
  assign array_update_77710[2] = add_77421 == 32'h0000_0002 ? array_update_77708 : array_update_77697[2];
  assign array_update_77710[3] = add_77421 == 32'h0000_0003 ? array_update_77708 : array_update_77697[3];
  assign array_update_77710[4] = add_77421 == 32'h0000_0004 ? array_update_77708 : array_update_77697[4];
  assign array_update_77710[5] = add_77421 == 32'h0000_0005 ? array_update_77708 : array_update_77697[5];
  assign array_update_77710[6] = add_77421 == 32'h0000_0006 ? array_update_77708 : array_update_77697[6];
  assign array_update_77710[7] = add_77421 == 32'h0000_0007 ? array_update_77708 : array_update_77697[7];
  assign array_update_77710[8] = add_77421 == 32'h0000_0008 ? array_update_77708 : array_update_77697[8];
  assign array_update_77710[9] = add_77421 == 32'h0000_0009 ? array_update_77708 : array_update_77697[9];
  assign array_index_77712 = array_update_72021[add_77709 > 32'h0000_0009 ? 4'h9 : add_77709[3:0]];
  assign array_index_77713 = array_update_77710[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_77717 = smul32b_32b_x_32b(array_index_77428[add_77709 > 32'h0000_0009 ? 4'h9 : add_77709[3:0]], array_index_77712[add_77694 > 32'h0000_0009 ? 4'h9 : add_77694[3:0]]);
  assign add_77719 = array_index_77713[add_77694 > 32'h0000_0009 ? 4'h9 : add_77694[3:0]] + smul_77717;
  assign array_update_77721[0] = add_77694 == 32'h0000_0000 ? add_77719 : array_index_77713[0];
  assign array_update_77721[1] = add_77694 == 32'h0000_0001 ? add_77719 : array_index_77713[1];
  assign array_update_77721[2] = add_77694 == 32'h0000_0002 ? add_77719 : array_index_77713[2];
  assign array_update_77721[3] = add_77694 == 32'h0000_0003 ? add_77719 : array_index_77713[3];
  assign array_update_77721[4] = add_77694 == 32'h0000_0004 ? add_77719 : array_index_77713[4];
  assign array_update_77721[5] = add_77694 == 32'h0000_0005 ? add_77719 : array_index_77713[5];
  assign array_update_77721[6] = add_77694 == 32'h0000_0006 ? add_77719 : array_index_77713[6];
  assign array_update_77721[7] = add_77694 == 32'h0000_0007 ? add_77719 : array_index_77713[7];
  assign array_update_77721[8] = add_77694 == 32'h0000_0008 ? add_77719 : array_index_77713[8];
  assign array_update_77721[9] = add_77694 == 32'h0000_0009 ? add_77719 : array_index_77713[9];
  assign add_77722 = add_77709 + 32'h0000_0001;
  assign array_update_77723[0] = add_77421 == 32'h0000_0000 ? array_update_77721 : array_update_77710[0];
  assign array_update_77723[1] = add_77421 == 32'h0000_0001 ? array_update_77721 : array_update_77710[1];
  assign array_update_77723[2] = add_77421 == 32'h0000_0002 ? array_update_77721 : array_update_77710[2];
  assign array_update_77723[3] = add_77421 == 32'h0000_0003 ? array_update_77721 : array_update_77710[3];
  assign array_update_77723[4] = add_77421 == 32'h0000_0004 ? array_update_77721 : array_update_77710[4];
  assign array_update_77723[5] = add_77421 == 32'h0000_0005 ? array_update_77721 : array_update_77710[5];
  assign array_update_77723[6] = add_77421 == 32'h0000_0006 ? array_update_77721 : array_update_77710[6];
  assign array_update_77723[7] = add_77421 == 32'h0000_0007 ? array_update_77721 : array_update_77710[7];
  assign array_update_77723[8] = add_77421 == 32'h0000_0008 ? array_update_77721 : array_update_77710[8];
  assign array_update_77723[9] = add_77421 == 32'h0000_0009 ? array_update_77721 : array_update_77710[9];
  assign array_index_77725 = array_update_72021[add_77722 > 32'h0000_0009 ? 4'h9 : add_77722[3:0]];
  assign array_index_77726 = array_update_77723[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_77730 = smul32b_32b_x_32b(array_index_77428[add_77722 > 32'h0000_0009 ? 4'h9 : add_77722[3:0]], array_index_77725[add_77694 > 32'h0000_0009 ? 4'h9 : add_77694[3:0]]);
  assign add_77732 = array_index_77726[add_77694 > 32'h0000_0009 ? 4'h9 : add_77694[3:0]] + smul_77730;
  assign array_update_77734[0] = add_77694 == 32'h0000_0000 ? add_77732 : array_index_77726[0];
  assign array_update_77734[1] = add_77694 == 32'h0000_0001 ? add_77732 : array_index_77726[1];
  assign array_update_77734[2] = add_77694 == 32'h0000_0002 ? add_77732 : array_index_77726[2];
  assign array_update_77734[3] = add_77694 == 32'h0000_0003 ? add_77732 : array_index_77726[3];
  assign array_update_77734[4] = add_77694 == 32'h0000_0004 ? add_77732 : array_index_77726[4];
  assign array_update_77734[5] = add_77694 == 32'h0000_0005 ? add_77732 : array_index_77726[5];
  assign array_update_77734[6] = add_77694 == 32'h0000_0006 ? add_77732 : array_index_77726[6];
  assign array_update_77734[7] = add_77694 == 32'h0000_0007 ? add_77732 : array_index_77726[7];
  assign array_update_77734[8] = add_77694 == 32'h0000_0008 ? add_77732 : array_index_77726[8];
  assign array_update_77734[9] = add_77694 == 32'h0000_0009 ? add_77732 : array_index_77726[9];
  assign add_77735 = add_77722 + 32'h0000_0001;
  assign array_update_77736[0] = add_77421 == 32'h0000_0000 ? array_update_77734 : array_update_77723[0];
  assign array_update_77736[1] = add_77421 == 32'h0000_0001 ? array_update_77734 : array_update_77723[1];
  assign array_update_77736[2] = add_77421 == 32'h0000_0002 ? array_update_77734 : array_update_77723[2];
  assign array_update_77736[3] = add_77421 == 32'h0000_0003 ? array_update_77734 : array_update_77723[3];
  assign array_update_77736[4] = add_77421 == 32'h0000_0004 ? array_update_77734 : array_update_77723[4];
  assign array_update_77736[5] = add_77421 == 32'h0000_0005 ? array_update_77734 : array_update_77723[5];
  assign array_update_77736[6] = add_77421 == 32'h0000_0006 ? array_update_77734 : array_update_77723[6];
  assign array_update_77736[7] = add_77421 == 32'h0000_0007 ? array_update_77734 : array_update_77723[7];
  assign array_update_77736[8] = add_77421 == 32'h0000_0008 ? array_update_77734 : array_update_77723[8];
  assign array_update_77736[9] = add_77421 == 32'h0000_0009 ? array_update_77734 : array_update_77723[9];
  assign array_index_77738 = array_update_72021[add_77735 > 32'h0000_0009 ? 4'h9 : add_77735[3:0]];
  assign array_index_77739 = array_update_77736[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_77743 = smul32b_32b_x_32b(array_index_77428[add_77735 > 32'h0000_0009 ? 4'h9 : add_77735[3:0]], array_index_77738[add_77694 > 32'h0000_0009 ? 4'h9 : add_77694[3:0]]);
  assign add_77745 = array_index_77739[add_77694 > 32'h0000_0009 ? 4'h9 : add_77694[3:0]] + smul_77743;
  assign array_update_77747[0] = add_77694 == 32'h0000_0000 ? add_77745 : array_index_77739[0];
  assign array_update_77747[1] = add_77694 == 32'h0000_0001 ? add_77745 : array_index_77739[1];
  assign array_update_77747[2] = add_77694 == 32'h0000_0002 ? add_77745 : array_index_77739[2];
  assign array_update_77747[3] = add_77694 == 32'h0000_0003 ? add_77745 : array_index_77739[3];
  assign array_update_77747[4] = add_77694 == 32'h0000_0004 ? add_77745 : array_index_77739[4];
  assign array_update_77747[5] = add_77694 == 32'h0000_0005 ? add_77745 : array_index_77739[5];
  assign array_update_77747[6] = add_77694 == 32'h0000_0006 ? add_77745 : array_index_77739[6];
  assign array_update_77747[7] = add_77694 == 32'h0000_0007 ? add_77745 : array_index_77739[7];
  assign array_update_77747[8] = add_77694 == 32'h0000_0008 ? add_77745 : array_index_77739[8];
  assign array_update_77747[9] = add_77694 == 32'h0000_0009 ? add_77745 : array_index_77739[9];
  assign add_77748 = add_77735 + 32'h0000_0001;
  assign array_update_77749[0] = add_77421 == 32'h0000_0000 ? array_update_77747 : array_update_77736[0];
  assign array_update_77749[1] = add_77421 == 32'h0000_0001 ? array_update_77747 : array_update_77736[1];
  assign array_update_77749[2] = add_77421 == 32'h0000_0002 ? array_update_77747 : array_update_77736[2];
  assign array_update_77749[3] = add_77421 == 32'h0000_0003 ? array_update_77747 : array_update_77736[3];
  assign array_update_77749[4] = add_77421 == 32'h0000_0004 ? array_update_77747 : array_update_77736[4];
  assign array_update_77749[5] = add_77421 == 32'h0000_0005 ? array_update_77747 : array_update_77736[5];
  assign array_update_77749[6] = add_77421 == 32'h0000_0006 ? array_update_77747 : array_update_77736[6];
  assign array_update_77749[7] = add_77421 == 32'h0000_0007 ? array_update_77747 : array_update_77736[7];
  assign array_update_77749[8] = add_77421 == 32'h0000_0008 ? array_update_77747 : array_update_77736[8];
  assign array_update_77749[9] = add_77421 == 32'h0000_0009 ? array_update_77747 : array_update_77736[9];
  assign array_index_77751 = array_update_72021[add_77748 > 32'h0000_0009 ? 4'h9 : add_77748[3:0]];
  assign array_index_77752 = array_update_77749[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_77756 = smul32b_32b_x_32b(array_index_77428[add_77748 > 32'h0000_0009 ? 4'h9 : add_77748[3:0]], array_index_77751[add_77694 > 32'h0000_0009 ? 4'h9 : add_77694[3:0]]);
  assign add_77758 = array_index_77752[add_77694 > 32'h0000_0009 ? 4'h9 : add_77694[3:0]] + smul_77756;
  assign array_update_77760[0] = add_77694 == 32'h0000_0000 ? add_77758 : array_index_77752[0];
  assign array_update_77760[1] = add_77694 == 32'h0000_0001 ? add_77758 : array_index_77752[1];
  assign array_update_77760[2] = add_77694 == 32'h0000_0002 ? add_77758 : array_index_77752[2];
  assign array_update_77760[3] = add_77694 == 32'h0000_0003 ? add_77758 : array_index_77752[3];
  assign array_update_77760[4] = add_77694 == 32'h0000_0004 ? add_77758 : array_index_77752[4];
  assign array_update_77760[5] = add_77694 == 32'h0000_0005 ? add_77758 : array_index_77752[5];
  assign array_update_77760[6] = add_77694 == 32'h0000_0006 ? add_77758 : array_index_77752[6];
  assign array_update_77760[7] = add_77694 == 32'h0000_0007 ? add_77758 : array_index_77752[7];
  assign array_update_77760[8] = add_77694 == 32'h0000_0008 ? add_77758 : array_index_77752[8];
  assign array_update_77760[9] = add_77694 == 32'h0000_0009 ? add_77758 : array_index_77752[9];
  assign add_77761 = add_77748 + 32'h0000_0001;
  assign array_update_77762[0] = add_77421 == 32'h0000_0000 ? array_update_77760 : array_update_77749[0];
  assign array_update_77762[1] = add_77421 == 32'h0000_0001 ? array_update_77760 : array_update_77749[1];
  assign array_update_77762[2] = add_77421 == 32'h0000_0002 ? array_update_77760 : array_update_77749[2];
  assign array_update_77762[3] = add_77421 == 32'h0000_0003 ? array_update_77760 : array_update_77749[3];
  assign array_update_77762[4] = add_77421 == 32'h0000_0004 ? array_update_77760 : array_update_77749[4];
  assign array_update_77762[5] = add_77421 == 32'h0000_0005 ? array_update_77760 : array_update_77749[5];
  assign array_update_77762[6] = add_77421 == 32'h0000_0006 ? array_update_77760 : array_update_77749[6];
  assign array_update_77762[7] = add_77421 == 32'h0000_0007 ? array_update_77760 : array_update_77749[7];
  assign array_update_77762[8] = add_77421 == 32'h0000_0008 ? array_update_77760 : array_update_77749[8];
  assign array_update_77762[9] = add_77421 == 32'h0000_0009 ? array_update_77760 : array_update_77749[9];
  assign array_index_77764 = array_update_72021[add_77761 > 32'h0000_0009 ? 4'h9 : add_77761[3:0]];
  assign array_index_77765 = array_update_77762[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_77769 = smul32b_32b_x_32b(array_index_77428[add_77761 > 32'h0000_0009 ? 4'h9 : add_77761[3:0]], array_index_77764[add_77694 > 32'h0000_0009 ? 4'h9 : add_77694[3:0]]);
  assign add_77771 = array_index_77765[add_77694 > 32'h0000_0009 ? 4'h9 : add_77694[3:0]] + smul_77769;
  assign array_update_77773[0] = add_77694 == 32'h0000_0000 ? add_77771 : array_index_77765[0];
  assign array_update_77773[1] = add_77694 == 32'h0000_0001 ? add_77771 : array_index_77765[1];
  assign array_update_77773[2] = add_77694 == 32'h0000_0002 ? add_77771 : array_index_77765[2];
  assign array_update_77773[3] = add_77694 == 32'h0000_0003 ? add_77771 : array_index_77765[3];
  assign array_update_77773[4] = add_77694 == 32'h0000_0004 ? add_77771 : array_index_77765[4];
  assign array_update_77773[5] = add_77694 == 32'h0000_0005 ? add_77771 : array_index_77765[5];
  assign array_update_77773[6] = add_77694 == 32'h0000_0006 ? add_77771 : array_index_77765[6];
  assign array_update_77773[7] = add_77694 == 32'h0000_0007 ? add_77771 : array_index_77765[7];
  assign array_update_77773[8] = add_77694 == 32'h0000_0008 ? add_77771 : array_index_77765[8];
  assign array_update_77773[9] = add_77694 == 32'h0000_0009 ? add_77771 : array_index_77765[9];
  assign add_77774 = add_77761 + 32'h0000_0001;
  assign array_update_77775[0] = add_77421 == 32'h0000_0000 ? array_update_77773 : array_update_77762[0];
  assign array_update_77775[1] = add_77421 == 32'h0000_0001 ? array_update_77773 : array_update_77762[1];
  assign array_update_77775[2] = add_77421 == 32'h0000_0002 ? array_update_77773 : array_update_77762[2];
  assign array_update_77775[3] = add_77421 == 32'h0000_0003 ? array_update_77773 : array_update_77762[3];
  assign array_update_77775[4] = add_77421 == 32'h0000_0004 ? array_update_77773 : array_update_77762[4];
  assign array_update_77775[5] = add_77421 == 32'h0000_0005 ? array_update_77773 : array_update_77762[5];
  assign array_update_77775[6] = add_77421 == 32'h0000_0006 ? array_update_77773 : array_update_77762[6];
  assign array_update_77775[7] = add_77421 == 32'h0000_0007 ? array_update_77773 : array_update_77762[7];
  assign array_update_77775[8] = add_77421 == 32'h0000_0008 ? array_update_77773 : array_update_77762[8];
  assign array_update_77775[9] = add_77421 == 32'h0000_0009 ? array_update_77773 : array_update_77762[9];
  assign array_index_77777 = array_update_72021[add_77774 > 32'h0000_0009 ? 4'h9 : add_77774[3:0]];
  assign array_index_77778 = array_update_77775[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_77782 = smul32b_32b_x_32b(array_index_77428[add_77774 > 32'h0000_0009 ? 4'h9 : add_77774[3:0]], array_index_77777[add_77694 > 32'h0000_0009 ? 4'h9 : add_77694[3:0]]);
  assign add_77784 = array_index_77778[add_77694 > 32'h0000_0009 ? 4'h9 : add_77694[3:0]] + smul_77782;
  assign array_update_77786[0] = add_77694 == 32'h0000_0000 ? add_77784 : array_index_77778[0];
  assign array_update_77786[1] = add_77694 == 32'h0000_0001 ? add_77784 : array_index_77778[1];
  assign array_update_77786[2] = add_77694 == 32'h0000_0002 ? add_77784 : array_index_77778[2];
  assign array_update_77786[3] = add_77694 == 32'h0000_0003 ? add_77784 : array_index_77778[3];
  assign array_update_77786[4] = add_77694 == 32'h0000_0004 ? add_77784 : array_index_77778[4];
  assign array_update_77786[5] = add_77694 == 32'h0000_0005 ? add_77784 : array_index_77778[5];
  assign array_update_77786[6] = add_77694 == 32'h0000_0006 ? add_77784 : array_index_77778[6];
  assign array_update_77786[7] = add_77694 == 32'h0000_0007 ? add_77784 : array_index_77778[7];
  assign array_update_77786[8] = add_77694 == 32'h0000_0008 ? add_77784 : array_index_77778[8];
  assign array_update_77786[9] = add_77694 == 32'h0000_0009 ? add_77784 : array_index_77778[9];
  assign add_77787 = add_77774 + 32'h0000_0001;
  assign array_update_77788[0] = add_77421 == 32'h0000_0000 ? array_update_77786 : array_update_77775[0];
  assign array_update_77788[1] = add_77421 == 32'h0000_0001 ? array_update_77786 : array_update_77775[1];
  assign array_update_77788[2] = add_77421 == 32'h0000_0002 ? array_update_77786 : array_update_77775[2];
  assign array_update_77788[3] = add_77421 == 32'h0000_0003 ? array_update_77786 : array_update_77775[3];
  assign array_update_77788[4] = add_77421 == 32'h0000_0004 ? array_update_77786 : array_update_77775[4];
  assign array_update_77788[5] = add_77421 == 32'h0000_0005 ? array_update_77786 : array_update_77775[5];
  assign array_update_77788[6] = add_77421 == 32'h0000_0006 ? array_update_77786 : array_update_77775[6];
  assign array_update_77788[7] = add_77421 == 32'h0000_0007 ? array_update_77786 : array_update_77775[7];
  assign array_update_77788[8] = add_77421 == 32'h0000_0008 ? array_update_77786 : array_update_77775[8];
  assign array_update_77788[9] = add_77421 == 32'h0000_0009 ? array_update_77786 : array_update_77775[9];
  assign array_index_77790 = array_update_72021[add_77787 > 32'h0000_0009 ? 4'h9 : add_77787[3:0]];
  assign array_index_77791 = array_update_77788[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_77795 = smul32b_32b_x_32b(array_index_77428[add_77787 > 32'h0000_0009 ? 4'h9 : add_77787[3:0]], array_index_77790[add_77694 > 32'h0000_0009 ? 4'h9 : add_77694[3:0]]);
  assign add_77797 = array_index_77791[add_77694 > 32'h0000_0009 ? 4'h9 : add_77694[3:0]] + smul_77795;
  assign array_update_77799[0] = add_77694 == 32'h0000_0000 ? add_77797 : array_index_77791[0];
  assign array_update_77799[1] = add_77694 == 32'h0000_0001 ? add_77797 : array_index_77791[1];
  assign array_update_77799[2] = add_77694 == 32'h0000_0002 ? add_77797 : array_index_77791[2];
  assign array_update_77799[3] = add_77694 == 32'h0000_0003 ? add_77797 : array_index_77791[3];
  assign array_update_77799[4] = add_77694 == 32'h0000_0004 ? add_77797 : array_index_77791[4];
  assign array_update_77799[5] = add_77694 == 32'h0000_0005 ? add_77797 : array_index_77791[5];
  assign array_update_77799[6] = add_77694 == 32'h0000_0006 ? add_77797 : array_index_77791[6];
  assign array_update_77799[7] = add_77694 == 32'h0000_0007 ? add_77797 : array_index_77791[7];
  assign array_update_77799[8] = add_77694 == 32'h0000_0008 ? add_77797 : array_index_77791[8];
  assign array_update_77799[9] = add_77694 == 32'h0000_0009 ? add_77797 : array_index_77791[9];
  assign add_77800 = add_77787 + 32'h0000_0001;
  assign array_update_77801[0] = add_77421 == 32'h0000_0000 ? array_update_77799 : array_update_77788[0];
  assign array_update_77801[1] = add_77421 == 32'h0000_0001 ? array_update_77799 : array_update_77788[1];
  assign array_update_77801[2] = add_77421 == 32'h0000_0002 ? array_update_77799 : array_update_77788[2];
  assign array_update_77801[3] = add_77421 == 32'h0000_0003 ? array_update_77799 : array_update_77788[3];
  assign array_update_77801[4] = add_77421 == 32'h0000_0004 ? array_update_77799 : array_update_77788[4];
  assign array_update_77801[5] = add_77421 == 32'h0000_0005 ? array_update_77799 : array_update_77788[5];
  assign array_update_77801[6] = add_77421 == 32'h0000_0006 ? array_update_77799 : array_update_77788[6];
  assign array_update_77801[7] = add_77421 == 32'h0000_0007 ? array_update_77799 : array_update_77788[7];
  assign array_update_77801[8] = add_77421 == 32'h0000_0008 ? array_update_77799 : array_update_77788[8];
  assign array_update_77801[9] = add_77421 == 32'h0000_0009 ? array_update_77799 : array_update_77788[9];
  assign array_index_77803 = array_update_72021[add_77800 > 32'h0000_0009 ? 4'h9 : add_77800[3:0]];
  assign array_index_77804 = array_update_77801[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_77808 = smul32b_32b_x_32b(array_index_77428[add_77800 > 32'h0000_0009 ? 4'h9 : add_77800[3:0]], array_index_77803[add_77694 > 32'h0000_0009 ? 4'h9 : add_77694[3:0]]);
  assign add_77810 = array_index_77804[add_77694 > 32'h0000_0009 ? 4'h9 : add_77694[3:0]] + smul_77808;
  assign array_update_77812[0] = add_77694 == 32'h0000_0000 ? add_77810 : array_index_77804[0];
  assign array_update_77812[1] = add_77694 == 32'h0000_0001 ? add_77810 : array_index_77804[1];
  assign array_update_77812[2] = add_77694 == 32'h0000_0002 ? add_77810 : array_index_77804[2];
  assign array_update_77812[3] = add_77694 == 32'h0000_0003 ? add_77810 : array_index_77804[3];
  assign array_update_77812[4] = add_77694 == 32'h0000_0004 ? add_77810 : array_index_77804[4];
  assign array_update_77812[5] = add_77694 == 32'h0000_0005 ? add_77810 : array_index_77804[5];
  assign array_update_77812[6] = add_77694 == 32'h0000_0006 ? add_77810 : array_index_77804[6];
  assign array_update_77812[7] = add_77694 == 32'h0000_0007 ? add_77810 : array_index_77804[7];
  assign array_update_77812[8] = add_77694 == 32'h0000_0008 ? add_77810 : array_index_77804[8];
  assign array_update_77812[9] = add_77694 == 32'h0000_0009 ? add_77810 : array_index_77804[9];
  assign add_77813 = add_77800 + 32'h0000_0001;
  assign array_update_77814[0] = add_77421 == 32'h0000_0000 ? array_update_77812 : array_update_77801[0];
  assign array_update_77814[1] = add_77421 == 32'h0000_0001 ? array_update_77812 : array_update_77801[1];
  assign array_update_77814[2] = add_77421 == 32'h0000_0002 ? array_update_77812 : array_update_77801[2];
  assign array_update_77814[3] = add_77421 == 32'h0000_0003 ? array_update_77812 : array_update_77801[3];
  assign array_update_77814[4] = add_77421 == 32'h0000_0004 ? array_update_77812 : array_update_77801[4];
  assign array_update_77814[5] = add_77421 == 32'h0000_0005 ? array_update_77812 : array_update_77801[5];
  assign array_update_77814[6] = add_77421 == 32'h0000_0006 ? array_update_77812 : array_update_77801[6];
  assign array_update_77814[7] = add_77421 == 32'h0000_0007 ? array_update_77812 : array_update_77801[7];
  assign array_update_77814[8] = add_77421 == 32'h0000_0008 ? array_update_77812 : array_update_77801[8];
  assign array_update_77814[9] = add_77421 == 32'h0000_0009 ? array_update_77812 : array_update_77801[9];
  assign array_index_77816 = array_update_72021[add_77813 > 32'h0000_0009 ? 4'h9 : add_77813[3:0]];
  assign array_index_77817 = array_update_77814[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_77821 = smul32b_32b_x_32b(array_index_77428[add_77813 > 32'h0000_0009 ? 4'h9 : add_77813[3:0]], array_index_77816[add_77694 > 32'h0000_0009 ? 4'h9 : add_77694[3:0]]);
  assign add_77823 = array_index_77817[add_77694 > 32'h0000_0009 ? 4'h9 : add_77694[3:0]] + smul_77821;
  assign array_update_77824[0] = add_77694 == 32'h0000_0000 ? add_77823 : array_index_77817[0];
  assign array_update_77824[1] = add_77694 == 32'h0000_0001 ? add_77823 : array_index_77817[1];
  assign array_update_77824[2] = add_77694 == 32'h0000_0002 ? add_77823 : array_index_77817[2];
  assign array_update_77824[3] = add_77694 == 32'h0000_0003 ? add_77823 : array_index_77817[3];
  assign array_update_77824[4] = add_77694 == 32'h0000_0004 ? add_77823 : array_index_77817[4];
  assign array_update_77824[5] = add_77694 == 32'h0000_0005 ? add_77823 : array_index_77817[5];
  assign array_update_77824[6] = add_77694 == 32'h0000_0006 ? add_77823 : array_index_77817[6];
  assign array_update_77824[7] = add_77694 == 32'h0000_0007 ? add_77823 : array_index_77817[7];
  assign array_update_77824[8] = add_77694 == 32'h0000_0008 ? add_77823 : array_index_77817[8];
  assign array_update_77824[9] = add_77694 == 32'h0000_0009 ? add_77823 : array_index_77817[9];
  assign array_update_77825[0] = add_77421 == 32'h0000_0000 ? array_update_77824 : array_update_77814[0];
  assign array_update_77825[1] = add_77421 == 32'h0000_0001 ? array_update_77824 : array_update_77814[1];
  assign array_update_77825[2] = add_77421 == 32'h0000_0002 ? array_update_77824 : array_update_77814[2];
  assign array_update_77825[3] = add_77421 == 32'h0000_0003 ? array_update_77824 : array_update_77814[3];
  assign array_update_77825[4] = add_77421 == 32'h0000_0004 ? array_update_77824 : array_update_77814[4];
  assign array_update_77825[5] = add_77421 == 32'h0000_0005 ? array_update_77824 : array_update_77814[5];
  assign array_update_77825[6] = add_77421 == 32'h0000_0006 ? array_update_77824 : array_update_77814[6];
  assign array_update_77825[7] = add_77421 == 32'h0000_0007 ? array_update_77824 : array_update_77814[7];
  assign array_update_77825[8] = add_77421 == 32'h0000_0008 ? array_update_77824 : array_update_77814[8];
  assign array_update_77825[9] = add_77421 == 32'h0000_0009 ? array_update_77824 : array_update_77814[9];
  assign array_index_77827 = array_update_77825[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign add_77829 = add_77694 + 32'h0000_0001;
  assign array_update_77830[0] = add_77829 == 32'h0000_0000 ? 32'h0000_0000 : array_index_77827[0];
  assign array_update_77830[1] = add_77829 == 32'h0000_0001 ? 32'h0000_0000 : array_index_77827[1];
  assign array_update_77830[2] = add_77829 == 32'h0000_0002 ? 32'h0000_0000 : array_index_77827[2];
  assign array_update_77830[3] = add_77829 == 32'h0000_0003 ? 32'h0000_0000 : array_index_77827[3];
  assign array_update_77830[4] = add_77829 == 32'h0000_0004 ? 32'h0000_0000 : array_index_77827[4];
  assign array_update_77830[5] = add_77829 == 32'h0000_0005 ? 32'h0000_0000 : array_index_77827[5];
  assign array_update_77830[6] = add_77829 == 32'h0000_0006 ? 32'h0000_0000 : array_index_77827[6];
  assign array_update_77830[7] = add_77829 == 32'h0000_0007 ? 32'h0000_0000 : array_index_77827[7];
  assign array_update_77830[8] = add_77829 == 32'h0000_0008 ? 32'h0000_0000 : array_index_77827[8];
  assign array_update_77830[9] = add_77829 == 32'h0000_0009 ? 32'h0000_0000 : array_index_77827[9];
  assign literal_77831 = 32'h0000_0000;
  assign array_update_77832[0] = add_77421 == 32'h0000_0000 ? array_update_77830 : array_update_77825[0];
  assign array_update_77832[1] = add_77421 == 32'h0000_0001 ? array_update_77830 : array_update_77825[1];
  assign array_update_77832[2] = add_77421 == 32'h0000_0002 ? array_update_77830 : array_update_77825[2];
  assign array_update_77832[3] = add_77421 == 32'h0000_0003 ? array_update_77830 : array_update_77825[3];
  assign array_update_77832[4] = add_77421 == 32'h0000_0004 ? array_update_77830 : array_update_77825[4];
  assign array_update_77832[5] = add_77421 == 32'h0000_0005 ? array_update_77830 : array_update_77825[5];
  assign array_update_77832[6] = add_77421 == 32'h0000_0006 ? array_update_77830 : array_update_77825[6];
  assign array_update_77832[7] = add_77421 == 32'h0000_0007 ? array_update_77830 : array_update_77825[7];
  assign array_update_77832[8] = add_77421 == 32'h0000_0008 ? array_update_77830 : array_update_77825[8];
  assign array_update_77832[9] = add_77421 == 32'h0000_0009 ? array_update_77830 : array_update_77825[9];
  assign array_index_77834 = array_update_72021[literal_77831 > 32'h0000_0009 ? 4'h9 : literal_77831[3:0]];
  assign array_index_77835 = array_update_77832[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_77839 = smul32b_32b_x_32b(array_index_77428[literal_77831 > 32'h0000_0009 ? 4'h9 : literal_77831[3:0]], array_index_77834[add_77829 > 32'h0000_0009 ? 4'h9 : add_77829[3:0]]);
  assign add_77841 = array_index_77835[add_77829 > 32'h0000_0009 ? 4'h9 : add_77829[3:0]] + smul_77839;
  assign array_update_77843[0] = add_77829 == 32'h0000_0000 ? add_77841 : array_index_77835[0];
  assign array_update_77843[1] = add_77829 == 32'h0000_0001 ? add_77841 : array_index_77835[1];
  assign array_update_77843[2] = add_77829 == 32'h0000_0002 ? add_77841 : array_index_77835[2];
  assign array_update_77843[3] = add_77829 == 32'h0000_0003 ? add_77841 : array_index_77835[3];
  assign array_update_77843[4] = add_77829 == 32'h0000_0004 ? add_77841 : array_index_77835[4];
  assign array_update_77843[5] = add_77829 == 32'h0000_0005 ? add_77841 : array_index_77835[5];
  assign array_update_77843[6] = add_77829 == 32'h0000_0006 ? add_77841 : array_index_77835[6];
  assign array_update_77843[7] = add_77829 == 32'h0000_0007 ? add_77841 : array_index_77835[7];
  assign array_update_77843[8] = add_77829 == 32'h0000_0008 ? add_77841 : array_index_77835[8];
  assign array_update_77843[9] = add_77829 == 32'h0000_0009 ? add_77841 : array_index_77835[9];
  assign add_77844 = literal_77831 + 32'h0000_0001;
  assign array_update_77845[0] = add_77421 == 32'h0000_0000 ? array_update_77843 : array_update_77832[0];
  assign array_update_77845[1] = add_77421 == 32'h0000_0001 ? array_update_77843 : array_update_77832[1];
  assign array_update_77845[2] = add_77421 == 32'h0000_0002 ? array_update_77843 : array_update_77832[2];
  assign array_update_77845[3] = add_77421 == 32'h0000_0003 ? array_update_77843 : array_update_77832[3];
  assign array_update_77845[4] = add_77421 == 32'h0000_0004 ? array_update_77843 : array_update_77832[4];
  assign array_update_77845[5] = add_77421 == 32'h0000_0005 ? array_update_77843 : array_update_77832[5];
  assign array_update_77845[6] = add_77421 == 32'h0000_0006 ? array_update_77843 : array_update_77832[6];
  assign array_update_77845[7] = add_77421 == 32'h0000_0007 ? array_update_77843 : array_update_77832[7];
  assign array_update_77845[8] = add_77421 == 32'h0000_0008 ? array_update_77843 : array_update_77832[8];
  assign array_update_77845[9] = add_77421 == 32'h0000_0009 ? array_update_77843 : array_update_77832[9];
  assign array_index_77847 = array_update_72021[add_77844 > 32'h0000_0009 ? 4'h9 : add_77844[3:0]];
  assign array_index_77848 = array_update_77845[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_77852 = smul32b_32b_x_32b(array_index_77428[add_77844 > 32'h0000_0009 ? 4'h9 : add_77844[3:0]], array_index_77847[add_77829 > 32'h0000_0009 ? 4'h9 : add_77829[3:0]]);
  assign add_77854 = array_index_77848[add_77829 > 32'h0000_0009 ? 4'h9 : add_77829[3:0]] + smul_77852;
  assign array_update_77856[0] = add_77829 == 32'h0000_0000 ? add_77854 : array_index_77848[0];
  assign array_update_77856[1] = add_77829 == 32'h0000_0001 ? add_77854 : array_index_77848[1];
  assign array_update_77856[2] = add_77829 == 32'h0000_0002 ? add_77854 : array_index_77848[2];
  assign array_update_77856[3] = add_77829 == 32'h0000_0003 ? add_77854 : array_index_77848[3];
  assign array_update_77856[4] = add_77829 == 32'h0000_0004 ? add_77854 : array_index_77848[4];
  assign array_update_77856[5] = add_77829 == 32'h0000_0005 ? add_77854 : array_index_77848[5];
  assign array_update_77856[6] = add_77829 == 32'h0000_0006 ? add_77854 : array_index_77848[6];
  assign array_update_77856[7] = add_77829 == 32'h0000_0007 ? add_77854 : array_index_77848[7];
  assign array_update_77856[8] = add_77829 == 32'h0000_0008 ? add_77854 : array_index_77848[8];
  assign array_update_77856[9] = add_77829 == 32'h0000_0009 ? add_77854 : array_index_77848[9];
  assign add_77857 = add_77844 + 32'h0000_0001;
  assign array_update_77858[0] = add_77421 == 32'h0000_0000 ? array_update_77856 : array_update_77845[0];
  assign array_update_77858[1] = add_77421 == 32'h0000_0001 ? array_update_77856 : array_update_77845[1];
  assign array_update_77858[2] = add_77421 == 32'h0000_0002 ? array_update_77856 : array_update_77845[2];
  assign array_update_77858[3] = add_77421 == 32'h0000_0003 ? array_update_77856 : array_update_77845[3];
  assign array_update_77858[4] = add_77421 == 32'h0000_0004 ? array_update_77856 : array_update_77845[4];
  assign array_update_77858[5] = add_77421 == 32'h0000_0005 ? array_update_77856 : array_update_77845[5];
  assign array_update_77858[6] = add_77421 == 32'h0000_0006 ? array_update_77856 : array_update_77845[6];
  assign array_update_77858[7] = add_77421 == 32'h0000_0007 ? array_update_77856 : array_update_77845[7];
  assign array_update_77858[8] = add_77421 == 32'h0000_0008 ? array_update_77856 : array_update_77845[8];
  assign array_update_77858[9] = add_77421 == 32'h0000_0009 ? array_update_77856 : array_update_77845[9];
  assign array_index_77860 = array_update_72021[add_77857 > 32'h0000_0009 ? 4'h9 : add_77857[3:0]];
  assign array_index_77861 = array_update_77858[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_77865 = smul32b_32b_x_32b(array_index_77428[add_77857 > 32'h0000_0009 ? 4'h9 : add_77857[3:0]], array_index_77860[add_77829 > 32'h0000_0009 ? 4'h9 : add_77829[3:0]]);
  assign add_77867 = array_index_77861[add_77829 > 32'h0000_0009 ? 4'h9 : add_77829[3:0]] + smul_77865;
  assign array_update_77869[0] = add_77829 == 32'h0000_0000 ? add_77867 : array_index_77861[0];
  assign array_update_77869[1] = add_77829 == 32'h0000_0001 ? add_77867 : array_index_77861[1];
  assign array_update_77869[2] = add_77829 == 32'h0000_0002 ? add_77867 : array_index_77861[2];
  assign array_update_77869[3] = add_77829 == 32'h0000_0003 ? add_77867 : array_index_77861[3];
  assign array_update_77869[4] = add_77829 == 32'h0000_0004 ? add_77867 : array_index_77861[4];
  assign array_update_77869[5] = add_77829 == 32'h0000_0005 ? add_77867 : array_index_77861[5];
  assign array_update_77869[6] = add_77829 == 32'h0000_0006 ? add_77867 : array_index_77861[6];
  assign array_update_77869[7] = add_77829 == 32'h0000_0007 ? add_77867 : array_index_77861[7];
  assign array_update_77869[8] = add_77829 == 32'h0000_0008 ? add_77867 : array_index_77861[8];
  assign array_update_77869[9] = add_77829 == 32'h0000_0009 ? add_77867 : array_index_77861[9];
  assign add_77870 = add_77857 + 32'h0000_0001;
  assign array_update_77871[0] = add_77421 == 32'h0000_0000 ? array_update_77869 : array_update_77858[0];
  assign array_update_77871[1] = add_77421 == 32'h0000_0001 ? array_update_77869 : array_update_77858[1];
  assign array_update_77871[2] = add_77421 == 32'h0000_0002 ? array_update_77869 : array_update_77858[2];
  assign array_update_77871[3] = add_77421 == 32'h0000_0003 ? array_update_77869 : array_update_77858[3];
  assign array_update_77871[4] = add_77421 == 32'h0000_0004 ? array_update_77869 : array_update_77858[4];
  assign array_update_77871[5] = add_77421 == 32'h0000_0005 ? array_update_77869 : array_update_77858[5];
  assign array_update_77871[6] = add_77421 == 32'h0000_0006 ? array_update_77869 : array_update_77858[6];
  assign array_update_77871[7] = add_77421 == 32'h0000_0007 ? array_update_77869 : array_update_77858[7];
  assign array_update_77871[8] = add_77421 == 32'h0000_0008 ? array_update_77869 : array_update_77858[8];
  assign array_update_77871[9] = add_77421 == 32'h0000_0009 ? array_update_77869 : array_update_77858[9];
  assign array_index_77873 = array_update_72021[add_77870 > 32'h0000_0009 ? 4'h9 : add_77870[3:0]];
  assign array_index_77874 = array_update_77871[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_77878 = smul32b_32b_x_32b(array_index_77428[add_77870 > 32'h0000_0009 ? 4'h9 : add_77870[3:0]], array_index_77873[add_77829 > 32'h0000_0009 ? 4'h9 : add_77829[3:0]]);
  assign add_77880 = array_index_77874[add_77829 > 32'h0000_0009 ? 4'h9 : add_77829[3:0]] + smul_77878;
  assign array_update_77882[0] = add_77829 == 32'h0000_0000 ? add_77880 : array_index_77874[0];
  assign array_update_77882[1] = add_77829 == 32'h0000_0001 ? add_77880 : array_index_77874[1];
  assign array_update_77882[2] = add_77829 == 32'h0000_0002 ? add_77880 : array_index_77874[2];
  assign array_update_77882[3] = add_77829 == 32'h0000_0003 ? add_77880 : array_index_77874[3];
  assign array_update_77882[4] = add_77829 == 32'h0000_0004 ? add_77880 : array_index_77874[4];
  assign array_update_77882[5] = add_77829 == 32'h0000_0005 ? add_77880 : array_index_77874[5];
  assign array_update_77882[6] = add_77829 == 32'h0000_0006 ? add_77880 : array_index_77874[6];
  assign array_update_77882[7] = add_77829 == 32'h0000_0007 ? add_77880 : array_index_77874[7];
  assign array_update_77882[8] = add_77829 == 32'h0000_0008 ? add_77880 : array_index_77874[8];
  assign array_update_77882[9] = add_77829 == 32'h0000_0009 ? add_77880 : array_index_77874[9];
  assign add_77883 = add_77870 + 32'h0000_0001;
  assign array_update_77884[0] = add_77421 == 32'h0000_0000 ? array_update_77882 : array_update_77871[0];
  assign array_update_77884[1] = add_77421 == 32'h0000_0001 ? array_update_77882 : array_update_77871[1];
  assign array_update_77884[2] = add_77421 == 32'h0000_0002 ? array_update_77882 : array_update_77871[2];
  assign array_update_77884[3] = add_77421 == 32'h0000_0003 ? array_update_77882 : array_update_77871[3];
  assign array_update_77884[4] = add_77421 == 32'h0000_0004 ? array_update_77882 : array_update_77871[4];
  assign array_update_77884[5] = add_77421 == 32'h0000_0005 ? array_update_77882 : array_update_77871[5];
  assign array_update_77884[6] = add_77421 == 32'h0000_0006 ? array_update_77882 : array_update_77871[6];
  assign array_update_77884[7] = add_77421 == 32'h0000_0007 ? array_update_77882 : array_update_77871[7];
  assign array_update_77884[8] = add_77421 == 32'h0000_0008 ? array_update_77882 : array_update_77871[8];
  assign array_update_77884[9] = add_77421 == 32'h0000_0009 ? array_update_77882 : array_update_77871[9];
  assign array_index_77886 = array_update_72021[add_77883 > 32'h0000_0009 ? 4'h9 : add_77883[3:0]];
  assign array_index_77887 = array_update_77884[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_77891 = smul32b_32b_x_32b(array_index_77428[add_77883 > 32'h0000_0009 ? 4'h9 : add_77883[3:0]], array_index_77886[add_77829 > 32'h0000_0009 ? 4'h9 : add_77829[3:0]]);
  assign add_77893 = array_index_77887[add_77829 > 32'h0000_0009 ? 4'h9 : add_77829[3:0]] + smul_77891;
  assign array_update_77895[0] = add_77829 == 32'h0000_0000 ? add_77893 : array_index_77887[0];
  assign array_update_77895[1] = add_77829 == 32'h0000_0001 ? add_77893 : array_index_77887[1];
  assign array_update_77895[2] = add_77829 == 32'h0000_0002 ? add_77893 : array_index_77887[2];
  assign array_update_77895[3] = add_77829 == 32'h0000_0003 ? add_77893 : array_index_77887[3];
  assign array_update_77895[4] = add_77829 == 32'h0000_0004 ? add_77893 : array_index_77887[4];
  assign array_update_77895[5] = add_77829 == 32'h0000_0005 ? add_77893 : array_index_77887[5];
  assign array_update_77895[6] = add_77829 == 32'h0000_0006 ? add_77893 : array_index_77887[6];
  assign array_update_77895[7] = add_77829 == 32'h0000_0007 ? add_77893 : array_index_77887[7];
  assign array_update_77895[8] = add_77829 == 32'h0000_0008 ? add_77893 : array_index_77887[8];
  assign array_update_77895[9] = add_77829 == 32'h0000_0009 ? add_77893 : array_index_77887[9];
  assign add_77896 = add_77883 + 32'h0000_0001;
  assign array_update_77897[0] = add_77421 == 32'h0000_0000 ? array_update_77895 : array_update_77884[0];
  assign array_update_77897[1] = add_77421 == 32'h0000_0001 ? array_update_77895 : array_update_77884[1];
  assign array_update_77897[2] = add_77421 == 32'h0000_0002 ? array_update_77895 : array_update_77884[2];
  assign array_update_77897[3] = add_77421 == 32'h0000_0003 ? array_update_77895 : array_update_77884[3];
  assign array_update_77897[4] = add_77421 == 32'h0000_0004 ? array_update_77895 : array_update_77884[4];
  assign array_update_77897[5] = add_77421 == 32'h0000_0005 ? array_update_77895 : array_update_77884[5];
  assign array_update_77897[6] = add_77421 == 32'h0000_0006 ? array_update_77895 : array_update_77884[6];
  assign array_update_77897[7] = add_77421 == 32'h0000_0007 ? array_update_77895 : array_update_77884[7];
  assign array_update_77897[8] = add_77421 == 32'h0000_0008 ? array_update_77895 : array_update_77884[8];
  assign array_update_77897[9] = add_77421 == 32'h0000_0009 ? array_update_77895 : array_update_77884[9];
  assign array_index_77899 = array_update_72021[add_77896 > 32'h0000_0009 ? 4'h9 : add_77896[3:0]];
  assign array_index_77900 = array_update_77897[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_77904 = smul32b_32b_x_32b(array_index_77428[add_77896 > 32'h0000_0009 ? 4'h9 : add_77896[3:0]], array_index_77899[add_77829 > 32'h0000_0009 ? 4'h9 : add_77829[3:0]]);
  assign add_77906 = array_index_77900[add_77829 > 32'h0000_0009 ? 4'h9 : add_77829[3:0]] + smul_77904;
  assign array_update_77908[0] = add_77829 == 32'h0000_0000 ? add_77906 : array_index_77900[0];
  assign array_update_77908[1] = add_77829 == 32'h0000_0001 ? add_77906 : array_index_77900[1];
  assign array_update_77908[2] = add_77829 == 32'h0000_0002 ? add_77906 : array_index_77900[2];
  assign array_update_77908[3] = add_77829 == 32'h0000_0003 ? add_77906 : array_index_77900[3];
  assign array_update_77908[4] = add_77829 == 32'h0000_0004 ? add_77906 : array_index_77900[4];
  assign array_update_77908[5] = add_77829 == 32'h0000_0005 ? add_77906 : array_index_77900[5];
  assign array_update_77908[6] = add_77829 == 32'h0000_0006 ? add_77906 : array_index_77900[6];
  assign array_update_77908[7] = add_77829 == 32'h0000_0007 ? add_77906 : array_index_77900[7];
  assign array_update_77908[8] = add_77829 == 32'h0000_0008 ? add_77906 : array_index_77900[8];
  assign array_update_77908[9] = add_77829 == 32'h0000_0009 ? add_77906 : array_index_77900[9];
  assign add_77909 = add_77896 + 32'h0000_0001;
  assign array_update_77910[0] = add_77421 == 32'h0000_0000 ? array_update_77908 : array_update_77897[0];
  assign array_update_77910[1] = add_77421 == 32'h0000_0001 ? array_update_77908 : array_update_77897[1];
  assign array_update_77910[2] = add_77421 == 32'h0000_0002 ? array_update_77908 : array_update_77897[2];
  assign array_update_77910[3] = add_77421 == 32'h0000_0003 ? array_update_77908 : array_update_77897[3];
  assign array_update_77910[4] = add_77421 == 32'h0000_0004 ? array_update_77908 : array_update_77897[4];
  assign array_update_77910[5] = add_77421 == 32'h0000_0005 ? array_update_77908 : array_update_77897[5];
  assign array_update_77910[6] = add_77421 == 32'h0000_0006 ? array_update_77908 : array_update_77897[6];
  assign array_update_77910[7] = add_77421 == 32'h0000_0007 ? array_update_77908 : array_update_77897[7];
  assign array_update_77910[8] = add_77421 == 32'h0000_0008 ? array_update_77908 : array_update_77897[8];
  assign array_update_77910[9] = add_77421 == 32'h0000_0009 ? array_update_77908 : array_update_77897[9];
  assign array_index_77912 = array_update_72021[add_77909 > 32'h0000_0009 ? 4'h9 : add_77909[3:0]];
  assign array_index_77913 = array_update_77910[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_77917 = smul32b_32b_x_32b(array_index_77428[add_77909 > 32'h0000_0009 ? 4'h9 : add_77909[3:0]], array_index_77912[add_77829 > 32'h0000_0009 ? 4'h9 : add_77829[3:0]]);
  assign add_77919 = array_index_77913[add_77829 > 32'h0000_0009 ? 4'h9 : add_77829[3:0]] + smul_77917;
  assign array_update_77921[0] = add_77829 == 32'h0000_0000 ? add_77919 : array_index_77913[0];
  assign array_update_77921[1] = add_77829 == 32'h0000_0001 ? add_77919 : array_index_77913[1];
  assign array_update_77921[2] = add_77829 == 32'h0000_0002 ? add_77919 : array_index_77913[2];
  assign array_update_77921[3] = add_77829 == 32'h0000_0003 ? add_77919 : array_index_77913[3];
  assign array_update_77921[4] = add_77829 == 32'h0000_0004 ? add_77919 : array_index_77913[4];
  assign array_update_77921[5] = add_77829 == 32'h0000_0005 ? add_77919 : array_index_77913[5];
  assign array_update_77921[6] = add_77829 == 32'h0000_0006 ? add_77919 : array_index_77913[6];
  assign array_update_77921[7] = add_77829 == 32'h0000_0007 ? add_77919 : array_index_77913[7];
  assign array_update_77921[8] = add_77829 == 32'h0000_0008 ? add_77919 : array_index_77913[8];
  assign array_update_77921[9] = add_77829 == 32'h0000_0009 ? add_77919 : array_index_77913[9];
  assign add_77922 = add_77909 + 32'h0000_0001;
  assign array_update_77923[0] = add_77421 == 32'h0000_0000 ? array_update_77921 : array_update_77910[0];
  assign array_update_77923[1] = add_77421 == 32'h0000_0001 ? array_update_77921 : array_update_77910[1];
  assign array_update_77923[2] = add_77421 == 32'h0000_0002 ? array_update_77921 : array_update_77910[2];
  assign array_update_77923[3] = add_77421 == 32'h0000_0003 ? array_update_77921 : array_update_77910[3];
  assign array_update_77923[4] = add_77421 == 32'h0000_0004 ? array_update_77921 : array_update_77910[4];
  assign array_update_77923[5] = add_77421 == 32'h0000_0005 ? array_update_77921 : array_update_77910[5];
  assign array_update_77923[6] = add_77421 == 32'h0000_0006 ? array_update_77921 : array_update_77910[6];
  assign array_update_77923[7] = add_77421 == 32'h0000_0007 ? array_update_77921 : array_update_77910[7];
  assign array_update_77923[8] = add_77421 == 32'h0000_0008 ? array_update_77921 : array_update_77910[8];
  assign array_update_77923[9] = add_77421 == 32'h0000_0009 ? array_update_77921 : array_update_77910[9];
  assign array_index_77925 = array_update_72021[add_77922 > 32'h0000_0009 ? 4'h9 : add_77922[3:0]];
  assign array_index_77926 = array_update_77923[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_77930 = smul32b_32b_x_32b(array_index_77428[add_77922 > 32'h0000_0009 ? 4'h9 : add_77922[3:0]], array_index_77925[add_77829 > 32'h0000_0009 ? 4'h9 : add_77829[3:0]]);
  assign add_77932 = array_index_77926[add_77829 > 32'h0000_0009 ? 4'h9 : add_77829[3:0]] + smul_77930;
  assign array_update_77934[0] = add_77829 == 32'h0000_0000 ? add_77932 : array_index_77926[0];
  assign array_update_77934[1] = add_77829 == 32'h0000_0001 ? add_77932 : array_index_77926[1];
  assign array_update_77934[2] = add_77829 == 32'h0000_0002 ? add_77932 : array_index_77926[2];
  assign array_update_77934[3] = add_77829 == 32'h0000_0003 ? add_77932 : array_index_77926[3];
  assign array_update_77934[4] = add_77829 == 32'h0000_0004 ? add_77932 : array_index_77926[4];
  assign array_update_77934[5] = add_77829 == 32'h0000_0005 ? add_77932 : array_index_77926[5];
  assign array_update_77934[6] = add_77829 == 32'h0000_0006 ? add_77932 : array_index_77926[6];
  assign array_update_77934[7] = add_77829 == 32'h0000_0007 ? add_77932 : array_index_77926[7];
  assign array_update_77934[8] = add_77829 == 32'h0000_0008 ? add_77932 : array_index_77926[8];
  assign array_update_77934[9] = add_77829 == 32'h0000_0009 ? add_77932 : array_index_77926[9];
  assign add_77935 = add_77922 + 32'h0000_0001;
  assign array_update_77936[0] = add_77421 == 32'h0000_0000 ? array_update_77934 : array_update_77923[0];
  assign array_update_77936[1] = add_77421 == 32'h0000_0001 ? array_update_77934 : array_update_77923[1];
  assign array_update_77936[2] = add_77421 == 32'h0000_0002 ? array_update_77934 : array_update_77923[2];
  assign array_update_77936[3] = add_77421 == 32'h0000_0003 ? array_update_77934 : array_update_77923[3];
  assign array_update_77936[4] = add_77421 == 32'h0000_0004 ? array_update_77934 : array_update_77923[4];
  assign array_update_77936[5] = add_77421 == 32'h0000_0005 ? array_update_77934 : array_update_77923[5];
  assign array_update_77936[6] = add_77421 == 32'h0000_0006 ? array_update_77934 : array_update_77923[6];
  assign array_update_77936[7] = add_77421 == 32'h0000_0007 ? array_update_77934 : array_update_77923[7];
  assign array_update_77936[8] = add_77421 == 32'h0000_0008 ? array_update_77934 : array_update_77923[8];
  assign array_update_77936[9] = add_77421 == 32'h0000_0009 ? array_update_77934 : array_update_77923[9];
  assign array_index_77938 = array_update_72021[add_77935 > 32'h0000_0009 ? 4'h9 : add_77935[3:0]];
  assign array_index_77939 = array_update_77936[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_77943 = smul32b_32b_x_32b(array_index_77428[add_77935 > 32'h0000_0009 ? 4'h9 : add_77935[3:0]], array_index_77938[add_77829 > 32'h0000_0009 ? 4'h9 : add_77829[3:0]]);
  assign add_77945 = array_index_77939[add_77829 > 32'h0000_0009 ? 4'h9 : add_77829[3:0]] + smul_77943;
  assign array_update_77947[0] = add_77829 == 32'h0000_0000 ? add_77945 : array_index_77939[0];
  assign array_update_77947[1] = add_77829 == 32'h0000_0001 ? add_77945 : array_index_77939[1];
  assign array_update_77947[2] = add_77829 == 32'h0000_0002 ? add_77945 : array_index_77939[2];
  assign array_update_77947[3] = add_77829 == 32'h0000_0003 ? add_77945 : array_index_77939[3];
  assign array_update_77947[4] = add_77829 == 32'h0000_0004 ? add_77945 : array_index_77939[4];
  assign array_update_77947[5] = add_77829 == 32'h0000_0005 ? add_77945 : array_index_77939[5];
  assign array_update_77947[6] = add_77829 == 32'h0000_0006 ? add_77945 : array_index_77939[6];
  assign array_update_77947[7] = add_77829 == 32'h0000_0007 ? add_77945 : array_index_77939[7];
  assign array_update_77947[8] = add_77829 == 32'h0000_0008 ? add_77945 : array_index_77939[8];
  assign array_update_77947[9] = add_77829 == 32'h0000_0009 ? add_77945 : array_index_77939[9];
  assign add_77948 = add_77935 + 32'h0000_0001;
  assign array_update_77949[0] = add_77421 == 32'h0000_0000 ? array_update_77947 : array_update_77936[0];
  assign array_update_77949[1] = add_77421 == 32'h0000_0001 ? array_update_77947 : array_update_77936[1];
  assign array_update_77949[2] = add_77421 == 32'h0000_0002 ? array_update_77947 : array_update_77936[2];
  assign array_update_77949[3] = add_77421 == 32'h0000_0003 ? array_update_77947 : array_update_77936[3];
  assign array_update_77949[4] = add_77421 == 32'h0000_0004 ? array_update_77947 : array_update_77936[4];
  assign array_update_77949[5] = add_77421 == 32'h0000_0005 ? array_update_77947 : array_update_77936[5];
  assign array_update_77949[6] = add_77421 == 32'h0000_0006 ? array_update_77947 : array_update_77936[6];
  assign array_update_77949[7] = add_77421 == 32'h0000_0007 ? array_update_77947 : array_update_77936[7];
  assign array_update_77949[8] = add_77421 == 32'h0000_0008 ? array_update_77947 : array_update_77936[8];
  assign array_update_77949[9] = add_77421 == 32'h0000_0009 ? array_update_77947 : array_update_77936[9];
  assign array_index_77951 = array_update_72021[add_77948 > 32'h0000_0009 ? 4'h9 : add_77948[3:0]];
  assign array_index_77952 = array_update_77949[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_77956 = smul32b_32b_x_32b(array_index_77428[add_77948 > 32'h0000_0009 ? 4'h9 : add_77948[3:0]], array_index_77951[add_77829 > 32'h0000_0009 ? 4'h9 : add_77829[3:0]]);
  assign add_77958 = array_index_77952[add_77829 > 32'h0000_0009 ? 4'h9 : add_77829[3:0]] + smul_77956;
  assign array_update_77959[0] = add_77829 == 32'h0000_0000 ? add_77958 : array_index_77952[0];
  assign array_update_77959[1] = add_77829 == 32'h0000_0001 ? add_77958 : array_index_77952[1];
  assign array_update_77959[2] = add_77829 == 32'h0000_0002 ? add_77958 : array_index_77952[2];
  assign array_update_77959[3] = add_77829 == 32'h0000_0003 ? add_77958 : array_index_77952[3];
  assign array_update_77959[4] = add_77829 == 32'h0000_0004 ? add_77958 : array_index_77952[4];
  assign array_update_77959[5] = add_77829 == 32'h0000_0005 ? add_77958 : array_index_77952[5];
  assign array_update_77959[6] = add_77829 == 32'h0000_0006 ? add_77958 : array_index_77952[6];
  assign array_update_77959[7] = add_77829 == 32'h0000_0007 ? add_77958 : array_index_77952[7];
  assign array_update_77959[8] = add_77829 == 32'h0000_0008 ? add_77958 : array_index_77952[8];
  assign array_update_77959[9] = add_77829 == 32'h0000_0009 ? add_77958 : array_index_77952[9];
  assign array_update_77960[0] = add_77421 == 32'h0000_0000 ? array_update_77959 : array_update_77949[0];
  assign array_update_77960[1] = add_77421 == 32'h0000_0001 ? array_update_77959 : array_update_77949[1];
  assign array_update_77960[2] = add_77421 == 32'h0000_0002 ? array_update_77959 : array_update_77949[2];
  assign array_update_77960[3] = add_77421 == 32'h0000_0003 ? array_update_77959 : array_update_77949[3];
  assign array_update_77960[4] = add_77421 == 32'h0000_0004 ? array_update_77959 : array_update_77949[4];
  assign array_update_77960[5] = add_77421 == 32'h0000_0005 ? array_update_77959 : array_update_77949[5];
  assign array_update_77960[6] = add_77421 == 32'h0000_0006 ? array_update_77959 : array_update_77949[6];
  assign array_update_77960[7] = add_77421 == 32'h0000_0007 ? array_update_77959 : array_update_77949[7];
  assign array_update_77960[8] = add_77421 == 32'h0000_0008 ? array_update_77959 : array_update_77949[8];
  assign array_update_77960[9] = add_77421 == 32'h0000_0009 ? array_update_77959 : array_update_77949[9];
  assign array_index_77962 = array_update_77960[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign add_77964 = add_77829 + 32'h0000_0001;
  assign array_update_77965[0] = add_77964 == 32'h0000_0000 ? 32'h0000_0000 : array_index_77962[0];
  assign array_update_77965[1] = add_77964 == 32'h0000_0001 ? 32'h0000_0000 : array_index_77962[1];
  assign array_update_77965[2] = add_77964 == 32'h0000_0002 ? 32'h0000_0000 : array_index_77962[2];
  assign array_update_77965[3] = add_77964 == 32'h0000_0003 ? 32'h0000_0000 : array_index_77962[3];
  assign array_update_77965[4] = add_77964 == 32'h0000_0004 ? 32'h0000_0000 : array_index_77962[4];
  assign array_update_77965[5] = add_77964 == 32'h0000_0005 ? 32'h0000_0000 : array_index_77962[5];
  assign array_update_77965[6] = add_77964 == 32'h0000_0006 ? 32'h0000_0000 : array_index_77962[6];
  assign array_update_77965[7] = add_77964 == 32'h0000_0007 ? 32'h0000_0000 : array_index_77962[7];
  assign array_update_77965[8] = add_77964 == 32'h0000_0008 ? 32'h0000_0000 : array_index_77962[8];
  assign array_update_77965[9] = add_77964 == 32'h0000_0009 ? 32'h0000_0000 : array_index_77962[9];
  assign literal_77966 = 32'h0000_0000;
  assign array_update_77967[0] = add_77421 == 32'h0000_0000 ? array_update_77965 : array_update_77960[0];
  assign array_update_77967[1] = add_77421 == 32'h0000_0001 ? array_update_77965 : array_update_77960[1];
  assign array_update_77967[2] = add_77421 == 32'h0000_0002 ? array_update_77965 : array_update_77960[2];
  assign array_update_77967[3] = add_77421 == 32'h0000_0003 ? array_update_77965 : array_update_77960[3];
  assign array_update_77967[4] = add_77421 == 32'h0000_0004 ? array_update_77965 : array_update_77960[4];
  assign array_update_77967[5] = add_77421 == 32'h0000_0005 ? array_update_77965 : array_update_77960[5];
  assign array_update_77967[6] = add_77421 == 32'h0000_0006 ? array_update_77965 : array_update_77960[6];
  assign array_update_77967[7] = add_77421 == 32'h0000_0007 ? array_update_77965 : array_update_77960[7];
  assign array_update_77967[8] = add_77421 == 32'h0000_0008 ? array_update_77965 : array_update_77960[8];
  assign array_update_77967[9] = add_77421 == 32'h0000_0009 ? array_update_77965 : array_update_77960[9];
  assign array_index_77969 = array_update_72021[literal_77966 > 32'h0000_0009 ? 4'h9 : literal_77966[3:0]];
  assign array_index_77970 = array_update_77967[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_77974 = smul32b_32b_x_32b(array_index_77428[literal_77966 > 32'h0000_0009 ? 4'h9 : literal_77966[3:0]], array_index_77969[add_77964 > 32'h0000_0009 ? 4'h9 : add_77964[3:0]]);
  assign add_77976 = array_index_77970[add_77964 > 32'h0000_0009 ? 4'h9 : add_77964[3:0]] + smul_77974;
  assign array_update_77978[0] = add_77964 == 32'h0000_0000 ? add_77976 : array_index_77970[0];
  assign array_update_77978[1] = add_77964 == 32'h0000_0001 ? add_77976 : array_index_77970[1];
  assign array_update_77978[2] = add_77964 == 32'h0000_0002 ? add_77976 : array_index_77970[2];
  assign array_update_77978[3] = add_77964 == 32'h0000_0003 ? add_77976 : array_index_77970[3];
  assign array_update_77978[4] = add_77964 == 32'h0000_0004 ? add_77976 : array_index_77970[4];
  assign array_update_77978[5] = add_77964 == 32'h0000_0005 ? add_77976 : array_index_77970[5];
  assign array_update_77978[6] = add_77964 == 32'h0000_0006 ? add_77976 : array_index_77970[6];
  assign array_update_77978[7] = add_77964 == 32'h0000_0007 ? add_77976 : array_index_77970[7];
  assign array_update_77978[8] = add_77964 == 32'h0000_0008 ? add_77976 : array_index_77970[8];
  assign array_update_77978[9] = add_77964 == 32'h0000_0009 ? add_77976 : array_index_77970[9];
  assign add_77979 = literal_77966 + 32'h0000_0001;
  assign array_update_77980[0] = add_77421 == 32'h0000_0000 ? array_update_77978 : array_update_77967[0];
  assign array_update_77980[1] = add_77421 == 32'h0000_0001 ? array_update_77978 : array_update_77967[1];
  assign array_update_77980[2] = add_77421 == 32'h0000_0002 ? array_update_77978 : array_update_77967[2];
  assign array_update_77980[3] = add_77421 == 32'h0000_0003 ? array_update_77978 : array_update_77967[3];
  assign array_update_77980[4] = add_77421 == 32'h0000_0004 ? array_update_77978 : array_update_77967[4];
  assign array_update_77980[5] = add_77421 == 32'h0000_0005 ? array_update_77978 : array_update_77967[5];
  assign array_update_77980[6] = add_77421 == 32'h0000_0006 ? array_update_77978 : array_update_77967[6];
  assign array_update_77980[7] = add_77421 == 32'h0000_0007 ? array_update_77978 : array_update_77967[7];
  assign array_update_77980[8] = add_77421 == 32'h0000_0008 ? array_update_77978 : array_update_77967[8];
  assign array_update_77980[9] = add_77421 == 32'h0000_0009 ? array_update_77978 : array_update_77967[9];
  assign array_index_77982 = array_update_72021[add_77979 > 32'h0000_0009 ? 4'h9 : add_77979[3:0]];
  assign array_index_77983 = array_update_77980[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_77987 = smul32b_32b_x_32b(array_index_77428[add_77979 > 32'h0000_0009 ? 4'h9 : add_77979[3:0]], array_index_77982[add_77964 > 32'h0000_0009 ? 4'h9 : add_77964[3:0]]);
  assign add_77989 = array_index_77983[add_77964 > 32'h0000_0009 ? 4'h9 : add_77964[3:0]] + smul_77987;
  assign array_update_77991[0] = add_77964 == 32'h0000_0000 ? add_77989 : array_index_77983[0];
  assign array_update_77991[1] = add_77964 == 32'h0000_0001 ? add_77989 : array_index_77983[1];
  assign array_update_77991[2] = add_77964 == 32'h0000_0002 ? add_77989 : array_index_77983[2];
  assign array_update_77991[3] = add_77964 == 32'h0000_0003 ? add_77989 : array_index_77983[3];
  assign array_update_77991[4] = add_77964 == 32'h0000_0004 ? add_77989 : array_index_77983[4];
  assign array_update_77991[5] = add_77964 == 32'h0000_0005 ? add_77989 : array_index_77983[5];
  assign array_update_77991[6] = add_77964 == 32'h0000_0006 ? add_77989 : array_index_77983[6];
  assign array_update_77991[7] = add_77964 == 32'h0000_0007 ? add_77989 : array_index_77983[7];
  assign array_update_77991[8] = add_77964 == 32'h0000_0008 ? add_77989 : array_index_77983[8];
  assign array_update_77991[9] = add_77964 == 32'h0000_0009 ? add_77989 : array_index_77983[9];
  assign add_77992 = add_77979 + 32'h0000_0001;
  assign array_update_77993[0] = add_77421 == 32'h0000_0000 ? array_update_77991 : array_update_77980[0];
  assign array_update_77993[1] = add_77421 == 32'h0000_0001 ? array_update_77991 : array_update_77980[1];
  assign array_update_77993[2] = add_77421 == 32'h0000_0002 ? array_update_77991 : array_update_77980[2];
  assign array_update_77993[3] = add_77421 == 32'h0000_0003 ? array_update_77991 : array_update_77980[3];
  assign array_update_77993[4] = add_77421 == 32'h0000_0004 ? array_update_77991 : array_update_77980[4];
  assign array_update_77993[5] = add_77421 == 32'h0000_0005 ? array_update_77991 : array_update_77980[5];
  assign array_update_77993[6] = add_77421 == 32'h0000_0006 ? array_update_77991 : array_update_77980[6];
  assign array_update_77993[7] = add_77421 == 32'h0000_0007 ? array_update_77991 : array_update_77980[7];
  assign array_update_77993[8] = add_77421 == 32'h0000_0008 ? array_update_77991 : array_update_77980[8];
  assign array_update_77993[9] = add_77421 == 32'h0000_0009 ? array_update_77991 : array_update_77980[9];
  assign array_index_77995 = array_update_72021[add_77992 > 32'h0000_0009 ? 4'h9 : add_77992[3:0]];
  assign array_index_77996 = array_update_77993[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_78000 = smul32b_32b_x_32b(array_index_77428[add_77992 > 32'h0000_0009 ? 4'h9 : add_77992[3:0]], array_index_77995[add_77964 > 32'h0000_0009 ? 4'h9 : add_77964[3:0]]);
  assign add_78002 = array_index_77996[add_77964 > 32'h0000_0009 ? 4'h9 : add_77964[3:0]] + smul_78000;
  assign array_update_78004[0] = add_77964 == 32'h0000_0000 ? add_78002 : array_index_77996[0];
  assign array_update_78004[1] = add_77964 == 32'h0000_0001 ? add_78002 : array_index_77996[1];
  assign array_update_78004[2] = add_77964 == 32'h0000_0002 ? add_78002 : array_index_77996[2];
  assign array_update_78004[3] = add_77964 == 32'h0000_0003 ? add_78002 : array_index_77996[3];
  assign array_update_78004[4] = add_77964 == 32'h0000_0004 ? add_78002 : array_index_77996[4];
  assign array_update_78004[5] = add_77964 == 32'h0000_0005 ? add_78002 : array_index_77996[5];
  assign array_update_78004[6] = add_77964 == 32'h0000_0006 ? add_78002 : array_index_77996[6];
  assign array_update_78004[7] = add_77964 == 32'h0000_0007 ? add_78002 : array_index_77996[7];
  assign array_update_78004[8] = add_77964 == 32'h0000_0008 ? add_78002 : array_index_77996[8];
  assign array_update_78004[9] = add_77964 == 32'h0000_0009 ? add_78002 : array_index_77996[9];
  assign add_78005 = add_77992 + 32'h0000_0001;
  assign array_update_78006[0] = add_77421 == 32'h0000_0000 ? array_update_78004 : array_update_77993[0];
  assign array_update_78006[1] = add_77421 == 32'h0000_0001 ? array_update_78004 : array_update_77993[1];
  assign array_update_78006[2] = add_77421 == 32'h0000_0002 ? array_update_78004 : array_update_77993[2];
  assign array_update_78006[3] = add_77421 == 32'h0000_0003 ? array_update_78004 : array_update_77993[3];
  assign array_update_78006[4] = add_77421 == 32'h0000_0004 ? array_update_78004 : array_update_77993[4];
  assign array_update_78006[5] = add_77421 == 32'h0000_0005 ? array_update_78004 : array_update_77993[5];
  assign array_update_78006[6] = add_77421 == 32'h0000_0006 ? array_update_78004 : array_update_77993[6];
  assign array_update_78006[7] = add_77421 == 32'h0000_0007 ? array_update_78004 : array_update_77993[7];
  assign array_update_78006[8] = add_77421 == 32'h0000_0008 ? array_update_78004 : array_update_77993[8];
  assign array_update_78006[9] = add_77421 == 32'h0000_0009 ? array_update_78004 : array_update_77993[9];
  assign array_index_78008 = array_update_72021[add_78005 > 32'h0000_0009 ? 4'h9 : add_78005[3:0]];
  assign array_index_78009 = array_update_78006[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_78013 = smul32b_32b_x_32b(array_index_77428[add_78005 > 32'h0000_0009 ? 4'h9 : add_78005[3:0]], array_index_78008[add_77964 > 32'h0000_0009 ? 4'h9 : add_77964[3:0]]);
  assign add_78015 = array_index_78009[add_77964 > 32'h0000_0009 ? 4'h9 : add_77964[3:0]] + smul_78013;
  assign array_update_78017[0] = add_77964 == 32'h0000_0000 ? add_78015 : array_index_78009[0];
  assign array_update_78017[1] = add_77964 == 32'h0000_0001 ? add_78015 : array_index_78009[1];
  assign array_update_78017[2] = add_77964 == 32'h0000_0002 ? add_78015 : array_index_78009[2];
  assign array_update_78017[3] = add_77964 == 32'h0000_0003 ? add_78015 : array_index_78009[3];
  assign array_update_78017[4] = add_77964 == 32'h0000_0004 ? add_78015 : array_index_78009[4];
  assign array_update_78017[5] = add_77964 == 32'h0000_0005 ? add_78015 : array_index_78009[5];
  assign array_update_78017[6] = add_77964 == 32'h0000_0006 ? add_78015 : array_index_78009[6];
  assign array_update_78017[7] = add_77964 == 32'h0000_0007 ? add_78015 : array_index_78009[7];
  assign array_update_78017[8] = add_77964 == 32'h0000_0008 ? add_78015 : array_index_78009[8];
  assign array_update_78017[9] = add_77964 == 32'h0000_0009 ? add_78015 : array_index_78009[9];
  assign add_78018 = add_78005 + 32'h0000_0001;
  assign array_update_78019[0] = add_77421 == 32'h0000_0000 ? array_update_78017 : array_update_78006[0];
  assign array_update_78019[1] = add_77421 == 32'h0000_0001 ? array_update_78017 : array_update_78006[1];
  assign array_update_78019[2] = add_77421 == 32'h0000_0002 ? array_update_78017 : array_update_78006[2];
  assign array_update_78019[3] = add_77421 == 32'h0000_0003 ? array_update_78017 : array_update_78006[3];
  assign array_update_78019[4] = add_77421 == 32'h0000_0004 ? array_update_78017 : array_update_78006[4];
  assign array_update_78019[5] = add_77421 == 32'h0000_0005 ? array_update_78017 : array_update_78006[5];
  assign array_update_78019[6] = add_77421 == 32'h0000_0006 ? array_update_78017 : array_update_78006[6];
  assign array_update_78019[7] = add_77421 == 32'h0000_0007 ? array_update_78017 : array_update_78006[7];
  assign array_update_78019[8] = add_77421 == 32'h0000_0008 ? array_update_78017 : array_update_78006[8];
  assign array_update_78019[9] = add_77421 == 32'h0000_0009 ? array_update_78017 : array_update_78006[9];
  assign array_index_78021 = array_update_72021[add_78018 > 32'h0000_0009 ? 4'h9 : add_78018[3:0]];
  assign array_index_78022 = array_update_78019[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_78026 = smul32b_32b_x_32b(array_index_77428[add_78018 > 32'h0000_0009 ? 4'h9 : add_78018[3:0]], array_index_78021[add_77964 > 32'h0000_0009 ? 4'h9 : add_77964[3:0]]);
  assign add_78028 = array_index_78022[add_77964 > 32'h0000_0009 ? 4'h9 : add_77964[3:0]] + smul_78026;
  assign array_update_78030[0] = add_77964 == 32'h0000_0000 ? add_78028 : array_index_78022[0];
  assign array_update_78030[1] = add_77964 == 32'h0000_0001 ? add_78028 : array_index_78022[1];
  assign array_update_78030[2] = add_77964 == 32'h0000_0002 ? add_78028 : array_index_78022[2];
  assign array_update_78030[3] = add_77964 == 32'h0000_0003 ? add_78028 : array_index_78022[3];
  assign array_update_78030[4] = add_77964 == 32'h0000_0004 ? add_78028 : array_index_78022[4];
  assign array_update_78030[5] = add_77964 == 32'h0000_0005 ? add_78028 : array_index_78022[5];
  assign array_update_78030[6] = add_77964 == 32'h0000_0006 ? add_78028 : array_index_78022[6];
  assign array_update_78030[7] = add_77964 == 32'h0000_0007 ? add_78028 : array_index_78022[7];
  assign array_update_78030[8] = add_77964 == 32'h0000_0008 ? add_78028 : array_index_78022[8];
  assign array_update_78030[9] = add_77964 == 32'h0000_0009 ? add_78028 : array_index_78022[9];
  assign add_78031 = add_78018 + 32'h0000_0001;
  assign array_update_78032[0] = add_77421 == 32'h0000_0000 ? array_update_78030 : array_update_78019[0];
  assign array_update_78032[1] = add_77421 == 32'h0000_0001 ? array_update_78030 : array_update_78019[1];
  assign array_update_78032[2] = add_77421 == 32'h0000_0002 ? array_update_78030 : array_update_78019[2];
  assign array_update_78032[3] = add_77421 == 32'h0000_0003 ? array_update_78030 : array_update_78019[3];
  assign array_update_78032[4] = add_77421 == 32'h0000_0004 ? array_update_78030 : array_update_78019[4];
  assign array_update_78032[5] = add_77421 == 32'h0000_0005 ? array_update_78030 : array_update_78019[5];
  assign array_update_78032[6] = add_77421 == 32'h0000_0006 ? array_update_78030 : array_update_78019[6];
  assign array_update_78032[7] = add_77421 == 32'h0000_0007 ? array_update_78030 : array_update_78019[7];
  assign array_update_78032[8] = add_77421 == 32'h0000_0008 ? array_update_78030 : array_update_78019[8];
  assign array_update_78032[9] = add_77421 == 32'h0000_0009 ? array_update_78030 : array_update_78019[9];
  assign array_index_78034 = array_update_72021[add_78031 > 32'h0000_0009 ? 4'h9 : add_78031[3:0]];
  assign array_index_78035 = array_update_78032[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_78039 = smul32b_32b_x_32b(array_index_77428[add_78031 > 32'h0000_0009 ? 4'h9 : add_78031[3:0]], array_index_78034[add_77964 > 32'h0000_0009 ? 4'h9 : add_77964[3:0]]);
  assign add_78041 = array_index_78035[add_77964 > 32'h0000_0009 ? 4'h9 : add_77964[3:0]] + smul_78039;
  assign array_update_78043[0] = add_77964 == 32'h0000_0000 ? add_78041 : array_index_78035[0];
  assign array_update_78043[1] = add_77964 == 32'h0000_0001 ? add_78041 : array_index_78035[1];
  assign array_update_78043[2] = add_77964 == 32'h0000_0002 ? add_78041 : array_index_78035[2];
  assign array_update_78043[3] = add_77964 == 32'h0000_0003 ? add_78041 : array_index_78035[3];
  assign array_update_78043[4] = add_77964 == 32'h0000_0004 ? add_78041 : array_index_78035[4];
  assign array_update_78043[5] = add_77964 == 32'h0000_0005 ? add_78041 : array_index_78035[5];
  assign array_update_78043[6] = add_77964 == 32'h0000_0006 ? add_78041 : array_index_78035[6];
  assign array_update_78043[7] = add_77964 == 32'h0000_0007 ? add_78041 : array_index_78035[7];
  assign array_update_78043[8] = add_77964 == 32'h0000_0008 ? add_78041 : array_index_78035[8];
  assign array_update_78043[9] = add_77964 == 32'h0000_0009 ? add_78041 : array_index_78035[9];
  assign add_78044 = add_78031 + 32'h0000_0001;
  assign array_update_78045[0] = add_77421 == 32'h0000_0000 ? array_update_78043 : array_update_78032[0];
  assign array_update_78045[1] = add_77421 == 32'h0000_0001 ? array_update_78043 : array_update_78032[1];
  assign array_update_78045[2] = add_77421 == 32'h0000_0002 ? array_update_78043 : array_update_78032[2];
  assign array_update_78045[3] = add_77421 == 32'h0000_0003 ? array_update_78043 : array_update_78032[3];
  assign array_update_78045[4] = add_77421 == 32'h0000_0004 ? array_update_78043 : array_update_78032[4];
  assign array_update_78045[5] = add_77421 == 32'h0000_0005 ? array_update_78043 : array_update_78032[5];
  assign array_update_78045[6] = add_77421 == 32'h0000_0006 ? array_update_78043 : array_update_78032[6];
  assign array_update_78045[7] = add_77421 == 32'h0000_0007 ? array_update_78043 : array_update_78032[7];
  assign array_update_78045[8] = add_77421 == 32'h0000_0008 ? array_update_78043 : array_update_78032[8];
  assign array_update_78045[9] = add_77421 == 32'h0000_0009 ? array_update_78043 : array_update_78032[9];
  assign array_index_78047 = array_update_72021[add_78044 > 32'h0000_0009 ? 4'h9 : add_78044[3:0]];
  assign array_index_78048 = array_update_78045[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_78052 = smul32b_32b_x_32b(array_index_77428[add_78044 > 32'h0000_0009 ? 4'h9 : add_78044[3:0]], array_index_78047[add_77964 > 32'h0000_0009 ? 4'h9 : add_77964[3:0]]);
  assign add_78054 = array_index_78048[add_77964 > 32'h0000_0009 ? 4'h9 : add_77964[3:0]] + smul_78052;
  assign array_update_78056[0] = add_77964 == 32'h0000_0000 ? add_78054 : array_index_78048[0];
  assign array_update_78056[1] = add_77964 == 32'h0000_0001 ? add_78054 : array_index_78048[1];
  assign array_update_78056[2] = add_77964 == 32'h0000_0002 ? add_78054 : array_index_78048[2];
  assign array_update_78056[3] = add_77964 == 32'h0000_0003 ? add_78054 : array_index_78048[3];
  assign array_update_78056[4] = add_77964 == 32'h0000_0004 ? add_78054 : array_index_78048[4];
  assign array_update_78056[5] = add_77964 == 32'h0000_0005 ? add_78054 : array_index_78048[5];
  assign array_update_78056[6] = add_77964 == 32'h0000_0006 ? add_78054 : array_index_78048[6];
  assign array_update_78056[7] = add_77964 == 32'h0000_0007 ? add_78054 : array_index_78048[7];
  assign array_update_78056[8] = add_77964 == 32'h0000_0008 ? add_78054 : array_index_78048[8];
  assign array_update_78056[9] = add_77964 == 32'h0000_0009 ? add_78054 : array_index_78048[9];
  assign add_78057 = add_78044 + 32'h0000_0001;
  assign array_update_78058[0] = add_77421 == 32'h0000_0000 ? array_update_78056 : array_update_78045[0];
  assign array_update_78058[1] = add_77421 == 32'h0000_0001 ? array_update_78056 : array_update_78045[1];
  assign array_update_78058[2] = add_77421 == 32'h0000_0002 ? array_update_78056 : array_update_78045[2];
  assign array_update_78058[3] = add_77421 == 32'h0000_0003 ? array_update_78056 : array_update_78045[3];
  assign array_update_78058[4] = add_77421 == 32'h0000_0004 ? array_update_78056 : array_update_78045[4];
  assign array_update_78058[5] = add_77421 == 32'h0000_0005 ? array_update_78056 : array_update_78045[5];
  assign array_update_78058[6] = add_77421 == 32'h0000_0006 ? array_update_78056 : array_update_78045[6];
  assign array_update_78058[7] = add_77421 == 32'h0000_0007 ? array_update_78056 : array_update_78045[7];
  assign array_update_78058[8] = add_77421 == 32'h0000_0008 ? array_update_78056 : array_update_78045[8];
  assign array_update_78058[9] = add_77421 == 32'h0000_0009 ? array_update_78056 : array_update_78045[9];
  assign array_index_78060 = array_update_72021[add_78057 > 32'h0000_0009 ? 4'h9 : add_78057[3:0]];
  assign array_index_78061 = array_update_78058[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_78065 = smul32b_32b_x_32b(array_index_77428[add_78057 > 32'h0000_0009 ? 4'h9 : add_78057[3:0]], array_index_78060[add_77964 > 32'h0000_0009 ? 4'h9 : add_77964[3:0]]);
  assign add_78067 = array_index_78061[add_77964 > 32'h0000_0009 ? 4'h9 : add_77964[3:0]] + smul_78065;
  assign array_update_78069[0] = add_77964 == 32'h0000_0000 ? add_78067 : array_index_78061[0];
  assign array_update_78069[1] = add_77964 == 32'h0000_0001 ? add_78067 : array_index_78061[1];
  assign array_update_78069[2] = add_77964 == 32'h0000_0002 ? add_78067 : array_index_78061[2];
  assign array_update_78069[3] = add_77964 == 32'h0000_0003 ? add_78067 : array_index_78061[3];
  assign array_update_78069[4] = add_77964 == 32'h0000_0004 ? add_78067 : array_index_78061[4];
  assign array_update_78069[5] = add_77964 == 32'h0000_0005 ? add_78067 : array_index_78061[5];
  assign array_update_78069[6] = add_77964 == 32'h0000_0006 ? add_78067 : array_index_78061[6];
  assign array_update_78069[7] = add_77964 == 32'h0000_0007 ? add_78067 : array_index_78061[7];
  assign array_update_78069[8] = add_77964 == 32'h0000_0008 ? add_78067 : array_index_78061[8];
  assign array_update_78069[9] = add_77964 == 32'h0000_0009 ? add_78067 : array_index_78061[9];
  assign add_78070 = add_78057 + 32'h0000_0001;
  assign array_update_78071[0] = add_77421 == 32'h0000_0000 ? array_update_78069 : array_update_78058[0];
  assign array_update_78071[1] = add_77421 == 32'h0000_0001 ? array_update_78069 : array_update_78058[1];
  assign array_update_78071[2] = add_77421 == 32'h0000_0002 ? array_update_78069 : array_update_78058[2];
  assign array_update_78071[3] = add_77421 == 32'h0000_0003 ? array_update_78069 : array_update_78058[3];
  assign array_update_78071[4] = add_77421 == 32'h0000_0004 ? array_update_78069 : array_update_78058[4];
  assign array_update_78071[5] = add_77421 == 32'h0000_0005 ? array_update_78069 : array_update_78058[5];
  assign array_update_78071[6] = add_77421 == 32'h0000_0006 ? array_update_78069 : array_update_78058[6];
  assign array_update_78071[7] = add_77421 == 32'h0000_0007 ? array_update_78069 : array_update_78058[7];
  assign array_update_78071[8] = add_77421 == 32'h0000_0008 ? array_update_78069 : array_update_78058[8];
  assign array_update_78071[9] = add_77421 == 32'h0000_0009 ? array_update_78069 : array_update_78058[9];
  assign array_index_78073 = array_update_72021[add_78070 > 32'h0000_0009 ? 4'h9 : add_78070[3:0]];
  assign array_index_78074 = array_update_78071[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_78078 = smul32b_32b_x_32b(array_index_77428[add_78070 > 32'h0000_0009 ? 4'h9 : add_78070[3:0]], array_index_78073[add_77964 > 32'h0000_0009 ? 4'h9 : add_77964[3:0]]);
  assign add_78080 = array_index_78074[add_77964 > 32'h0000_0009 ? 4'h9 : add_77964[3:0]] + smul_78078;
  assign array_update_78082[0] = add_77964 == 32'h0000_0000 ? add_78080 : array_index_78074[0];
  assign array_update_78082[1] = add_77964 == 32'h0000_0001 ? add_78080 : array_index_78074[1];
  assign array_update_78082[2] = add_77964 == 32'h0000_0002 ? add_78080 : array_index_78074[2];
  assign array_update_78082[3] = add_77964 == 32'h0000_0003 ? add_78080 : array_index_78074[3];
  assign array_update_78082[4] = add_77964 == 32'h0000_0004 ? add_78080 : array_index_78074[4];
  assign array_update_78082[5] = add_77964 == 32'h0000_0005 ? add_78080 : array_index_78074[5];
  assign array_update_78082[6] = add_77964 == 32'h0000_0006 ? add_78080 : array_index_78074[6];
  assign array_update_78082[7] = add_77964 == 32'h0000_0007 ? add_78080 : array_index_78074[7];
  assign array_update_78082[8] = add_77964 == 32'h0000_0008 ? add_78080 : array_index_78074[8];
  assign array_update_78082[9] = add_77964 == 32'h0000_0009 ? add_78080 : array_index_78074[9];
  assign add_78083 = add_78070 + 32'h0000_0001;
  assign array_update_78084[0] = add_77421 == 32'h0000_0000 ? array_update_78082 : array_update_78071[0];
  assign array_update_78084[1] = add_77421 == 32'h0000_0001 ? array_update_78082 : array_update_78071[1];
  assign array_update_78084[2] = add_77421 == 32'h0000_0002 ? array_update_78082 : array_update_78071[2];
  assign array_update_78084[3] = add_77421 == 32'h0000_0003 ? array_update_78082 : array_update_78071[3];
  assign array_update_78084[4] = add_77421 == 32'h0000_0004 ? array_update_78082 : array_update_78071[4];
  assign array_update_78084[5] = add_77421 == 32'h0000_0005 ? array_update_78082 : array_update_78071[5];
  assign array_update_78084[6] = add_77421 == 32'h0000_0006 ? array_update_78082 : array_update_78071[6];
  assign array_update_78084[7] = add_77421 == 32'h0000_0007 ? array_update_78082 : array_update_78071[7];
  assign array_update_78084[8] = add_77421 == 32'h0000_0008 ? array_update_78082 : array_update_78071[8];
  assign array_update_78084[9] = add_77421 == 32'h0000_0009 ? array_update_78082 : array_update_78071[9];
  assign array_index_78086 = array_update_72021[add_78083 > 32'h0000_0009 ? 4'h9 : add_78083[3:0]];
  assign array_index_78087 = array_update_78084[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_78091 = smul32b_32b_x_32b(array_index_77428[add_78083 > 32'h0000_0009 ? 4'h9 : add_78083[3:0]], array_index_78086[add_77964 > 32'h0000_0009 ? 4'h9 : add_77964[3:0]]);
  assign add_78093 = array_index_78087[add_77964 > 32'h0000_0009 ? 4'h9 : add_77964[3:0]] + smul_78091;
  assign array_update_78094[0] = add_77964 == 32'h0000_0000 ? add_78093 : array_index_78087[0];
  assign array_update_78094[1] = add_77964 == 32'h0000_0001 ? add_78093 : array_index_78087[1];
  assign array_update_78094[2] = add_77964 == 32'h0000_0002 ? add_78093 : array_index_78087[2];
  assign array_update_78094[3] = add_77964 == 32'h0000_0003 ? add_78093 : array_index_78087[3];
  assign array_update_78094[4] = add_77964 == 32'h0000_0004 ? add_78093 : array_index_78087[4];
  assign array_update_78094[5] = add_77964 == 32'h0000_0005 ? add_78093 : array_index_78087[5];
  assign array_update_78094[6] = add_77964 == 32'h0000_0006 ? add_78093 : array_index_78087[6];
  assign array_update_78094[7] = add_77964 == 32'h0000_0007 ? add_78093 : array_index_78087[7];
  assign array_update_78094[8] = add_77964 == 32'h0000_0008 ? add_78093 : array_index_78087[8];
  assign array_update_78094[9] = add_77964 == 32'h0000_0009 ? add_78093 : array_index_78087[9];
  assign array_update_78095[0] = add_77421 == 32'h0000_0000 ? array_update_78094 : array_update_78084[0];
  assign array_update_78095[1] = add_77421 == 32'h0000_0001 ? array_update_78094 : array_update_78084[1];
  assign array_update_78095[2] = add_77421 == 32'h0000_0002 ? array_update_78094 : array_update_78084[2];
  assign array_update_78095[3] = add_77421 == 32'h0000_0003 ? array_update_78094 : array_update_78084[3];
  assign array_update_78095[4] = add_77421 == 32'h0000_0004 ? array_update_78094 : array_update_78084[4];
  assign array_update_78095[5] = add_77421 == 32'h0000_0005 ? array_update_78094 : array_update_78084[5];
  assign array_update_78095[6] = add_77421 == 32'h0000_0006 ? array_update_78094 : array_update_78084[6];
  assign array_update_78095[7] = add_77421 == 32'h0000_0007 ? array_update_78094 : array_update_78084[7];
  assign array_update_78095[8] = add_77421 == 32'h0000_0008 ? array_update_78094 : array_update_78084[8];
  assign array_update_78095[9] = add_77421 == 32'h0000_0009 ? array_update_78094 : array_update_78084[9];
  assign array_index_78097 = array_update_78095[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign add_78099 = add_77964 + 32'h0000_0001;
  assign array_update_78100[0] = add_78099 == 32'h0000_0000 ? 32'h0000_0000 : array_index_78097[0];
  assign array_update_78100[1] = add_78099 == 32'h0000_0001 ? 32'h0000_0000 : array_index_78097[1];
  assign array_update_78100[2] = add_78099 == 32'h0000_0002 ? 32'h0000_0000 : array_index_78097[2];
  assign array_update_78100[3] = add_78099 == 32'h0000_0003 ? 32'h0000_0000 : array_index_78097[3];
  assign array_update_78100[4] = add_78099 == 32'h0000_0004 ? 32'h0000_0000 : array_index_78097[4];
  assign array_update_78100[5] = add_78099 == 32'h0000_0005 ? 32'h0000_0000 : array_index_78097[5];
  assign array_update_78100[6] = add_78099 == 32'h0000_0006 ? 32'h0000_0000 : array_index_78097[6];
  assign array_update_78100[7] = add_78099 == 32'h0000_0007 ? 32'h0000_0000 : array_index_78097[7];
  assign array_update_78100[8] = add_78099 == 32'h0000_0008 ? 32'h0000_0000 : array_index_78097[8];
  assign array_update_78100[9] = add_78099 == 32'h0000_0009 ? 32'h0000_0000 : array_index_78097[9];
  assign literal_78101 = 32'h0000_0000;
  assign array_update_78102[0] = add_77421 == 32'h0000_0000 ? array_update_78100 : array_update_78095[0];
  assign array_update_78102[1] = add_77421 == 32'h0000_0001 ? array_update_78100 : array_update_78095[1];
  assign array_update_78102[2] = add_77421 == 32'h0000_0002 ? array_update_78100 : array_update_78095[2];
  assign array_update_78102[3] = add_77421 == 32'h0000_0003 ? array_update_78100 : array_update_78095[3];
  assign array_update_78102[4] = add_77421 == 32'h0000_0004 ? array_update_78100 : array_update_78095[4];
  assign array_update_78102[5] = add_77421 == 32'h0000_0005 ? array_update_78100 : array_update_78095[5];
  assign array_update_78102[6] = add_77421 == 32'h0000_0006 ? array_update_78100 : array_update_78095[6];
  assign array_update_78102[7] = add_77421 == 32'h0000_0007 ? array_update_78100 : array_update_78095[7];
  assign array_update_78102[8] = add_77421 == 32'h0000_0008 ? array_update_78100 : array_update_78095[8];
  assign array_update_78102[9] = add_77421 == 32'h0000_0009 ? array_update_78100 : array_update_78095[9];
  assign array_index_78104 = array_update_72021[literal_78101 > 32'h0000_0009 ? 4'h9 : literal_78101[3:0]];
  assign array_index_78105 = array_update_78102[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_78109 = smul32b_32b_x_32b(array_index_77428[literal_78101 > 32'h0000_0009 ? 4'h9 : literal_78101[3:0]], array_index_78104[add_78099 > 32'h0000_0009 ? 4'h9 : add_78099[3:0]]);
  assign add_78111 = array_index_78105[add_78099 > 32'h0000_0009 ? 4'h9 : add_78099[3:0]] + smul_78109;
  assign array_update_78113[0] = add_78099 == 32'h0000_0000 ? add_78111 : array_index_78105[0];
  assign array_update_78113[1] = add_78099 == 32'h0000_0001 ? add_78111 : array_index_78105[1];
  assign array_update_78113[2] = add_78099 == 32'h0000_0002 ? add_78111 : array_index_78105[2];
  assign array_update_78113[3] = add_78099 == 32'h0000_0003 ? add_78111 : array_index_78105[3];
  assign array_update_78113[4] = add_78099 == 32'h0000_0004 ? add_78111 : array_index_78105[4];
  assign array_update_78113[5] = add_78099 == 32'h0000_0005 ? add_78111 : array_index_78105[5];
  assign array_update_78113[6] = add_78099 == 32'h0000_0006 ? add_78111 : array_index_78105[6];
  assign array_update_78113[7] = add_78099 == 32'h0000_0007 ? add_78111 : array_index_78105[7];
  assign array_update_78113[8] = add_78099 == 32'h0000_0008 ? add_78111 : array_index_78105[8];
  assign array_update_78113[9] = add_78099 == 32'h0000_0009 ? add_78111 : array_index_78105[9];
  assign add_78114 = literal_78101 + 32'h0000_0001;
  assign array_update_78115[0] = add_77421 == 32'h0000_0000 ? array_update_78113 : array_update_78102[0];
  assign array_update_78115[1] = add_77421 == 32'h0000_0001 ? array_update_78113 : array_update_78102[1];
  assign array_update_78115[2] = add_77421 == 32'h0000_0002 ? array_update_78113 : array_update_78102[2];
  assign array_update_78115[3] = add_77421 == 32'h0000_0003 ? array_update_78113 : array_update_78102[3];
  assign array_update_78115[4] = add_77421 == 32'h0000_0004 ? array_update_78113 : array_update_78102[4];
  assign array_update_78115[5] = add_77421 == 32'h0000_0005 ? array_update_78113 : array_update_78102[5];
  assign array_update_78115[6] = add_77421 == 32'h0000_0006 ? array_update_78113 : array_update_78102[6];
  assign array_update_78115[7] = add_77421 == 32'h0000_0007 ? array_update_78113 : array_update_78102[7];
  assign array_update_78115[8] = add_77421 == 32'h0000_0008 ? array_update_78113 : array_update_78102[8];
  assign array_update_78115[9] = add_77421 == 32'h0000_0009 ? array_update_78113 : array_update_78102[9];
  assign array_index_78117 = array_update_72021[add_78114 > 32'h0000_0009 ? 4'h9 : add_78114[3:0]];
  assign array_index_78118 = array_update_78115[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_78122 = smul32b_32b_x_32b(array_index_77428[add_78114 > 32'h0000_0009 ? 4'h9 : add_78114[3:0]], array_index_78117[add_78099 > 32'h0000_0009 ? 4'h9 : add_78099[3:0]]);
  assign add_78124 = array_index_78118[add_78099 > 32'h0000_0009 ? 4'h9 : add_78099[3:0]] + smul_78122;
  assign array_update_78126[0] = add_78099 == 32'h0000_0000 ? add_78124 : array_index_78118[0];
  assign array_update_78126[1] = add_78099 == 32'h0000_0001 ? add_78124 : array_index_78118[1];
  assign array_update_78126[2] = add_78099 == 32'h0000_0002 ? add_78124 : array_index_78118[2];
  assign array_update_78126[3] = add_78099 == 32'h0000_0003 ? add_78124 : array_index_78118[3];
  assign array_update_78126[4] = add_78099 == 32'h0000_0004 ? add_78124 : array_index_78118[4];
  assign array_update_78126[5] = add_78099 == 32'h0000_0005 ? add_78124 : array_index_78118[5];
  assign array_update_78126[6] = add_78099 == 32'h0000_0006 ? add_78124 : array_index_78118[6];
  assign array_update_78126[7] = add_78099 == 32'h0000_0007 ? add_78124 : array_index_78118[7];
  assign array_update_78126[8] = add_78099 == 32'h0000_0008 ? add_78124 : array_index_78118[8];
  assign array_update_78126[9] = add_78099 == 32'h0000_0009 ? add_78124 : array_index_78118[9];
  assign add_78127 = add_78114 + 32'h0000_0001;
  assign array_update_78128[0] = add_77421 == 32'h0000_0000 ? array_update_78126 : array_update_78115[0];
  assign array_update_78128[1] = add_77421 == 32'h0000_0001 ? array_update_78126 : array_update_78115[1];
  assign array_update_78128[2] = add_77421 == 32'h0000_0002 ? array_update_78126 : array_update_78115[2];
  assign array_update_78128[3] = add_77421 == 32'h0000_0003 ? array_update_78126 : array_update_78115[3];
  assign array_update_78128[4] = add_77421 == 32'h0000_0004 ? array_update_78126 : array_update_78115[4];
  assign array_update_78128[5] = add_77421 == 32'h0000_0005 ? array_update_78126 : array_update_78115[5];
  assign array_update_78128[6] = add_77421 == 32'h0000_0006 ? array_update_78126 : array_update_78115[6];
  assign array_update_78128[7] = add_77421 == 32'h0000_0007 ? array_update_78126 : array_update_78115[7];
  assign array_update_78128[8] = add_77421 == 32'h0000_0008 ? array_update_78126 : array_update_78115[8];
  assign array_update_78128[9] = add_77421 == 32'h0000_0009 ? array_update_78126 : array_update_78115[9];
  assign array_index_78130 = array_update_72021[add_78127 > 32'h0000_0009 ? 4'h9 : add_78127[3:0]];
  assign array_index_78131 = array_update_78128[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_78135 = smul32b_32b_x_32b(array_index_77428[add_78127 > 32'h0000_0009 ? 4'h9 : add_78127[3:0]], array_index_78130[add_78099 > 32'h0000_0009 ? 4'h9 : add_78099[3:0]]);
  assign add_78137 = array_index_78131[add_78099 > 32'h0000_0009 ? 4'h9 : add_78099[3:0]] + smul_78135;
  assign array_update_78139[0] = add_78099 == 32'h0000_0000 ? add_78137 : array_index_78131[0];
  assign array_update_78139[1] = add_78099 == 32'h0000_0001 ? add_78137 : array_index_78131[1];
  assign array_update_78139[2] = add_78099 == 32'h0000_0002 ? add_78137 : array_index_78131[2];
  assign array_update_78139[3] = add_78099 == 32'h0000_0003 ? add_78137 : array_index_78131[3];
  assign array_update_78139[4] = add_78099 == 32'h0000_0004 ? add_78137 : array_index_78131[4];
  assign array_update_78139[5] = add_78099 == 32'h0000_0005 ? add_78137 : array_index_78131[5];
  assign array_update_78139[6] = add_78099 == 32'h0000_0006 ? add_78137 : array_index_78131[6];
  assign array_update_78139[7] = add_78099 == 32'h0000_0007 ? add_78137 : array_index_78131[7];
  assign array_update_78139[8] = add_78099 == 32'h0000_0008 ? add_78137 : array_index_78131[8];
  assign array_update_78139[9] = add_78099 == 32'h0000_0009 ? add_78137 : array_index_78131[9];
  assign add_78140 = add_78127 + 32'h0000_0001;
  assign array_update_78141[0] = add_77421 == 32'h0000_0000 ? array_update_78139 : array_update_78128[0];
  assign array_update_78141[1] = add_77421 == 32'h0000_0001 ? array_update_78139 : array_update_78128[1];
  assign array_update_78141[2] = add_77421 == 32'h0000_0002 ? array_update_78139 : array_update_78128[2];
  assign array_update_78141[3] = add_77421 == 32'h0000_0003 ? array_update_78139 : array_update_78128[3];
  assign array_update_78141[4] = add_77421 == 32'h0000_0004 ? array_update_78139 : array_update_78128[4];
  assign array_update_78141[5] = add_77421 == 32'h0000_0005 ? array_update_78139 : array_update_78128[5];
  assign array_update_78141[6] = add_77421 == 32'h0000_0006 ? array_update_78139 : array_update_78128[6];
  assign array_update_78141[7] = add_77421 == 32'h0000_0007 ? array_update_78139 : array_update_78128[7];
  assign array_update_78141[8] = add_77421 == 32'h0000_0008 ? array_update_78139 : array_update_78128[8];
  assign array_update_78141[9] = add_77421 == 32'h0000_0009 ? array_update_78139 : array_update_78128[9];
  assign array_index_78143 = array_update_72021[add_78140 > 32'h0000_0009 ? 4'h9 : add_78140[3:0]];
  assign array_index_78144 = array_update_78141[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_78148 = smul32b_32b_x_32b(array_index_77428[add_78140 > 32'h0000_0009 ? 4'h9 : add_78140[3:0]], array_index_78143[add_78099 > 32'h0000_0009 ? 4'h9 : add_78099[3:0]]);
  assign add_78150 = array_index_78144[add_78099 > 32'h0000_0009 ? 4'h9 : add_78099[3:0]] + smul_78148;
  assign array_update_78152[0] = add_78099 == 32'h0000_0000 ? add_78150 : array_index_78144[0];
  assign array_update_78152[1] = add_78099 == 32'h0000_0001 ? add_78150 : array_index_78144[1];
  assign array_update_78152[2] = add_78099 == 32'h0000_0002 ? add_78150 : array_index_78144[2];
  assign array_update_78152[3] = add_78099 == 32'h0000_0003 ? add_78150 : array_index_78144[3];
  assign array_update_78152[4] = add_78099 == 32'h0000_0004 ? add_78150 : array_index_78144[4];
  assign array_update_78152[5] = add_78099 == 32'h0000_0005 ? add_78150 : array_index_78144[5];
  assign array_update_78152[6] = add_78099 == 32'h0000_0006 ? add_78150 : array_index_78144[6];
  assign array_update_78152[7] = add_78099 == 32'h0000_0007 ? add_78150 : array_index_78144[7];
  assign array_update_78152[8] = add_78099 == 32'h0000_0008 ? add_78150 : array_index_78144[8];
  assign array_update_78152[9] = add_78099 == 32'h0000_0009 ? add_78150 : array_index_78144[9];
  assign add_78153 = add_78140 + 32'h0000_0001;
  assign array_update_78154[0] = add_77421 == 32'h0000_0000 ? array_update_78152 : array_update_78141[0];
  assign array_update_78154[1] = add_77421 == 32'h0000_0001 ? array_update_78152 : array_update_78141[1];
  assign array_update_78154[2] = add_77421 == 32'h0000_0002 ? array_update_78152 : array_update_78141[2];
  assign array_update_78154[3] = add_77421 == 32'h0000_0003 ? array_update_78152 : array_update_78141[3];
  assign array_update_78154[4] = add_77421 == 32'h0000_0004 ? array_update_78152 : array_update_78141[4];
  assign array_update_78154[5] = add_77421 == 32'h0000_0005 ? array_update_78152 : array_update_78141[5];
  assign array_update_78154[6] = add_77421 == 32'h0000_0006 ? array_update_78152 : array_update_78141[6];
  assign array_update_78154[7] = add_77421 == 32'h0000_0007 ? array_update_78152 : array_update_78141[7];
  assign array_update_78154[8] = add_77421 == 32'h0000_0008 ? array_update_78152 : array_update_78141[8];
  assign array_update_78154[9] = add_77421 == 32'h0000_0009 ? array_update_78152 : array_update_78141[9];
  assign array_index_78156 = array_update_72021[add_78153 > 32'h0000_0009 ? 4'h9 : add_78153[3:0]];
  assign array_index_78157 = array_update_78154[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_78161 = smul32b_32b_x_32b(array_index_77428[add_78153 > 32'h0000_0009 ? 4'h9 : add_78153[3:0]], array_index_78156[add_78099 > 32'h0000_0009 ? 4'h9 : add_78099[3:0]]);
  assign add_78163 = array_index_78157[add_78099 > 32'h0000_0009 ? 4'h9 : add_78099[3:0]] + smul_78161;
  assign array_update_78165[0] = add_78099 == 32'h0000_0000 ? add_78163 : array_index_78157[0];
  assign array_update_78165[1] = add_78099 == 32'h0000_0001 ? add_78163 : array_index_78157[1];
  assign array_update_78165[2] = add_78099 == 32'h0000_0002 ? add_78163 : array_index_78157[2];
  assign array_update_78165[3] = add_78099 == 32'h0000_0003 ? add_78163 : array_index_78157[3];
  assign array_update_78165[4] = add_78099 == 32'h0000_0004 ? add_78163 : array_index_78157[4];
  assign array_update_78165[5] = add_78099 == 32'h0000_0005 ? add_78163 : array_index_78157[5];
  assign array_update_78165[6] = add_78099 == 32'h0000_0006 ? add_78163 : array_index_78157[6];
  assign array_update_78165[7] = add_78099 == 32'h0000_0007 ? add_78163 : array_index_78157[7];
  assign array_update_78165[8] = add_78099 == 32'h0000_0008 ? add_78163 : array_index_78157[8];
  assign array_update_78165[9] = add_78099 == 32'h0000_0009 ? add_78163 : array_index_78157[9];
  assign add_78166 = add_78153 + 32'h0000_0001;
  assign array_update_78167[0] = add_77421 == 32'h0000_0000 ? array_update_78165 : array_update_78154[0];
  assign array_update_78167[1] = add_77421 == 32'h0000_0001 ? array_update_78165 : array_update_78154[1];
  assign array_update_78167[2] = add_77421 == 32'h0000_0002 ? array_update_78165 : array_update_78154[2];
  assign array_update_78167[3] = add_77421 == 32'h0000_0003 ? array_update_78165 : array_update_78154[3];
  assign array_update_78167[4] = add_77421 == 32'h0000_0004 ? array_update_78165 : array_update_78154[4];
  assign array_update_78167[5] = add_77421 == 32'h0000_0005 ? array_update_78165 : array_update_78154[5];
  assign array_update_78167[6] = add_77421 == 32'h0000_0006 ? array_update_78165 : array_update_78154[6];
  assign array_update_78167[7] = add_77421 == 32'h0000_0007 ? array_update_78165 : array_update_78154[7];
  assign array_update_78167[8] = add_77421 == 32'h0000_0008 ? array_update_78165 : array_update_78154[8];
  assign array_update_78167[9] = add_77421 == 32'h0000_0009 ? array_update_78165 : array_update_78154[9];
  assign array_index_78169 = array_update_72021[add_78166 > 32'h0000_0009 ? 4'h9 : add_78166[3:0]];
  assign array_index_78170 = array_update_78167[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_78174 = smul32b_32b_x_32b(array_index_77428[add_78166 > 32'h0000_0009 ? 4'h9 : add_78166[3:0]], array_index_78169[add_78099 > 32'h0000_0009 ? 4'h9 : add_78099[3:0]]);
  assign add_78176 = array_index_78170[add_78099 > 32'h0000_0009 ? 4'h9 : add_78099[3:0]] + smul_78174;
  assign array_update_78178[0] = add_78099 == 32'h0000_0000 ? add_78176 : array_index_78170[0];
  assign array_update_78178[1] = add_78099 == 32'h0000_0001 ? add_78176 : array_index_78170[1];
  assign array_update_78178[2] = add_78099 == 32'h0000_0002 ? add_78176 : array_index_78170[2];
  assign array_update_78178[3] = add_78099 == 32'h0000_0003 ? add_78176 : array_index_78170[3];
  assign array_update_78178[4] = add_78099 == 32'h0000_0004 ? add_78176 : array_index_78170[4];
  assign array_update_78178[5] = add_78099 == 32'h0000_0005 ? add_78176 : array_index_78170[5];
  assign array_update_78178[6] = add_78099 == 32'h0000_0006 ? add_78176 : array_index_78170[6];
  assign array_update_78178[7] = add_78099 == 32'h0000_0007 ? add_78176 : array_index_78170[7];
  assign array_update_78178[8] = add_78099 == 32'h0000_0008 ? add_78176 : array_index_78170[8];
  assign array_update_78178[9] = add_78099 == 32'h0000_0009 ? add_78176 : array_index_78170[9];
  assign add_78179 = add_78166 + 32'h0000_0001;
  assign array_update_78180[0] = add_77421 == 32'h0000_0000 ? array_update_78178 : array_update_78167[0];
  assign array_update_78180[1] = add_77421 == 32'h0000_0001 ? array_update_78178 : array_update_78167[1];
  assign array_update_78180[2] = add_77421 == 32'h0000_0002 ? array_update_78178 : array_update_78167[2];
  assign array_update_78180[3] = add_77421 == 32'h0000_0003 ? array_update_78178 : array_update_78167[3];
  assign array_update_78180[4] = add_77421 == 32'h0000_0004 ? array_update_78178 : array_update_78167[4];
  assign array_update_78180[5] = add_77421 == 32'h0000_0005 ? array_update_78178 : array_update_78167[5];
  assign array_update_78180[6] = add_77421 == 32'h0000_0006 ? array_update_78178 : array_update_78167[6];
  assign array_update_78180[7] = add_77421 == 32'h0000_0007 ? array_update_78178 : array_update_78167[7];
  assign array_update_78180[8] = add_77421 == 32'h0000_0008 ? array_update_78178 : array_update_78167[8];
  assign array_update_78180[9] = add_77421 == 32'h0000_0009 ? array_update_78178 : array_update_78167[9];
  assign array_index_78182 = array_update_72021[add_78179 > 32'h0000_0009 ? 4'h9 : add_78179[3:0]];
  assign array_index_78183 = array_update_78180[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_78187 = smul32b_32b_x_32b(array_index_77428[add_78179 > 32'h0000_0009 ? 4'h9 : add_78179[3:0]], array_index_78182[add_78099 > 32'h0000_0009 ? 4'h9 : add_78099[3:0]]);
  assign add_78189 = array_index_78183[add_78099 > 32'h0000_0009 ? 4'h9 : add_78099[3:0]] + smul_78187;
  assign array_update_78191[0] = add_78099 == 32'h0000_0000 ? add_78189 : array_index_78183[0];
  assign array_update_78191[1] = add_78099 == 32'h0000_0001 ? add_78189 : array_index_78183[1];
  assign array_update_78191[2] = add_78099 == 32'h0000_0002 ? add_78189 : array_index_78183[2];
  assign array_update_78191[3] = add_78099 == 32'h0000_0003 ? add_78189 : array_index_78183[3];
  assign array_update_78191[4] = add_78099 == 32'h0000_0004 ? add_78189 : array_index_78183[4];
  assign array_update_78191[5] = add_78099 == 32'h0000_0005 ? add_78189 : array_index_78183[5];
  assign array_update_78191[6] = add_78099 == 32'h0000_0006 ? add_78189 : array_index_78183[6];
  assign array_update_78191[7] = add_78099 == 32'h0000_0007 ? add_78189 : array_index_78183[7];
  assign array_update_78191[8] = add_78099 == 32'h0000_0008 ? add_78189 : array_index_78183[8];
  assign array_update_78191[9] = add_78099 == 32'h0000_0009 ? add_78189 : array_index_78183[9];
  assign add_78192 = add_78179 + 32'h0000_0001;
  assign array_update_78193[0] = add_77421 == 32'h0000_0000 ? array_update_78191 : array_update_78180[0];
  assign array_update_78193[1] = add_77421 == 32'h0000_0001 ? array_update_78191 : array_update_78180[1];
  assign array_update_78193[2] = add_77421 == 32'h0000_0002 ? array_update_78191 : array_update_78180[2];
  assign array_update_78193[3] = add_77421 == 32'h0000_0003 ? array_update_78191 : array_update_78180[3];
  assign array_update_78193[4] = add_77421 == 32'h0000_0004 ? array_update_78191 : array_update_78180[4];
  assign array_update_78193[5] = add_77421 == 32'h0000_0005 ? array_update_78191 : array_update_78180[5];
  assign array_update_78193[6] = add_77421 == 32'h0000_0006 ? array_update_78191 : array_update_78180[6];
  assign array_update_78193[7] = add_77421 == 32'h0000_0007 ? array_update_78191 : array_update_78180[7];
  assign array_update_78193[8] = add_77421 == 32'h0000_0008 ? array_update_78191 : array_update_78180[8];
  assign array_update_78193[9] = add_77421 == 32'h0000_0009 ? array_update_78191 : array_update_78180[9];
  assign array_index_78195 = array_update_72021[add_78192 > 32'h0000_0009 ? 4'h9 : add_78192[3:0]];
  assign array_index_78196 = array_update_78193[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_78200 = smul32b_32b_x_32b(array_index_77428[add_78192 > 32'h0000_0009 ? 4'h9 : add_78192[3:0]], array_index_78195[add_78099 > 32'h0000_0009 ? 4'h9 : add_78099[3:0]]);
  assign add_78202 = array_index_78196[add_78099 > 32'h0000_0009 ? 4'h9 : add_78099[3:0]] + smul_78200;
  assign array_update_78204[0] = add_78099 == 32'h0000_0000 ? add_78202 : array_index_78196[0];
  assign array_update_78204[1] = add_78099 == 32'h0000_0001 ? add_78202 : array_index_78196[1];
  assign array_update_78204[2] = add_78099 == 32'h0000_0002 ? add_78202 : array_index_78196[2];
  assign array_update_78204[3] = add_78099 == 32'h0000_0003 ? add_78202 : array_index_78196[3];
  assign array_update_78204[4] = add_78099 == 32'h0000_0004 ? add_78202 : array_index_78196[4];
  assign array_update_78204[5] = add_78099 == 32'h0000_0005 ? add_78202 : array_index_78196[5];
  assign array_update_78204[6] = add_78099 == 32'h0000_0006 ? add_78202 : array_index_78196[6];
  assign array_update_78204[7] = add_78099 == 32'h0000_0007 ? add_78202 : array_index_78196[7];
  assign array_update_78204[8] = add_78099 == 32'h0000_0008 ? add_78202 : array_index_78196[8];
  assign array_update_78204[9] = add_78099 == 32'h0000_0009 ? add_78202 : array_index_78196[9];
  assign add_78205 = add_78192 + 32'h0000_0001;
  assign array_update_78206[0] = add_77421 == 32'h0000_0000 ? array_update_78204 : array_update_78193[0];
  assign array_update_78206[1] = add_77421 == 32'h0000_0001 ? array_update_78204 : array_update_78193[1];
  assign array_update_78206[2] = add_77421 == 32'h0000_0002 ? array_update_78204 : array_update_78193[2];
  assign array_update_78206[3] = add_77421 == 32'h0000_0003 ? array_update_78204 : array_update_78193[3];
  assign array_update_78206[4] = add_77421 == 32'h0000_0004 ? array_update_78204 : array_update_78193[4];
  assign array_update_78206[5] = add_77421 == 32'h0000_0005 ? array_update_78204 : array_update_78193[5];
  assign array_update_78206[6] = add_77421 == 32'h0000_0006 ? array_update_78204 : array_update_78193[6];
  assign array_update_78206[7] = add_77421 == 32'h0000_0007 ? array_update_78204 : array_update_78193[7];
  assign array_update_78206[8] = add_77421 == 32'h0000_0008 ? array_update_78204 : array_update_78193[8];
  assign array_update_78206[9] = add_77421 == 32'h0000_0009 ? array_update_78204 : array_update_78193[9];
  assign array_index_78208 = array_update_72021[add_78205 > 32'h0000_0009 ? 4'h9 : add_78205[3:0]];
  assign array_index_78209 = array_update_78206[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_78213 = smul32b_32b_x_32b(array_index_77428[add_78205 > 32'h0000_0009 ? 4'h9 : add_78205[3:0]], array_index_78208[add_78099 > 32'h0000_0009 ? 4'h9 : add_78099[3:0]]);
  assign add_78215 = array_index_78209[add_78099 > 32'h0000_0009 ? 4'h9 : add_78099[3:0]] + smul_78213;
  assign array_update_78217[0] = add_78099 == 32'h0000_0000 ? add_78215 : array_index_78209[0];
  assign array_update_78217[1] = add_78099 == 32'h0000_0001 ? add_78215 : array_index_78209[1];
  assign array_update_78217[2] = add_78099 == 32'h0000_0002 ? add_78215 : array_index_78209[2];
  assign array_update_78217[3] = add_78099 == 32'h0000_0003 ? add_78215 : array_index_78209[3];
  assign array_update_78217[4] = add_78099 == 32'h0000_0004 ? add_78215 : array_index_78209[4];
  assign array_update_78217[5] = add_78099 == 32'h0000_0005 ? add_78215 : array_index_78209[5];
  assign array_update_78217[6] = add_78099 == 32'h0000_0006 ? add_78215 : array_index_78209[6];
  assign array_update_78217[7] = add_78099 == 32'h0000_0007 ? add_78215 : array_index_78209[7];
  assign array_update_78217[8] = add_78099 == 32'h0000_0008 ? add_78215 : array_index_78209[8];
  assign array_update_78217[9] = add_78099 == 32'h0000_0009 ? add_78215 : array_index_78209[9];
  assign add_78218 = add_78205 + 32'h0000_0001;
  assign array_update_78219[0] = add_77421 == 32'h0000_0000 ? array_update_78217 : array_update_78206[0];
  assign array_update_78219[1] = add_77421 == 32'h0000_0001 ? array_update_78217 : array_update_78206[1];
  assign array_update_78219[2] = add_77421 == 32'h0000_0002 ? array_update_78217 : array_update_78206[2];
  assign array_update_78219[3] = add_77421 == 32'h0000_0003 ? array_update_78217 : array_update_78206[3];
  assign array_update_78219[4] = add_77421 == 32'h0000_0004 ? array_update_78217 : array_update_78206[4];
  assign array_update_78219[5] = add_77421 == 32'h0000_0005 ? array_update_78217 : array_update_78206[5];
  assign array_update_78219[6] = add_77421 == 32'h0000_0006 ? array_update_78217 : array_update_78206[6];
  assign array_update_78219[7] = add_77421 == 32'h0000_0007 ? array_update_78217 : array_update_78206[7];
  assign array_update_78219[8] = add_77421 == 32'h0000_0008 ? array_update_78217 : array_update_78206[8];
  assign array_update_78219[9] = add_77421 == 32'h0000_0009 ? array_update_78217 : array_update_78206[9];
  assign array_index_78221 = array_update_72021[add_78218 > 32'h0000_0009 ? 4'h9 : add_78218[3:0]];
  assign array_index_78222 = array_update_78219[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_78226 = smul32b_32b_x_32b(array_index_77428[add_78218 > 32'h0000_0009 ? 4'h9 : add_78218[3:0]], array_index_78221[add_78099 > 32'h0000_0009 ? 4'h9 : add_78099[3:0]]);
  assign add_78228 = array_index_78222[add_78099 > 32'h0000_0009 ? 4'h9 : add_78099[3:0]] + smul_78226;
  assign array_update_78229[0] = add_78099 == 32'h0000_0000 ? add_78228 : array_index_78222[0];
  assign array_update_78229[1] = add_78099 == 32'h0000_0001 ? add_78228 : array_index_78222[1];
  assign array_update_78229[2] = add_78099 == 32'h0000_0002 ? add_78228 : array_index_78222[2];
  assign array_update_78229[3] = add_78099 == 32'h0000_0003 ? add_78228 : array_index_78222[3];
  assign array_update_78229[4] = add_78099 == 32'h0000_0004 ? add_78228 : array_index_78222[4];
  assign array_update_78229[5] = add_78099 == 32'h0000_0005 ? add_78228 : array_index_78222[5];
  assign array_update_78229[6] = add_78099 == 32'h0000_0006 ? add_78228 : array_index_78222[6];
  assign array_update_78229[7] = add_78099 == 32'h0000_0007 ? add_78228 : array_index_78222[7];
  assign array_update_78229[8] = add_78099 == 32'h0000_0008 ? add_78228 : array_index_78222[8];
  assign array_update_78229[9] = add_78099 == 32'h0000_0009 ? add_78228 : array_index_78222[9];
  assign array_update_78230[0] = add_77421 == 32'h0000_0000 ? array_update_78229 : array_update_78219[0];
  assign array_update_78230[1] = add_77421 == 32'h0000_0001 ? array_update_78229 : array_update_78219[1];
  assign array_update_78230[2] = add_77421 == 32'h0000_0002 ? array_update_78229 : array_update_78219[2];
  assign array_update_78230[3] = add_77421 == 32'h0000_0003 ? array_update_78229 : array_update_78219[3];
  assign array_update_78230[4] = add_77421 == 32'h0000_0004 ? array_update_78229 : array_update_78219[4];
  assign array_update_78230[5] = add_77421 == 32'h0000_0005 ? array_update_78229 : array_update_78219[5];
  assign array_update_78230[6] = add_77421 == 32'h0000_0006 ? array_update_78229 : array_update_78219[6];
  assign array_update_78230[7] = add_77421 == 32'h0000_0007 ? array_update_78229 : array_update_78219[7];
  assign array_update_78230[8] = add_77421 == 32'h0000_0008 ? array_update_78229 : array_update_78219[8];
  assign array_update_78230[9] = add_77421 == 32'h0000_0009 ? array_update_78229 : array_update_78219[9];
  assign array_index_78232 = array_update_78230[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign add_78234 = add_78099 + 32'h0000_0001;
  assign array_update_78235[0] = add_78234 == 32'h0000_0000 ? 32'h0000_0000 : array_index_78232[0];
  assign array_update_78235[1] = add_78234 == 32'h0000_0001 ? 32'h0000_0000 : array_index_78232[1];
  assign array_update_78235[2] = add_78234 == 32'h0000_0002 ? 32'h0000_0000 : array_index_78232[2];
  assign array_update_78235[3] = add_78234 == 32'h0000_0003 ? 32'h0000_0000 : array_index_78232[3];
  assign array_update_78235[4] = add_78234 == 32'h0000_0004 ? 32'h0000_0000 : array_index_78232[4];
  assign array_update_78235[5] = add_78234 == 32'h0000_0005 ? 32'h0000_0000 : array_index_78232[5];
  assign array_update_78235[6] = add_78234 == 32'h0000_0006 ? 32'h0000_0000 : array_index_78232[6];
  assign array_update_78235[7] = add_78234 == 32'h0000_0007 ? 32'h0000_0000 : array_index_78232[7];
  assign array_update_78235[8] = add_78234 == 32'h0000_0008 ? 32'h0000_0000 : array_index_78232[8];
  assign array_update_78235[9] = add_78234 == 32'h0000_0009 ? 32'h0000_0000 : array_index_78232[9];
  assign literal_78236 = 32'h0000_0000;
  assign array_update_78237[0] = add_77421 == 32'h0000_0000 ? array_update_78235 : array_update_78230[0];
  assign array_update_78237[1] = add_77421 == 32'h0000_0001 ? array_update_78235 : array_update_78230[1];
  assign array_update_78237[2] = add_77421 == 32'h0000_0002 ? array_update_78235 : array_update_78230[2];
  assign array_update_78237[3] = add_77421 == 32'h0000_0003 ? array_update_78235 : array_update_78230[3];
  assign array_update_78237[4] = add_77421 == 32'h0000_0004 ? array_update_78235 : array_update_78230[4];
  assign array_update_78237[5] = add_77421 == 32'h0000_0005 ? array_update_78235 : array_update_78230[5];
  assign array_update_78237[6] = add_77421 == 32'h0000_0006 ? array_update_78235 : array_update_78230[6];
  assign array_update_78237[7] = add_77421 == 32'h0000_0007 ? array_update_78235 : array_update_78230[7];
  assign array_update_78237[8] = add_77421 == 32'h0000_0008 ? array_update_78235 : array_update_78230[8];
  assign array_update_78237[9] = add_77421 == 32'h0000_0009 ? array_update_78235 : array_update_78230[9];
  assign array_index_78239 = array_update_72021[literal_78236 > 32'h0000_0009 ? 4'h9 : literal_78236[3:0]];
  assign array_index_78240 = array_update_78237[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_78244 = smul32b_32b_x_32b(array_index_77428[literal_78236 > 32'h0000_0009 ? 4'h9 : literal_78236[3:0]], array_index_78239[add_78234 > 32'h0000_0009 ? 4'h9 : add_78234[3:0]]);
  assign add_78246 = array_index_78240[add_78234 > 32'h0000_0009 ? 4'h9 : add_78234[3:0]] + smul_78244;
  assign array_update_78248[0] = add_78234 == 32'h0000_0000 ? add_78246 : array_index_78240[0];
  assign array_update_78248[1] = add_78234 == 32'h0000_0001 ? add_78246 : array_index_78240[1];
  assign array_update_78248[2] = add_78234 == 32'h0000_0002 ? add_78246 : array_index_78240[2];
  assign array_update_78248[3] = add_78234 == 32'h0000_0003 ? add_78246 : array_index_78240[3];
  assign array_update_78248[4] = add_78234 == 32'h0000_0004 ? add_78246 : array_index_78240[4];
  assign array_update_78248[5] = add_78234 == 32'h0000_0005 ? add_78246 : array_index_78240[5];
  assign array_update_78248[6] = add_78234 == 32'h0000_0006 ? add_78246 : array_index_78240[6];
  assign array_update_78248[7] = add_78234 == 32'h0000_0007 ? add_78246 : array_index_78240[7];
  assign array_update_78248[8] = add_78234 == 32'h0000_0008 ? add_78246 : array_index_78240[8];
  assign array_update_78248[9] = add_78234 == 32'h0000_0009 ? add_78246 : array_index_78240[9];
  assign add_78249 = literal_78236 + 32'h0000_0001;
  assign array_update_78250[0] = add_77421 == 32'h0000_0000 ? array_update_78248 : array_update_78237[0];
  assign array_update_78250[1] = add_77421 == 32'h0000_0001 ? array_update_78248 : array_update_78237[1];
  assign array_update_78250[2] = add_77421 == 32'h0000_0002 ? array_update_78248 : array_update_78237[2];
  assign array_update_78250[3] = add_77421 == 32'h0000_0003 ? array_update_78248 : array_update_78237[3];
  assign array_update_78250[4] = add_77421 == 32'h0000_0004 ? array_update_78248 : array_update_78237[4];
  assign array_update_78250[5] = add_77421 == 32'h0000_0005 ? array_update_78248 : array_update_78237[5];
  assign array_update_78250[6] = add_77421 == 32'h0000_0006 ? array_update_78248 : array_update_78237[6];
  assign array_update_78250[7] = add_77421 == 32'h0000_0007 ? array_update_78248 : array_update_78237[7];
  assign array_update_78250[8] = add_77421 == 32'h0000_0008 ? array_update_78248 : array_update_78237[8];
  assign array_update_78250[9] = add_77421 == 32'h0000_0009 ? array_update_78248 : array_update_78237[9];
  assign array_index_78252 = array_update_72021[add_78249 > 32'h0000_0009 ? 4'h9 : add_78249[3:0]];
  assign array_index_78253 = array_update_78250[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_78257 = smul32b_32b_x_32b(array_index_77428[add_78249 > 32'h0000_0009 ? 4'h9 : add_78249[3:0]], array_index_78252[add_78234 > 32'h0000_0009 ? 4'h9 : add_78234[3:0]]);
  assign add_78259 = array_index_78253[add_78234 > 32'h0000_0009 ? 4'h9 : add_78234[3:0]] + smul_78257;
  assign array_update_78261[0] = add_78234 == 32'h0000_0000 ? add_78259 : array_index_78253[0];
  assign array_update_78261[1] = add_78234 == 32'h0000_0001 ? add_78259 : array_index_78253[1];
  assign array_update_78261[2] = add_78234 == 32'h0000_0002 ? add_78259 : array_index_78253[2];
  assign array_update_78261[3] = add_78234 == 32'h0000_0003 ? add_78259 : array_index_78253[3];
  assign array_update_78261[4] = add_78234 == 32'h0000_0004 ? add_78259 : array_index_78253[4];
  assign array_update_78261[5] = add_78234 == 32'h0000_0005 ? add_78259 : array_index_78253[5];
  assign array_update_78261[6] = add_78234 == 32'h0000_0006 ? add_78259 : array_index_78253[6];
  assign array_update_78261[7] = add_78234 == 32'h0000_0007 ? add_78259 : array_index_78253[7];
  assign array_update_78261[8] = add_78234 == 32'h0000_0008 ? add_78259 : array_index_78253[8];
  assign array_update_78261[9] = add_78234 == 32'h0000_0009 ? add_78259 : array_index_78253[9];
  assign add_78262 = add_78249 + 32'h0000_0001;
  assign array_update_78263[0] = add_77421 == 32'h0000_0000 ? array_update_78261 : array_update_78250[0];
  assign array_update_78263[1] = add_77421 == 32'h0000_0001 ? array_update_78261 : array_update_78250[1];
  assign array_update_78263[2] = add_77421 == 32'h0000_0002 ? array_update_78261 : array_update_78250[2];
  assign array_update_78263[3] = add_77421 == 32'h0000_0003 ? array_update_78261 : array_update_78250[3];
  assign array_update_78263[4] = add_77421 == 32'h0000_0004 ? array_update_78261 : array_update_78250[4];
  assign array_update_78263[5] = add_77421 == 32'h0000_0005 ? array_update_78261 : array_update_78250[5];
  assign array_update_78263[6] = add_77421 == 32'h0000_0006 ? array_update_78261 : array_update_78250[6];
  assign array_update_78263[7] = add_77421 == 32'h0000_0007 ? array_update_78261 : array_update_78250[7];
  assign array_update_78263[8] = add_77421 == 32'h0000_0008 ? array_update_78261 : array_update_78250[8];
  assign array_update_78263[9] = add_77421 == 32'h0000_0009 ? array_update_78261 : array_update_78250[9];
  assign array_index_78265 = array_update_72021[add_78262 > 32'h0000_0009 ? 4'h9 : add_78262[3:0]];
  assign array_index_78266 = array_update_78263[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_78270 = smul32b_32b_x_32b(array_index_77428[add_78262 > 32'h0000_0009 ? 4'h9 : add_78262[3:0]], array_index_78265[add_78234 > 32'h0000_0009 ? 4'h9 : add_78234[3:0]]);
  assign add_78272 = array_index_78266[add_78234 > 32'h0000_0009 ? 4'h9 : add_78234[3:0]] + smul_78270;
  assign array_update_78274[0] = add_78234 == 32'h0000_0000 ? add_78272 : array_index_78266[0];
  assign array_update_78274[1] = add_78234 == 32'h0000_0001 ? add_78272 : array_index_78266[1];
  assign array_update_78274[2] = add_78234 == 32'h0000_0002 ? add_78272 : array_index_78266[2];
  assign array_update_78274[3] = add_78234 == 32'h0000_0003 ? add_78272 : array_index_78266[3];
  assign array_update_78274[4] = add_78234 == 32'h0000_0004 ? add_78272 : array_index_78266[4];
  assign array_update_78274[5] = add_78234 == 32'h0000_0005 ? add_78272 : array_index_78266[5];
  assign array_update_78274[6] = add_78234 == 32'h0000_0006 ? add_78272 : array_index_78266[6];
  assign array_update_78274[7] = add_78234 == 32'h0000_0007 ? add_78272 : array_index_78266[7];
  assign array_update_78274[8] = add_78234 == 32'h0000_0008 ? add_78272 : array_index_78266[8];
  assign array_update_78274[9] = add_78234 == 32'h0000_0009 ? add_78272 : array_index_78266[9];
  assign add_78275 = add_78262 + 32'h0000_0001;
  assign array_update_78276[0] = add_77421 == 32'h0000_0000 ? array_update_78274 : array_update_78263[0];
  assign array_update_78276[1] = add_77421 == 32'h0000_0001 ? array_update_78274 : array_update_78263[1];
  assign array_update_78276[2] = add_77421 == 32'h0000_0002 ? array_update_78274 : array_update_78263[2];
  assign array_update_78276[3] = add_77421 == 32'h0000_0003 ? array_update_78274 : array_update_78263[3];
  assign array_update_78276[4] = add_77421 == 32'h0000_0004 ? array_update_78274 : array_update_78263[4];
  assign array_update_78276[5] = add_77421 == 32'h0000_0005 ? array_update_78274 : array_update_78263[5];
  assign array_update_78276[6] = add_77421 == 32'h0000_0006 ? array_update_78274 : array_update_78263[6];
  assign array_update_78276[7] = add_77421 == 32'h0000_0007 ? array_update_78274 : array_update_78263[7];
  assign array_update_78276[8] = add_77421 == 32'h0000_0008 ? array_update_78274 : array_update_78263[8];
  assign array_update_78276[9] = add_77421 == 32'h0000_0009 ? array_update_78274 : array_update_78263[9];
  assign array_index_78278 = array_update_72021[add_78275 > 32'h0000_0009 ? 4'h9 : add_78275[3:0]];
  assign array_index_78279 = array_update_78276[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_78283 = smul32b_32b_x_32b(array_index_77428[add_78275 > 32'h0000_0009 ? 4'h9 : add_78275[3:0]], array_index_78278[add_78234 > 32'h0000_0009 ? 4'h9 : add_78234[3:0]]);
  assign add_78285 = array_index_78279[add_78234 > 32'h0000_0009 ? 4'h9 : add_78234[3:0]] + smul_78283;
  assign array_update_78287[0] = add_78234 == 32'h0000_0000 ? add_78285 : array_index_78279[0];
  assign array_update_78287[1] = add_78234 == 32'h0000_0001 ? add_78285 : array_index_78279[1];
  assign array_update_78287[2] = add_78234 == 32'h0000_0002 ? add_78285 : array_index_78279[2];
  assign array_update_78287[3] = add_78234 == 32'h0000_0003 ? add_78285 : array_index_78279[3];
  assign array_update_78287[4] = add_78234 == 32'h0000_0004 ? add_78285 : array_index_78279[4];
  assign array_update_78287[5] = add_78234 == 32'h0000_0005 ? add_78285 : array_index_78279[5];
  assign array_update_78287[6] = add_78234 == 32'h0000_0006 ? add_78285 : array_index_78279[6];
  assign array_update_78287[7] = add_78234 == 32'h0000_0007 ? add_78285 : array_index_78279[7];
  assign array_update_78287[8] = add_78234 == 32'h0000_0008 ? add_78285 : array_index_78279[8];
  assign array_update_78287[9] = add_78234 == 32'h0000_0009 ? add_78285 : array_index_78279[9];
  assign add_78288 = add_78275 + 32'h0000_0001;
  assign array_update_78289[0] = add_77421 == 32'h0000_0000 ? array_update_78287 : array_update_78276[0];
  assign array_update_78289[1] = add_77421 == 32'h0000_0001 ? array_update_78287 : array_update_78276[1];
  assign array_update_78289[2] = add_77421 == 32'h0000_0002 ? array_update_78287 : array_update_78276[2];
  assign array_update_78289[3] = add_77421 == 32'h0000_0003 ? array_update_78287 : array_update_78276[3];
  assign array_update_78289[4] = add_77421 == 32'h0000_0004 ? array_update_78287 : array_update_78276[4];
  assign array_update_78289[5] = add_77421 == 32'h0000_0005 ? array_update_78287 : array_update_78276[5];
  assign array_update_78289[6] = add_77421 == 32'h0000_0006 ? array_update_78287 : array_update_78276[6];
  assign array_update_78289[7] = add_77421 == 32'h0000_0007 ? array_update_78287 : array_update_78276[7];
  assign array_update_78289[8] = add_77421 == 32'h0000_0008 ? array_update_78287 : array_update_78276[8];
  assign array_update_78289[9] = add_77421 == 32'h0000_0009 ? array_update_78287 : array_update_78276[9];
  assign array_index_78291 = array_update_72021[add_78288 > 32'h0000_0009 ? 4'h9 : add_78288[3:0]];
  assign array_index_78292 = array_update_78289[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_78296 = smul32b_32b_x_32b(array_index_77428[add_78288 > 32'h0000_0009 ? 4'h9 : add_78288[3:0]], array_index_78291[add_78234 > 32'h0000_0009 ? 4'h9 : add_78234[3:0]]);
  assign add_78298 = array_index_78292[add_78234 > 32'h0000_0009 ? 4'h9 : add_78234[3:0]] + smul_78296;
  assign array_update_78300[0] = add_78234 == 32'h0000_0000 ? add_78298 : array_index_78292[0];
  assign array_update_78300[1] = add_78234 == 32'h0000_0001 ? add_78298 : array_index_78292[1];
  assign array_update_78300[2] = add_78234 == 32'h0000_0002 ? add_78298 : array_index_78292[2];
  assign array_update_78300[3] = add_78234 == 32'h0000_0003 ? add_78298 : array_index_78292[3];
  assign array_update_78300[4] = add_78234 == 32'h0000_0004 ? add_78298 : array_index_78292[4];
  assign array_update_78300[5] = add_78234 == 32'h0000_0005 ? add_78298 : array_index_78292[5];
  assign array_update_78300[6] = add_78234 == 32'h0000_0006 ? add_78298 : array_index_78292[6];
  assign array_update_78300[7] = add_78234 == 32'h0000_0007 ? add_78298 : array_index_78292[7];
  assign array_update_78300[8] = add_78234 == 32'h0000_0008 ? add_78298 : array_index_78292[8];
  assign array_update_78300[9] = add_78234 == 32'h0000_0009 ? add_78298 : array_index_78292[9];
  assign add_78301 = add_78288 + 32'h0000_0001;
  assign array_update_78302[0] = add_77421 == 32'h0000_0000 ? array_update_78300 : array_update_78289[0];
  assign array_update_78302[1] = add_77421 == 32'h0000_0001 ? array_update_78300 : array_update_78289[1];
  assign array_update_78302[2] = add_77421 == 32'h0000_0002 ? array_update_78300 : array_update_78289[2];
  assign array_update_78302[3] = add_77421 == 32'h0000_0003 ? array_update_78300 : array_update_78289[3];
  assign array_update_78302[4] = add_77421 == 32'h0000_0004 ? array_update_78300 : array_update_78289[4];
  assign array_update_78302[5] = add_77421 == 32'h0000_0005 ? array_update_78300 : array_update_78289[5];
  assign array_update_78302[6] = add_77421 == 32'h0000_0006 ? array_update_78300 : array_update_78289[6];
  assign array_update_78302[7] = add_77421 == 32'h0000_0007 ? array_update_78300 : array_update_78289[7];
  assign array_update_78302[8] = add_77421 == 32'h0000_0008 ? array_update_78300 : array_update_78289[8];
  assign array_update_78302[9] = add_77421 == 32'h0000_0009 ? array_update_78300 : array_update_78289[9];
  assign array_index_78304 = array_update_72021[add_78301 > 32'h0000_0009 ? 4'h9 : add_78301[3:0]];
  assign array_index_78305 = array_update_78302[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_78309 = smul32b_32b_x_32b(array_index_77428[add_78301 > 32'h0000_0009 ? 4'h9 : add_78301[3:0]], array_index_78304[add_78234 > 32'h0000_0009 ? 4'h9 : add_78234[3:0]]);
  assign add_78311 = array_index_78305[add_78234 > 32'h0000_0009 ? 4'h9 : add_78234[3:0]] + smul_78309;
  assign array_update_78313[0] = add_78234 == 32'h0000_0000 ? add_78311 : array_index_78305[0];
  assign array_update_78313[1] = add_78234 == 32'h0000_0001 ? add_78311 : array_index_78305[1];
  assign array_update_78313[2] = add_78234 == 32'h0000_0002 ? add_78311 : array_index_78305[2];
  assign array_update_78313[3] = add_78234 == 32'h0000_0003 ? add_78311 : array_index_78305[3];
  assign array_update_78313[4] = add_78234 == 32'h0000_0004 ? add_78311 : array_index_78305[4];
  assign array_update_78313[5] = add_78234 == 32'h0000_0005 ? add_78311 : array_index_78305[5];
  assign array_update_78313[6] = add_78234 == 32'h0000_0006 ? add_78311 : array_index_78305[6];
  assign array_update_78313[7] = add_78234 == 32'h0000_0007 ? add_78311 : array_index_78305[7];
  assign array_update_78313[8] = add_78234 == 32'h0000_0008 ? add_78311 : array_index_78305[8];
  assign array_update_78313[9] = add_78234 == 32'h0000_0009 ? add_78311 : array_index_78305[9];
  assign add_78314 = add_78301 + 32'h0000_0001;
  assign array_update_78315[0] = add_77421 == 32'h0000_0000 ? array_update_78313 : array_update_78302[0];
  assign array_update_78315[1] = add_77421 == 32'h0000_0001 ? array_update_78313 : array_update_78302[1];
  assign array_update_78315[2] = add_77421 == 32'h0000_0002 ? array_update_78313 : array_update_78302[2];
  assign array_update_78315[3] = add_77421 == 32'h0000_0003 ? array_update_78313 : array_update_78302[3];
  assign array_update_78315[4] = add_77421 == 32'h0000_0004 ? array_update_78313 : array_update_78302[4];
  assign array_update_78315[5] = add_77421 == 32'h0000_0005 ? array_update_78313 : array_update_78302[5];
  assign array_update_78315[6] = add_77421 == 32'h0000_0006 ? array_update_78313 : array_update_78302[6];
  assign array_update_78315[7] = add_77421 == 32'h0000_0007 ? array_update_78313 : array_update_78302[7];
  assign array_update_78315[8] = add_77421 == 32'h0000_0008 ? array_update_78313 : array_update_78302[8];
  assign array_update_78315[9] = add_77421 == 32'h0000_0009 ? array_update_78313 : array_update_78302[9];
  assign array_index_78317 = array_update_72021[add_78314 > 32'h0000_0009 ? 4'h9 : add_78314[3:0]];
  assign array_index_78318 = array_update_78315[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_78322 = smul32b_32b_x_32b(array_index_77428[add_78314 > 32'h0000_0009 ? 4'h9 : add_78314[3:0]], array_index_78317[add_78234 > 32'h0000_0009 ? 4'h9 : add_78234[3:0]]);
  assign add_78324 = array_index_78318[add_78234 > 32'h0000_0009 ? 4'h9 : add_78234[3:0]] + smul_78322;
  assign array_update_78326[0] = add_78234 == 32'h0000_0000 ? add_78324 : array_index_78318[0];
  assign array_update_78326[1] = add_78234 == 32'h0000_0001 ? add_78324 : array_index_78318[1];
  assign array_update_78326[2] = add_78234 == 32'h0000_0002 ? add_78324 : array_index_78318[2];
  assign array_update_78326[3] = add_78234 == 32'h0000_0003 ? add_78324 : array_index_78318[3];
  assign array_update_78326[4] = add_78234 == 32'h0000_0004 ? add_78324 : array_index_78318[4];
  assign array_update_78326[5] = add_78234 == 32'h0000_0005 ? add_78324 : array_index_78318[5];
  assign array_update_78326[6] = add_78234 == 32'h0000_0006 ? add_78324 : array_index_78318[6];
  assign array_update_78326[7] = add_78234 == 32'h0000_0007 ? add_78324 : array_index_78318[7];
  assign array_update_78326[8] = add_78234 == 32'h0000_0008 ? add_78324 : array_index_78318[8];
  assign array_update_78326[9] = add_78234 == 32'h0000_0009 ? add_78324 : array_index_78318[9];
  assign add_78327 = add_78314 + 32'h0000_0001;
  assign array_update_78328[0] = add_77421 == 32'h0000_0000 ? array_update_78326 : array_update_78315[0];
  assign array_update_78328[1] = add_77421 == 32'h0000_0001 ? array_update_78326 : array_update_78315[1];
  assign array_update_78328[2] = add_77421 == 32'h0000_0002 ? array_update_78326 : array_update_78315[2];
  assign array_update_78328[3] = add_77421 == 32'h0000_0003 ? array_update_78326 : array_update_78315[3];
  assign array_update_78328[4] = add_77421 == 32'h0000_0004 ? array_update_78326 : array_update_78315[4];
  assign array_update_78328[5] = add_77421 == 32'h0000_0005 ? array_update_78326 : array_update_78315[5];
  assign array_update_78328[6] = add_77421 == 32'h0000_0006 ? array_update_78326 : array_update_78315[6];
  assign array_update_78328[7] = add_77421 == 32'h0000_0007 ? array_update_78326 : array_update_78315[7];
  assign array_update_78328[8] = add_77421 == 32'h0000_0008 ? array_update_78326 : array_update_78315[8];
  assign array_update_78328[9] = add_77421 == 32'h0000_0009 ? array_update_78326 : array_update_78315[9];
  assign array_index_78330 = array_update_72021[add_78327 > 32'h0000_0009 ? 4'h9 : add_78327[3:0]];
  assign array_index_78331 = array_update_78328[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_78335 = smul32b_32b_x_32b(array_index_77428[add_78327 > 32'h0000_0009 ? 4'h9 : add_78327[3:0]], array_index_78330[add_78234 > 32'h0000_0009 ? 4'h9 : add_78234[3:0]]);
  assign add_78337 = array_index_78331[add_78234 > 32'h0000_0009 ? 4'h9 : add_78234[3:0]] + smul_78335;
  assign array_update_78339[0] = add_78234 == 32'h0000_0000 ? add_78337 : array_index_78331[0];
  assign array_update_78339[1] = add_78234 == 32'h0000_0001 ? add_78337 : array_index_78331[1];
  assign array_update_78339[2] = add_78234 == 32'h0000_0002 ? add_78337 : array_index_78331[2];
  assign array_update_78339[3] = add_78234 == 32'h0000_0003 ? add_78337 : array_index_78331[3];
  assign array_update_78339[4] = add_78234 == 32'h0000_0004 ? add_78337 : array_index_78331[4];
  assign array_update_78339[5] = add_78234 == 32'h0000_0005 ? add_78337 : array_index_78331[5];
  assign array_update_78339[6] = add_78234 == 32'h0000_0006 ? add_78337 : array_index_78331[6];
  assign array_update_78339[7] = add_78234 == 32'h0000_0007 ? add_78337 : array_index_78331[7];
  assign array_update_78339[8] = add_78234 == 32'h0000_0008 ? add_78337 : array_index_78331[8];
  assign array_update_78339[9] = add_78234 == 32'h0000_0009 ? add_78337 : array_index_78331[9];
  assign add_78340 = add_78327 + 32'h0000_0001;
  assign array_update_78341[0] = add_77421 == 32'h0000_0000 ? array_update_78339 : array_update_78328[0];
  assign array_update_78341[1] = add_77421 == 32'h0000_0001 ? array_update_78339 : array_update_78328[1];
  assign array_update_78341[2] = add_77421 == 32'h0000_0002 ? array_update_78339 : array_update_78328[2];
  assign array_update_78341[3] = add_77421 == 32'h0000_0003 ? array_update_78339 : array_update_78328[3];
  assign array_update_78341[4] = add_77421 == 32'h0000_0004 ? array_update_78339 : array_update_78328[4];
  assign array_update_78341[5] = add_77421 == 32'h0000_0005 ? array_update_78339 : array_update_78328[5];
  assign array_update_78341[6] = add_77421 == 32'h0000_0006 ? array_update_78339 : array_update_78328[6];
  assign array_update_78341[7] = add_77421 == 32'h0000_0007 ? array_update_78339 : array_update_78328[7];
  assign array_update_78341[8] = add_77421 == 32'h0000_0008 ? array_update_78339 : array_update_78328[8];
  assign array_update_78341[9] = add_77421 == 32'h0000_0009 ? array_update_78339 : array_update_78328[9];
  assign array_index_78343 = array_update_72021[add_78340 > 32'h0000_0009 ? 4'h9 : add_78340[3:0]];
  assign array_index_78344 = array_update_78341[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_78348 = smul32b_32b_x_32b(array_index_77428[add_78340 > 32'h0000_0009 ? 4'h9 : add_78340[3:0]], array_index_78343[add_78234 > 32'h0000_0009 ? 4'h9 : add_78234[3:0]]);
  assign add_78350 = array_index_78344[add_78234 > 32'h0000_0009 ? 4'h9 : add_78234[3:0]] + smul_78348;
  assign array_update_78352[0] = add_78234 == 32'h0000_0000 ? add_78350 : array_index_78344[0];
  assign array_update_78352[1] = add_78234 == 32'h0000_0001 ? add_78350 : array_index_78344[1];
  assign array_update_78352[2] = add_78234 == 32'h0000_0002 ? add_78350 : array_index_78344[2];
  assign array_update_78352[3] = add_78234 == 32'h0000_0003 ? add_78350 : array_index_78344[3];
  assign array_update_78352[4] = add_78234 == 32'h0000_0004 ? add_78350 : array_index_78344[4];
  assign array_update_78352[5] = add_78234 == 32'h0000_0005 ? add_78350 : array_index_78344[5];
  assign array_update_78352[6] = add_78234 == 32'h0000_0006 ? add_78350 : array_index_78344[6];
  assign array_update_78352[7] = add_78234 == 32'h0000_0007 ? add_78350 : array_index_78344[7];
  assign array_update_78352[8] = add_78234 == 32'h0000_0008 ? add_78350 : array_index_78344[8];
  assign array_update_78352[9] = add_78234 == 32'h0000_0009 ? add_78350 : array_index_78344[9];
  assign add_78353 = add_78340 + 32'h0000_0001;
  assign array_update_78354[0] = add_77421 == 32'h0000_0000 ? array_update_78352 : array_update_78341[0];
  assign array_update_78354[1] = add_77421 == 32'h0000_0001 ? array_update_78352 : array_update_78341[1];
  assign array_update_78354[2] = add_77421 == 32'h0000_0002 ? array_update_78352 : array_update_78341[2];
  assign array_update_78354[3] = add_77421 == 32'h0000_0003 ? array_update_78352 : array_update_78341[3];
  assign array_update_78354[4] = add_77421 == 32'h0000_0004 ? array_update_78352 : array_update_78341[4];
  assign array_update_78354[5] = add_77421 == 32'h0000_0005 ? array_update_78352 : array_update_78341[5];
  assign array_update_78354[6] = add_77421 == 32'h0000_0006 ? array_update_78352 : array_update_78341[6];
  assign array_update_78354[7] = add_77421 == 32'h0000_0007 ? array_update_78352 : array_update_78341[7];
  assign array_update_78354[8] = add_77421 == 32'h0000_0008 ? array_update_78352 : array_update_78341[8];
  assign array_update_78354[9] = add_77421 == 32'h0000_0009 ? array_update_78352 : array_update_78341[9];
  assign array_index_78356 = array_update_72021[add_78353 > 32'h0000_0009 ? 4'h9 : add_78353[3:0]];
  assign array_index_78357 = array_update_78354[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_78361 = smul32b_32b_x_32b(array_index_77428[add_78353 > 32'h0000_0009 ? 4'h9 : add_78353[3:0]], array_index_78356[add_78234 > 32'h0000_0009 ? 4'h9 : add_78234[3:0]]);
  assign add_78363 = array_index_78357[add_78234 > 32'h0000_0009 ? 4'h9 : add_78234[3:0]] + smul_78361;
  assign array_update_78364[0] = add_78234 == 32'h0000_0000 ? add_78363 : array_index_78357[0];
  assign array_update_78364[1] = add_78234 == 32'h0000_0001 ? add_78363 : array_index_78357[1];
  assign array_update_78364[2] = add_78234 == 32'h0000_0002 ? add_78363 : array_index_78357[2];
  assign array_update_78364[3] = add_78234 == 32'h0000_0003 ? add_78363 : array_index_78357[3];
  assign array_update_78364[4] = add_78234 == 32'h0000_0004 ? add_78363 : array_index_78357[4];
  assign array_update_78364[5] = add_78234 == 32'h0000_0005 ? add_78363 : array_index_78357[5];
  assign array_update_78364[6] = add_78234 == 32'h0000_0006 ? add_78363 : array_index_78357[6];
  assign array_update_78364[7] = add_78234 == 32'h0000_0007 ? add_78363 : array_index_78357[7];
  assign array_update_78364[8] = add_78234 == 32'h0000_0008 ? add_78363 : array_index_78357[8];
  assign array_update_78364[9] = add_78234 == 32'h0000_0009 ? add_78363 : array_index_78357[9];
  assign array_update_78365[0] = add_77421 == 32'h0000_0000 ? array_update_78364 : array_update_78354[0];
  assign array_update_78365[1] = add_77421 == 32'h0000_0001 ? array_update_78364 : array_update_78354[1];
  assign array_update_78365[2] = add_77421 == 32'h0000_0002 ? array_update_78364 : array_update_78354[2];
  assign array_update_78365[3] = add_77421 == 32'h0000_0003 ? array_update_78364 : array_update_78354[3];
  assign array_update_78365[4] = add_77421 == 32'h0000_0004 ? array_update_78364 : array_update_78354[4];
  assign array_update_78365[5] = add_77421 == 32'h0000_0005 ? array_update_78364 : array_update_78354[5];
  assign array_update_78365[6] = add_77421 == 32'h0000_0006 ? array_update_78364 : array_update_78354[6];
  assign array_update_78365[7] = add_77421 == 32'h0000_0007 ? array_update_78364 : array_update_78354[7];
  assign array_update_78365[8] = add_77421 == 32'h0000_0008 ? array_update_78364 : array_update_78354[8];
  assign array_update_78365[9] = add_77421 == 32'h0000_0009 ? array_update_78364 : array_update_78354[9];
  assign array_index_78367 = array_update_78365[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign add_78369 = add_78234 + 32'h0000_0001;
  assign array_update_78370[0] = add_78369 == 32'h0000_0000 ? 32'h0000_0000 : array_index_78367[0];
  assign array_update_78370[1] = add_78369 == 32'h0000_0001 ? 32'h0000_0000 : array_index_78367[1];
  assign array_update_78370[2] = add_78369 == 32'h0000_0002 ? 32'h0000_0000 : array_index_78367[2];
  assign array_update_78370[3] = add_78369 == 32'h0000_0003 ? 32'h0000_0000 : array_index_78367[3];
  assign array_update_78370[4] = add_78369 == 32'h0000_0004 ? 32'h0000_0000 : array_index_78367[4];
  assign array_update_78370[5] = add_78369 == 32'h0000_0005 ? 32'h0000_0000 : array_index_78367[5];
  assign array_update_78370[6] = add_78369 == 32'h0000_0006 ? 32'h0000_0000 : array_index_78367[6];
  assign array_update_78370[7] = add_78369 == 32'h0000_0007 ? 32'h0000_0000 : array_index_78367[7];
  assign array_update_78370[8] = add_78369 == 32'h0000_0008 ? 32'h0000_0000 : array_index_78367[8];
  assign array_update_78370[9] = add_78369 == 32'h0000_0009 ? 32'h0000_0000 : array_index_78367[9];
  assign literal_78371 = 32'h0000_0000;
  assign array_update_78372[0] = add_77421 == 32'h0000_0000 ? array_update_78370 : array_update_78365[0];
  assign array_update_78372[1] = add_77421 == 32'h0000_0001 ? array_update_78370 : array_update_78365[1];
  assign array_update_78372[2] = add_77421 == 32'h0000_0002 ? array_update_78370 : array_update_78365[2];
  assign array_update_78372[3] = add_77421 == 32'h0000_0003 ? array_update_78370 : array_update_78365[3];
  assign array_update_78372[4] = add_77421 == 32'h0000_0004 ? array_update_78370 : array_update_78365[4];
  assign array_update_78372[5] = add_77421 == 32'h0000_0005 ? array_update_78370 : array_update_78365[5];
  assign array_update_78372[6] = add_77421 == 32'h0000_0006 ? array_update_78370 : array_update_78365[6];
  assign array_update_78372[7] = add_77421 == 32'h0000_0007 ? array_update_78370 : array_update_78365[7];
  assign array_update_78372[8] = add_77421 == 32'h0000_0008 ? array_update_78370 : array_update_78365[8];
  assign array_update_78372[9] = add_77421 == 32'h0000_0009 ? array_update_78370 : array_update_78365[9];
  assign array_index_78374 = array_update_72021[literal_78371 > 32'h0000_0009 ? 4'h9 : literal_78371[3:0]];
  assign array_index_78375 = array_update_78372[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_78379 = smul32b_32b_x_32b(array_index_77428[literal_78371 > 32'h0000_0009 ? 4'h9 : literal_78371[3:0]], array_index_78374[add_78369 > 32'h0000_0009 ? 4'h9 : add_78369[3:0]]);
  assign add_78381 = array_index_78375[add_78369 > 32'h0000_0009 ? 4'h9 : add_78369[3:0]] + smul_78379;
  assign array_update_78383[0] = add_78369 == 32'h0000_0000 ? add_78381 : array_index_78375[0];
  assign array_update_78383[1] = add_78369 == 32'h0000_0001 ? add_78381 : array_index_78375[1];
  assign array_update_78383[2] = add_78369 == 32'h0000_0002 ? add_78381 : array_index_78375[2];
  assign array_update_78383[3] = add_78369 == 32'h0000_0003 ? add_78381 : array_index_78375[3];
  assign array_update_78383[4] = add_78369 == 32'h0000_0004 ? add_78381 : array_index_78375[4];
  assign array_update_78383[5] = add_78369 == 32'h0000_0005 ? add_78381 : array_index_78375[5];
  assign array_update_78383[6] = add_78369 == 32'h0000_0006 ? add_78381 : array_index_78375[6];
  assign array_update_78383[7] = add_78369 == 32'h0000_0007 ? add_78381 : array_index_78375[7];
  assign array_update_78383[8] = add_78369 == 32'h0000_0008 ? add_78381 : array_index_78375[8];
  assign array_update_78383[9] = add_78369 == 32'h0000_0009 ? add_78381 : array_index_78375[9];
  assign add_78384 = literal_78371 + 32'h0000_0001;
  assign array_update_78385[0] = add_77421 == 32'h0000_0000 ? array_update_78383 : array_update_78372[0];
  assign array_update_78385[1] = add_77421 == 32'h0000_0001 ? array_update_78383 : array_update_78372[1];
  assign array_update_78385[2] = add_77421 == 32'h0000_0002 ? array_update_78383 : array_update_78372[2];
  assign array_update_78385[3] = add_77421 == 32'h0000_0003 ? array_update_78383 : array_update_78372[3];
  assign array_update_78385[4] = add_77421 == 32'h0000_0004 ? array_update_78383 : array_update_78372[4];
  assign array_update_78385[5] = add_77421 == 32'h0000_0005 ? array_update_78383 : array_update_78372[5];
  assign array_update_78385[6] = add_77421 == 32'h0000_0006 ? array_update_78383 : array_update_78372[6];
  assign array_update_78385[7] = add_77421 == 32'h0000_0007 ? array_update_78383 : array_update_78372[7];
  assign array_update_78385[8] = add_77421 == 32'h0000_0008 ? array_update_78383 : array_update_78372[8];
  assign array_update_78385[9] = add_77421 == 32'h0000_0009 ? array_update_78383 : array_update_78372[9];
  assign array_index_78387 = array_update_72021[add_78384 > 32'h0000_0009 ? 4'h9 : add_78384[3:0]];
  assign array_index_78388 = array_update_78385[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_78392 = smul32b_32b_x_32b(array_index_77428[add_78384 > 32'h0000_0009 ? 4'h9 : add_78384[3:0]], array_index_78387[add_78369 > 32'h0000_0009 ? 4'h9 : add_78369[3:0]]);
  assign add_78394 = array_index_78388[add_78369 > 32'h0000_0009 ? 4'h9 : add_78369[3:0]] + smul_78392;
  assign array_update_78396[0] = add_78369 == 32'h0000_0000 ? add_78394 : array_index_78388[0];
  assign array_update_78396[1] = add_78369 == 32'h0000_0001 ? add_78394 : array_index_78388[1];
  assign array_update_78396[2] = add_78369 == 32'h0000_0002 ? add_78394 : array_index_78388[2];
  assign array_update_78396[3] = add_78369 == 32'h0000_0003 ? add_78394 : array_index_78388[3];
  assign array_update_78396[4] = add_78369 == 32'h0000_0004 ? add_78394 : array_index_78388[4];
  assign array_update_78396[5] = add_78369 == 32'h0000_0005 ? add_78394 : array_index_78388[5];
  assign array_update_78396[6] = add_78369 == 32'h0000_0006 ? add_78394 : array_index_78388[6];
  assign array_update_78396[7] = add_78369 == 32'h0000_0007 ? add_78394 : array_index_78388[7];
  assign array_update_78396[8] = add_78369 == 32'h0000_0008 ? add_78394 : array_index_78388[8];
  assign array_update_78396[9] = add_78369 == 32'h0000_0009 ? add_78394 : array_index_78388[9];
  assign add_78397 = add_78384 + 32'h0000_0001;
  assign array_update_78398[0] = add_77421 == 32'h0000_0000 ? array_update_78396 : array_update_78385[0];
  assign array_update_78398[1] = add_77421 == 32'h0000_0001 ? array_update_78396 : array_update_78385[1];
  assign array_update_78398[2] = add_77421 == 32'h0000_0002 ? array_update_78396 : array_update_78385[2];
  assign array_update_78398[3] = add_77421 == 32'h0000_0003 ? array_update_78396 : array_update_78385[3];
  assign array_update_78398[4] = add_77421 == 32'h0000_0004 ? array_update_78396 : array_update_78385[4];
  assign array_update_78398[5] = add_77421 == 32'h0000_0005 ? array_update_78396 : array_update_78385[5];
  assign array_update_78398[6] = add_77421 == 32'h0000_0006 ? array_update_78396 : array_update_78385[6];
  assign array_update_78398[7] = add_77421 == 32'h0000_0007 ? array_update_78396 : array_update_78385[7];
  assign array_update_78398[8] = add_77421 == 32'h0000_0008 ? array_update_78396 : array_update_78385[8];
  assign array_update_78398[9] = add_77421 == 32'h0000_0009 ? array_update_78396 : array_update_78385[9];
  assign array_index_78400 = array_update_72021[add_78397 > 32'h0000_0009 ? 4'h9 : add_78397[3:0]];
  assign array_index_78401 = array_update_78398[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_78405 = smul32b_32b_x_32b(array_index_77428[add_78397 > 32'h0000_0009 ? 4'h9 : add_78397[3:0]], array_index_78400[add_78369 > 32'h0000_0009 ? 4'h9 : add_78369[3:0]]);
  assign add_78407 = array_index_78401[add_78369 > 32'h0000_0009 ? 4'h9 : add_78369[3:0]] + smul_78405;
  assign array_update_78409[0] = add_78369 == 32'h0000_0000 ? add_78407 : array_index_78401[0];
  assign array_update_78409[1] = add_78369 == 32'h0000_0001 ? add_78407 : array_index_78401[1];
  assign array_update_78409[2] = add_78369 == 32'h0000_0002 ? add_78407 : array_index_78401[2];
  assign array_update_78409[3] = add_78369 == 32'h0000_0003 ? add_78407 : array_index_78401[3];
  assign array_update_78409[4] = add_78369 == 32'h0000_0004 ? add_78407 : array_index_78401[4];
  assign array_update_78409[5] = add_78369 == 32'h0000_0005 ? add_78407 : array_index_78401[5];
  assign array_update_78409[6] = add_78369 == 32'h0000_0006 ? add_78407 : array_index_78401[6];
  assign array_update_78409[7] = add_78369 == 32'h0000_0007 ? add_78407 : array_index_78401[7];
  assign array_update_78409[8] = add_78369 == 32'h0000_0008 ? add_78407 : array_index_78401[8];
  assign array_update_78409[9] = add_78369 == 32'h0000_0009 ? add_78407 : array_index_78401[9];
  assign add_78410 = add_78397 + 32'h0000_0001;
  assign array_update_78411[0] = add_77421 == 32'h0000_0000 ? array_update_78409 : array_update_78398[0];
  assign array_update_78411[1] = add_77421 == 32'h0000_0001 ? array_update_78409 : array_update_78398[1];
  assign array_update_78411[2] = add_77421 == 32'h0000_0002 ? array_update_78409 : array_update_78398[2];
  assign array_update_78411[3] = add_77421 == 32'h0000_0003 ? array_update_78409 : array_update_78398[3];
  assign array_update_78411[4] = add_77421 == 32'h0000_0004 ? array_update_78409 : array_update_78398[4];
  assign array_update_78411[5] = add_77421 == 32'h0000_0005 ? array_update_78409 : array_update_78398[5];
  assign array_update_78411[6] = add_77421 == 32'h0000_0006 ? array_update_78409 : array_update_78398[6];
  assign array_update_78411[7] = add_77421 == 32'h0000_0007 ? array_update_78409 : array_update_78398[7];
  assign array_update_78411[8] = add_77421 == 32'h0000_0008 ? array_update_78409 : array_update_78398[8];
  assign array_update_78411[9] = add_77421 == 32'h0000_0009 ? array_update_78409 : array_update_78398[9];
  assign array_index_78413 = array_update_72021[add_78410 > 32'h0000_0009 ? 4'h9 : add_78410[3:0]];
  assign array_index_78414 = array_update_78411[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_78418 = smul32b_32b_x_32b(array_index_77428[add_78410 > 32'h0000_0009 ? 4'h9 : add_78410[3:0]], array_index_78413[add_78369 > 32'h0000_0009 ? 4'h9 : add_78369[3:0]]);
  assign add_78420 = array_index_78414[add_78369 > 32'h0000_0009 ? 4'h9 : add_78369[3:0]] + smul_78418;
  assign array_update_78422[0] = add_78369 == 32'h0000_0000 ? add_78420 : array_index_78414[0];
  assign array_update_78422[1] = add_78369 == 32'h0000_0001 ? add_78420 : array_index_78414[1];
  assign array_update_78422[2] = add_78369 == 32'h0000_0002 ? add_78420 : array_index_78414[2];
  assign array_update_78422[3] = add_78369 == 32'h0000_0003 ? add_78420 : array_index_78414[3];
  assign array_update_78422[4] = add_78369 == 32'h0000_0004 ? add_78420 : array_index_78414[4];
  assign array_update_78422[5] = add_78369 == 32'h0000_0005 ? add_78420 : array_index_78414[5];
  assign array_update_78422[6] = add_78369 == 32'h0000_0006 ? add_78420 : array_index_78414[6];
  assign array_update_78422[7] = add_78369 == 32'h0000_0007 ? add_78420 : array_index_78414[7];
  assign array_update_78422[8] = add_78369 == 32'h0000_0008 ? add_78420 : array_index_78414[8];
  assign array_update_78422[9] = add_78369 == 32'h0000_0009 ? add_78420 : array_index_78414[9];
  assign add_78423 = add_78410 + 32'h0000_0001;
  assign array_update_78424[0] = add_77421 == 32'h0000_0000 ? array_update_78422 : array_update_78411[0];
  assign array_update_78424[1] = add_77421 == 32'h0000_0001 ? array_update_78422 : array_update_78411[1];
  assign array_update_78424[2] = add_77421 == 32'h0000_0002 ? array_update_78422 : array_update_78411[2];
  assign array_update_78424[3] = add_77421 == 32'h0000_0003 ? array_update_78422 : array_update_78411[3];
  assign array_update_78424[4] = add_77421 == 32'h0000_0004 ? array_update_78422 : array_update_78411[4];
  assign array_update_78424[5] = add_77421 == 32'h0000_0005 ? array_update_78422 : array_update_78411[5];
  assign array_update_78424[6] = add_77421 == 32'h0000_0006 ? array_update_78422 : array_update_78411[6];
  assign array_update_78424[7] = add_77421 == 32'h0000_0007 ? array_update_78422 : array_update_78411[7];
  assign array_update_78424[8] = add_77421 == 32'h0000_0008 ? array_update_78422 : array_update_78411[8];
  assign array_update_78424[9] = add_77421 == 32'h0000_0009 ? array_update_78422 : array_update_78411[9];
  assign array_index_78426 = array_update_72021[add_78423 > 32'h0000_0009 ? 4'h9 : add_78423[3:0]];
  assign array_index_78427 = array_update_78424[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_78431 = smul32b_32b_x_32b(array_index_77428[add_78423 > 32'h0000_0009 ? 4'h9 : add_78423[3:0]], array_index_78426[add_78369 > 32'h0000_0009 ? 4'h9 : add_78369[3:0]]);
  assign add_78433 = array_index_78427[add_78369 > 32'h0000_0009 ? 4'h9 : add_78369[3:0]] + smul_78431;
  assign array_update_78435[0] = add_78369 == 32'h0000_0000 ? add_78433 : array_index_78427[0];
  assign array_update_78435[1] = add_78369 == 32'h0000_0001 ? add_78433 : array_index_78427[1];
  assign array_update_78435[2] = add_78369 == 32'h0000_0002 ? add_78433 : array_index_78427[2];
  assign array_update_78435[3] = add_78369 == 32'h0000_0003 ? add_78433 : array_index_78427[3];
  assign array_update_78435[4] = add_78369 == 32'h0000_0004 ? add_78433 : array_index_78427[4];
  assign array_update_78435[5] = add_78369 == 32'h0000_0005 ? add_78433 : array_index_78427[5];
  assign array_update_78435[6] = add_78369 == 32'h0000_0006 ? add_78433 : array_index_78427[6];
  assign array_update_78435[7] = add_78369 == 32'h0000_0007 ? add_78433 : array_index_78427[7];
  assign array_update_78435[8] = add_78369 == 32'h0000_0008 ? add_78433 : array_index_78427[8];
  assign array_update_78435[9] = add_78369 == 32'h0000_0009 ? add_78433 : array_index_78427[9];
  assign add_78436 = add_78423 + 32'h0000_0001;
  assign array_update_78437[0] = add_77421 == 32'h0000_0000 ? array_update_78435 : array_update_78424[0];
  assign array_update_78437[1] = add_77421 == 32'h0000_0001 ? array_update_78435 : array_update_78424[1];
  assign array_update_78437[2] = add_77421 == 32'h0000_0002 ? array_update_78435 : array_update_78424[2];
  assign array_update_78437[3] = add_77421 == 32'h0000_0003 ? array_update_78435 : array_update_78424[3];
  assign array_update_78437[4] = add_77421 == 32'h0000_0004 ? array_update_78435 : array_update_78424[4];
  assign array_update_78437[5] = add_77421 == 32'h0000_0005 ? array_update_78435 : array_update_78424[5];
  assign array_update_78437[6] = add_77421 == 32'h0000_0006 ? array_update_78435 : array_update_78424[6];
  assign array_update_78437[7] = add_77421 == 32'h0000_0007 ? array_update_78435 : array_update_78424[7];
  assign array_update_78437[8] = add_77421 == 32'h0000_0008 ? array_update_78435 : array_update_78424[8];
  assign array_update_78437[9] = add_77421 == 32'h0000_0009 ? array_update_78435 : array_update_78424[9];
  assign array_index_78439 = array_update_72021[add_78436 > 32'h0000_0009 ? 4'h9 : add_78436[3:0]];
  assign array_index_78440 = array_update_78437[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_78444 = smul32b_32b_x_32b(array_index_77428[add_78436 > 32'h0000_0009 ? 4'h9 : add_78436[3:0]], array_index_78439[add_78369 > 32'h0000_0009 ? 4'h9 : add_78369[3:0]]);
  assign add_78446 = array_index_78440[add_78369 > 32'h0000_0009 ? 4'h9 : add_78369[3:0]] + smul_78444;
  assign array_update_78448[0] = add_78369 == 32'h0000_0000 ? add_78446 : array_index_78440[0];
  assign array_update_78448[1] = add_78369 == 32'h0000_0001 ? add_78446 : array_index_78440[1];
  assign array_update_78448[2] = add_78369 == 32'h0000_0002 ? add_78446 : array_index_78440[2];
  assign array_update_78448[3] = add_78369 == 32'h0000_0003 ? add_78446 : array_index_78440[3];
  assign array_update_78448[4] = add_78369 == 32'h0000_0004 ? add_78446 : array_index_78440[4];
  assign array_update_78448[5] = add_78369 == 32'h0000_0005 ? add_78446 : array_index_78440[5];
  assign array_update_78448[6] = add_78369 == 32'h0000_0006 ? add_78446 : array_index_78440[6];
  assign array_update_78448[7] = add_78369 == 32'h0000_0007 ? add_78446 : array_index_78440[7];
  assign array_update_78448[8] = add_78369 == 32'h0000_0008 ? add_78446 : array_index_78440[8];
  assign array_update_78448[9] = add_78369 == 32'h0000_0009 ? add_78446 : array_index_78440[9];
  assign add_78449 = add_78436 + 32'h0000_0001;
  assign array_update_78450[0] = add_77421 == 32'h0000_0000 ? array_update_78448 : array_update_78437[0];
  assign array_update_78450[1] = add_77421 == 32'h0000_0001 ? array_update_78448 : array_update_78437[1];
  assign array_update_78450[2] = add_77421 == 32'h0000_0002 ? array_update_78448 : array_update_78437[2];
  assign array_update_78450[3] = add_77421 == 32'h0000_0003 ? array_update_78448 : array_update_78437[3];
  assign array_update_78450[4] = add_77421 == 32'h0000_0004 ? array_update_78448 : array_update_78437[4];
  assign array_update_78450[5] = add_77421 == 32'h0000_0005 ? array_update_78448 : array_update_78437[5];
  assign array_update_78450[6] = add_77421 == 32'h0000_0006 ? array_update_78448 : array_update_78437[6];
  assign array_update_78450[7] = add_77421 == 32'h0000_0007 ? array_update_78448 : array_update_78437[7];
  assign array_update_78450[8] = add_77421 == 32'h0000_0008 ? array_update_78448 : array_update_78437[8];
  assign array_update_78450[9] = add_77421 == 32'h0000_0009 ? array_update_78448 : array_update_78437[9];
  assign array_index_78452 = array_update_72021[add_78449 > 32'h0000_0009 ? 4'h9 : add_78449[3:0]];
  assign array_index_78453 = array_update_78450[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_78457 = smul32b_32b_x_32b(array_index_77428[add_78449 > 32'h0000_0009 ? 4'h9 : add_78449[3:0]], array_index_78452[add_78369 > 32'h0000_0009 ? 4'h9 : add_78369[3:0]]);
  assign add_78459 = array_index_78453[add_78369 > 32'h0000_0009 ? 4'h9 : add_78369[3:0]] + smul_78457;
  assign array_update_78461[0] = add_78369 == 32'h0000_0000 ? add_78459 : array_index_78453[0];
  assign array_update_78461[1] = add_78369 == 32'h0000_0001 ? add_78459 : array_index_78453[1];
  assign array_update_78461[2] = add_78369 == 32'h0000_0002 ? add_78459 : array_index_78453[2];
  assign array_update_78461[3] = add_78369 == 32'h0000_0003 ? add_78459 : array_index_78453[3];
  assign array_update_78461[4] = add_78369 == 32'h0000_0004 ? add_78459 : array_index_78453[4];
  assign array_update_78461[5] = add_78369 == 32'h0000_0005 ? add_78459 : array_index_78453[5];
  assign array_update_78461[6] = add_78369 == 32'h0000_0006 ? add_78459 : array_index_78453[6];
  assign array_update_78461[7] = add_78369 == 32'h0000_0007 ? add_78459 : array_index_78453[7];
  assign array_update_78461[8] = add_78369 == 32'h0000_0008 ? add_78459 : array_index_78453[8];
  assign array_update_78461[9] = add_78369 == 32'h0000_0009 ? add_78459 : array_index_78453[9];
  assign add_78462 = add_78449 + 32'h0000_0001;
  assign array_update_78463[0] = add_77421 == 32'h0000_0000 ? array_update_78461 : array_update_78450[0];
  assign array_update_78463[1] = add_77421 == 32'h0000_0001 ? array_update_78461 : array_update_78450[1];
  assign array_update_78463[2] = add_77421 == 32'h0000_0002 ? array_update_78461 : array_update_78450[2];
  assign array_update_78463[3] = add_77421 == 32'h0000_0003 ? array_update_78461 : array_update_78450[3];
  assign array_update_78463[4] = add_77421 == 32'h0000_0004 ? array_update_78461 : array_update_78450[4];
  assign array_update_78463[5] = add_77421 == 32'h0000_0005 ? array_update_78461 : array_update_78450[5];
  assign array_update_78463[6] = add_77421 == 32'h0000_0006 ? array_update_78461 : array_update_78450[6];
  assign array_update_78463[7] = add_77421 == 32'h0000_0007 ? array_update_78461 : array_update_78450[7];
  assign array_update_78463[8] = add_77421 == 32'h0000_0008 ? array_update_78461 : array_update_78450[8];
  assign array_update_78463[9] = add_77421 == 32'h0000_0009 ? array_update_78461 : array_update_78450[9];
  assign array_index_78465 = array_update_72021[add_78462 > 32'h0000_0009 ? 4'h9 : add_78462[3:0]];
  assign array_index_78466 = array_update_78463[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_78470 = smul32b_32b_x_32b(array_index_77428[add_78462 > 32'h0000_0009 ? 4'h9 : add_78462[3:0]], array_index_78465[add_78369 > 32'h0000_0009 ? 4'h9 : add_78369[3:0]]);
  assign add_78472 = array_index_78466[add_78369 > 32'h0000_0009 ? 4'h9 : add_78369[3:0]] + smul_78470;
  assign array_update_78474[0] = add_78369 == 32'h0000_0000 ? add_78472 : array_index_78466[0];
  assign array_update_78474[1] = add_78369 == 32'h0000_0001 ? add_78472 : array_index_78466[1];
  assign array_update_78474[2] = add_78369 == 32'h0000_0002 ? add_78472 : array_index_78466[2];
  assign array_update_78474[3] = add_78369 == 32'h0000_0003 ? add_78472 : array_index_78466[3];
  assign array_update_78474[4] = add_78369 == 32'h0000_0004 ? add_78472 : array_index_78466[4];
  assign array_update_78474[5] = add_78369 == 32'h0000_0005 ? add_78472 : array_index_78466[5];
  assign array_update_78474[6] = add_78369 == 32'h0000_0006 ? add_78472 : array_index_78466[6];
  assign array_update_78474[7] = add_78369 == 32'h0000_0007 ? add_78472 : array_index_78466[7];
  assign array_update_78474[8] = add_78369 == 32'h0000_0008 ? add_78472 : array_index_78466[8];
  assign array_update_78474[9] = add_78369 == 32'h0000_0009 ? add_78472 : array_index_78466[9];
  assign add_78475 = add_78462 + 32'h0000_0001;
  assign array_update_78476[0] = add_77421 == 32'h0000_0000 ? array_update_78474 : array_update_78463[0];
  assign array_update_78476[1] = add_77421 == 32'h0000_0001 ? array_update_78474 : array_update_78463[1];
  assign array_update_78476[2] = add_77421 == 32'h0000_0002 ? array_update_78474 : array_update_78463[2];
  assign array_update_78476[3] = add_77421 == 32'h0000_0003 ? array_update_78474 : array_update_78463[3];
  assign array_update_78476[4] = add_77421 == 32'h0000_0004 ? array_update_78474 : array_update_78463[4];
  assign array_update_78476[5] = add_77421 == 32'h0000_0005 ? array_update_78474 : array_update_78463[5];
  assign array_update_78476[6] = add_77421 == 32'h0000_0006 ? array_update_78474 : array_update_78463[6];
  assign array_update_78476[7] = add_77421 == 32'h0000_0007 ? array_update_78474 : array_update_78463[7];
  assign array_update_78476[8] = add_77421 == 32'h0000_0008 ? array_update_78474 : array_update_78463[8];
  assign array_update_78476[9] = add_77421 == 32'h0000_0009 ? array_update_78474 : array_update_78463[9];
  assign array_index_78478 = array_update_72021[add_78475 > 32'h0000_0009 ? 4'h9 : add_78475[3:0]];
  assign array_index_78479 = array_update_78476[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_78483 = smul32b_32b_x_32b(array_index_77428[add_78475 > 32'h0000_0009 ? 4'h9 : add_78475[3:0]], array_index_78478[add_78369 > 32'h0000_0009 ? 4'h9 : add_78369[3:0]]);
  assign add_78485 = array_index_78479[add_78369 > 32'h0000_0009 ? 4'h9 : add_78369[3:0]] + smul_78483;
  assign array_update_78487[0] = add_78369 == 32'h0000_0000 ? add_78485 : array_index_78479[0];
  assign array_update_78487[1] = add_78369 == 32'h0000_0001 ? add_78485 : array_index_78479[1];
  assign array_update_78487[2] = add_78369 == 32'h0000_0002 ? add_78485 : array_index_78479[2];
  assign array_update_78487[3] = add_78369 == 32'h0000_0003 ? add_78485 : array_index_78479[3];
  assign array_update_78487[4] = add_78369 == 32'h0000_0004 ? add_78485 : array_index_78479[4];
  assign array_update_78487[5] = add_78369 == 32'h0000_0005 ? add_78485 : array_index_78479[5];
  assign array_update_78487[6] = add_78369 == 32'h0000_0006 ? add_78485 : array_index_78479[6];
  assign array_update_78487[7] = add_78369 == 32'h0000_0007 ? add_78485 : array_index_78479[7];
  assign array_update_78487[8] = add_78369 == 32'h0000_0008 ? add_78485 : array_index_78479[8];
  assign array_update_78487[9] = add_78369 == 32'h0000_0009 ? add_78485 : array_index_78479[9];
  assign add_78488 = add_78475 + 32'h0000_0001;
  assign array_update_78489[0] = add_77421 == 32'h0000_0000 ? array_update_78487 : array_update_78476[0];
  assign array_update_78489[1] = add_77421 == 32'h0000_0001 ? array_update_78487 : array_update_78476[1];
  assign array_update_78489[2] = add_77421 == 32'h0000_0002 ? array_update_78487 : array_update_78476[2];
  assign array_update_78489[3] = add_77421 == 32'h0000_0003 ? array_update_78487 : array_update_78476[3];
  assign array_update_78489[4] = add_77421 == 32'h0000_0004 ? array_update_78487 : array_update_78476[4];
  assign array_update_78489[5] = add_77421 == 32'h0000_0005 ? array_update_78487 : array_update_78476[5];
  assign array_update_78489[6] = add_77421 == 32'h0000_0006 ? array_update_78487 : array_update_78476[6];
  assign array_update_78489[7] = add_77421 == 32'h0000_0007 ? array_update_78487 : array_update_78476[7];
  assign array_update_78489[8] = add_77421 == 32'h0000_0008 ? array_update_78487 : array_update_78476[8];
  assign array_update_78489[9] = add_77421 == 32'h0000_0009 ? array_update_78487 : array_update_78476[9];
  assign array_index_78491 = array_update_72021[add_78488 > 32'h0000_0009 ? 4'h9 : add_78488[3:0]];
  assign array_index_78492 = array_update_78489[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_78496 = smul32b_32b_x_32b(array_index_77428[add_78488 > 32'h0000_0009 ? 4'h9 : add_78488[3:0]], array_index_78491[add_78369 > 32'h0000_0009 ? 4'h9 : add_78369[3:0]]);
  assign add_78498 = array_index_78492[add_78369 > 32'h0000_0009 ? 4'h9 : add_78369[3:0]] + smul_78496;
  assign array_update_78499[0] = add_78369 == 32'h0000_0000 ? add_78498 : array_index_78492[0];
  assign array_update_78499[1] = add_78369 == 32'h0000_0001 ? add_78498 : array_index_78492[1];
  assign array_update_78499[2] = add_78369 == 32'h0000_0002 ? add_78498 : array_index_78492[2];
  assign array_update_78499[3] = add_78369 == 32'h0000_0003 ? add_78498 : array_index_78492[3];
  assign array_update_78499[4] = add_78369 == 32'h0000_0004 ? add_78498 : array_index_78492[4];
  assign array_update_78499[5] = add_78369 == 32'h0000_0005 ? add_78498 : array_index_78492[5];
  assign array_update_78499[6] = add_78369 == 32'h0000_0006 ? add_78498 : array_index_78492[6];
  assign array_update_78499[7] = add_78369 == 32'h0000_0007 ? add_78498 : array_index_78492[7];
  assign array_update_78499[8] = add_78369 == 32'h0000_0008 ? add_78498 : array_index_78492[8];
  assign array_update_78499[9] = add_78369 == 32'h0000_0009 ? add_78498 : array_index_78492[9];
  assign array_update_78500[0] = add_77421 == 32'h0000_0000 ? array_update_78499 : array_update_78489[0];
  assign array_update_78500[1] = add_77421 == 32'h0000_0001 ? array_update_78499 : array_update_78489[1];
  assign array_update_78500[2] = add_77421 == 32'h0000_0002 ? array_update_78499 : array_update_78489[2];
  assign array_update_78500[3] = add_77421 == 32'h0000_0003 ? array_update_78499 : array_update_78489[3];
  assign array_update_78500[4] = add_77421 == 32'h0000_0004 ? array_update_78499 : array_update_78489[4];
  assign array_update_78500[5] = add_77421 == 32'h0000_0005 ? array_update_78499 : array_update_78489[5];
  assign array_update_78500[6] = add_77421 == 32'h0000_0006 ? array_update_78499 : array_update_78489[6];
  assign array_update_78500[7] = add_77421 == 32'h0000_0007 ? array_update_78499 : array_update_78489[7];
  assign array_update_78500[8] = add_77421 == 32'h0000_0008 ? array_update_78499 : array_update_78489[8];
  assign array_update_78500[9] = add_77421 == 32'h0000_0009 ? array_update_78499 : array_update_78489[9];
  assign array_index_78502 = array_update_78500[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign add_78504 = add_78369 + 32'h0000_0001;
  assign array_update_78505[0] = add_78504 == 32'h0000_0000 ? 32'h0000_0000 : array_index_78502[0];
  assign array_update_78505[1] = add_78504 == 32'h0000_0001 ? 32'h0000_0000 : array_index_78502[1];
  assign array_update_78505[2] = add_78504 == 32'h0000_0002 ? 32'h0000_0000 : array_index_78502[2];
  assign array_update_78505[3] = add_78504 == 32'h0000_0003 ? 32'h0000_0000 : array_index_78502[3];
  assign array_update_78505[4] = add_78504 == 32'h0000_0004 ? 32'h0000_0000 : array_index_78502[4];
  assign array_update_78505[5] = add_78504 == 32'h0000_0005 ? 32'h0000_0000 : array_index_78502[5];
  assign array_update_78505[6] = add_78504 == 32'h0000_0006 ? 32'h0000_0000 : array_index_78502[6];
  assign array_update_78505[7] = add_78504 == 32'h0000_0007 ? 32'h0000_0000 : array_index_78502[7];
  assign array_update_78505[8] = add_78504 == 32'h0000_0008 ? 32'h0000_0000 : array_index_78502[8];
  assign array_update_78505[9] = add_78504 == 32'h0000_0009 ? 32'h0000_0000 : array_index_78502[9];
  assign literal_78506 = 32'h0000_0000;
  assign array_update_78507[0] = add_77421 == 32'h0000_0000 ? array_update_78505 : array_update_78500[0];
  assign array_update_78507[1] = add_77421 == 32'h0000_0001 ? array_update_78505 : array_update_78500[1];
  assign array_update_78507[2] = add_77421 == 32'h0000_0002 ? array_update_78505 : array_update_78500[2];
  assign array_update_78507[3] = add_77421 == 32'h0000_0003 ? array_update_78505 : array_update_78500[3];
  assign array_update_78507[4] = add_77421 == 32'h0000_0004 ? array_update_78505 : array_update_78500[4];
  assign array_update_78507[5] = add_77421 == 32'h0000_0005 ? array_update_78505 : array_update_78500[5];
  assign array_update_78507[6] = add_77421 == 32'h0000_0006 ? array_update_78505 : array_update_78500[6];
  assign array_update_78507[7] = add_77421 == 32'h0000_0007 ? array_update_78505 : array_update_78500[7];
  assign array_update_78507[8] = add_77421 == 32'h0000_0008 ? array_update_78505 : array_update_78500[8];
  assign array_update_78507[9] = add_77421 == 32'h0000_0009 ? array_update_78505 : array_update_78500[9];
  assign array_index_78509 = array_update_72021[literal_78506 > 32'h0000_0009 ? 4'h9 : literal_78506[3:0]];
  assign array_index_78510 = array_update_78507[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_78514 = smul32b_32b_x_32b(array_index_77428[literal_78506 > 32'h0000_0009 ? 4'h9 : literal_78506[3:0]], array_index_78509[add_78504 > 32'h0000_0009 ? 4'h9 : add_78504[3:0]]);
  assign add_78516 = array_index_78510[add_78504 > 32'h0000_0009 ? 4'h9 : add_78504[3:0]] + smul_78514;
  assign array_update_78518[0] = add_78504 == 32'h0000_0000 ? add_78516 : array_index_78510[0];
  assign array_update_78518[1] = add_78504 == 32'h0000_0001 ? add_78516 : array_index_78510[1];
  assign array_update_78518[2] = add_78504 == 32'h0000_0002 ? add_78516 : array_index_78510[2];
  assign array_update_78518[3] = add_78504 == 32'h0000_0003 ? add_78516 : array_index_78510[3];
  assign array_update_78518[4] = add_78504 == 32'h0000_0004 ? add_78516 : array_index_78510[4];
  assign array_update_78518[5] = add_78504 == 32'h0000_0005 ? add_78516 : array_index_78510[5];
  assign array_update_78518[6] = add_78504 == 32'h0000_0006 ? add_78516 : array_index_78510[6];
  assign array_update_78518[7] = add_78504 == 32'h0000_0007 ? add_78516 : array_index_78510[7];
  assign array_update_78518[8] = add_78504 == 32'h0000_0008 ? add_78516 : array_index_78510[8];
  assign array_update_78518[9] = add_78504 == 32'h0000_0009 ? add_78516 : array_index_78510[9];
  assign add_78519 = literal_78506 + 32'h0000_0001;
  assign array_update_78520[0] = add_77421 == 32'h0000_0000 ? array_update_78518 : array_update_78507[0];
  assign array_update_78520[1] = add_77421 == 32'h0000_0001 ? array_update_78518 : array_update_78507[1];
  assign array_update_78520[2] = add_77421 == 32'h0000_0002 ? array_update_78518 : array_update_78507[2];
  assign array_update_78520[3] = add_77421 == 32'h0000_0003 ? array_update_78518 : array_update_78507[3];
  assign array_update_78520[4] = add_77421 == 32'h0000_0004 ? array_update_78518 : array_update_78507[4];
  assign array_update_78520[5] = add_77421 == 32'h0000_0005 ? array_update_78518 : array_update_78507[5];
  assign array_update_78520[6] = add_77421 == 32'h0000_0006 ? array_update_78518 : array_update_78507[6];
  assign array_update_78520[7] = add_77421 == 32'h0000_0007 ? array_update_78518 : array_update_78507[7];
  assign array_update_78520[8] = add_77421 == 32'h0000_0008 ? array_update_78518 : array_update_78507[8];
  assign array_update_78520[9] = add_77421 == 32'h0000_0009 ? array_update_78518 : array_update_78507[9];
  assign array_index_78522 = array_update_72021[add_78519 > 32'h0000_0009 ? 4'h9 : add_78519[3:0]];
  assign array_index_78523 = array_update_78520[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_78527 = smul32b_32b_x_32b(array_index_77428[add_78519 > 32'h0000_0009 ? 4'h9 : add_78519[3:0]], array_index_78522[add_78504 > 32'h0000_0009 ? 4'h9 : add_78504[3:0]]);
  assign add_78529 = array_index_78523[add_78504 > 32'h0000_0009 ? 4'h9 : add_78504[3:0]] + smul_78527;
  assign array_update_78531[0] = add_78504 == 32'h0000_0000 ? add_78529 : array_index_78523[0];
  assign array_update_78531[1] = add_78504 == 32'h0000_0001 ? add_78529 : array_index_78523[1];
  assign array_update_78531[2] = add_78504 == 32'h0000_0002 ? add_78529 : array_index_78523[2];
  assign array_update_78531[3] = add_78504 == 32'h0000_0003 ? add_78529 : array_index_78523[3];
  assign array_update_78531[4] = add_78504 == 32'h0000_0004 ? add_78529 : array_index_78523[4];
  assign array_update_78531[5] = add_78504 == 32'h0000_0005 ? add_78529 : array_index_78523[5];
  assign array_update_78531[6] = add_78504 == 32'h0000_0006 ? add_78529 : array_index_78523[6];
  assign array_update_78531[7] = add_78504 == 32'h0000_0007 ? add_78529 : array_index_78523[7];
  assign array_update_78531[8] = add_78504 == 32'h0000_0008 ? add_78529 : array_index_78523[8];
  assign array_update_78531[9] = add_78504 == 32'h0000_0009 ? add_78529 : array_index_78523[9];
  assign add_78532 = add_78519 + 32'h0000_0001;
  assign array_update_78533[0] = add_77421 == 32'h0000_0000 ? array_update_78531 : array_update_78520[0];
  assign array_update_78533[1] = add_77421 == 32'h0000_0001 ? array_update_78531 : array_update_78520[1];
  assign array_update_78533[2] = add_77421 == 32'h0000_0002 ? array_update_78531 : array_update_78520[2];
  assign array_update_78533[3] = add_77421 == 32'h0000_0003 ? array_update_78531 : array_update_78520[3];
  assign array_update_78533[4] = add_77421 == 32'h0000_0004 ? array_update_78531 : array_update_78520[4];
  assign array_update_78533[5] = add_77421 == 32'h0000_0005 ? array_update_78531 : array_update_78520[5];
  assign array_update_78533[6] = add_77421 == 32'h0000_0006 ? array_update_78531 : array_update_78520[6];
  assign array_update_78533[7] = add_77421 == 32'h0000_0007 ? array_update_78531 : array_update_78520[7];
  assign array_update_78533[8] = add_77421 == 32'h0000_0008 ? array_update_78531 : array_update_78520[8];
  assign array_update_78533[9] = add_77421 == 32'h0000_0009 ? array_update_78531 : array_update_78520[9];
  assign array_index_78535 = array_update_72021[add_78532 > 32'h0000_0009 ? 4'h9 : add_78532[3:0]];
  assign array_index_78536 = array_update_78533[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_78540 = smul32b_32b_x_32b(array_index_77428[add_78532 > 32'h0000_0009 ? 4'h9 : add_78532[3:0]], array_index_78535[add_78504 > 32'h0000_0009 ? 4'h9 : add_78504[3:0]]);
  assign add_78542 = array_index_78536[add_78504 > 32'h0000_0009 ? 4'h9 : add_78504[3:0]] + smul_78540;
  assign array_update_78544[0] = add_78504 == 32'h0000_0000 ? add_78542 : array_index_78536[0];
  assign array_update_78544[1] = add_78504 == 32'h0000_0001 ? add_78542 : array_index_78536[1];
  assign array_update_78544[2] = add_78504 == 32'h0000_0002 ? add_78542 : array_index_78536[2];
  assign array_update_78544[3] = add_78504 == 32'h0000_0003 ? add_78542 : array_index_78536[3];
  assign array_update_78544[4] = add_78504 == 32'h0000_0004 ? add_78542 : array_index_78536[4];
  assign array_update_78544[5] = add_78504 == 32'h0000_0005 ? add_78542 : array_index_78536[5];
  assign array_update_78544[6] = add_78504 == 32'h0000_0006 ? add_78542 : array_index_78536[6];
  assign array_update_78544[7] = add_78504 == 32'h0000_0007 ? add_78542 : array_index_78536[7];
  assign array_update_78544[8] = add_78504 == 32'h0000_0008 ? add_78542 : array_index_78536[8];
  assign array_update_78544[9] = add_78504 == 32'h0000_0009 ? add_78542 : array_index_78536[9];
  assign add_78545 = add_78532 + 32'h0000_0001;
  assign array_update_78546[0] = add_77421 == 32'h0000_0000 ? array_update_78544 : array_update_78533[0];
  assign array_update_78546[1] = add_77421 == 32'h0000_0001 ? array_update_78544 : array_update_78533[1];
  assign array_update_78546[2] = add_77421 == 32'h0000_0002 ? array_update_78544 : array_update_78533[2];
  assign array_update_78546[3] = add_77421 == 32'h0000_0003 ? array_update_78544 : array_update_78533[3];
  assign array_update_78546[4] = add_77421 == 32'h0000_0004 ? array_update_78544 : array_update_78533[4];
  assign array_update_78546[5] = add_77421 == 32'h0000_0005 ? array_update_78544 : array_update_78533[5];
  assign array_update_78546[6] = add_77421 == 32'h0000_0006 ? array_update_78544 : array_update_78533[6];
  assign array_update_78546[7] = add_77421 == 32'h0000_0007 ? array_update_78544 : array_update_78533[7];
  assign array_update_78546[8] = add_77421 == 32'h0000_0008 ? array_update_78544 : array_update_78533[8];
  assign array_update_78546[9] = add_77421 == 32'h0000_0009 ? array_update_78544 : array_update_78533[9];
  assign array_index_78548 = array_update_72021[add_78545 > 32'h0000_0009 ? 4'h9 : add_78545[3:0]];
  assign array_index_78549 = array_update_78546[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_78553 = smul32b_32b_x_32b(array_index_77428[add_78545 > 32'h0000_0009 ? 4'h9 : add_78545[3:0]], array_index_78548[add_78504 > 32'h0000_0009 ? 4'h9 : add_78504[3:0]]);
  assign add_78555 = array_index_78549[add_78504 > 32'h0000_0009 ? 4'h9 : add_78504[3:0]] + smul_78553;
  assign array_update_78557[0] = add_78504 == 32'h0000_0000 ? add_78555 : array_index_78549[0];
  assign array_update_78557[1] = add_78504 == 32'h0000_0001 ? add_78555 : array_index_78549[1];
  assign array_update_78557[2] = add_78504 == 32'h0000_0002 ? add_78555 : array_index_78549[2];
  assign array_update_78557[3] = add_78504 == 32'h0000_0003 ? add_78555 : array_index_78549[3];
  assign array_update_78557[4] = add_78504 == 32'h0000_0004 ? add_78555 : array_index_78549[4];
  assign array_update_78557[5] = add_78504 == 32'h0000_0005 ? add_78555 : array_index_78549[5];
  assign array_update_78557[6] = add_78504 == 32'h0000_0006 ? add_78555 : array_index_78549[6];
  assign array_update_78557[7] = add_78504 == 32'h0000_0007 ? add_78555 : array_index_78549[7];
  assign array_update_78557[8] = add_78504 == 32'h0000_0008 ? add_78555 : array_index_78549[8];
  assign array_update_78557[9] = add_78504 == 32'h0000_0009 ? add_78555 : array_index_78549[9];
  assign add_78558 = add_78545 + 32'h0000_0001;
  assign array_update_78559[0] = add_77421 == 32'h0000_0000 ? array_update_78557 : array_update_78546[0];
  assign array_update_78559[1] = add_77421 == 32'h0000_0001 ? array_update_78557 : array_update_78546[1];
  assign array_update_78559[2] = add_77421 == 32'h0000_0002 ? array_update_78557 : array_update_78546[2];
  assign array_update_78559[3] = add_77421 == 32'h0000_0003 ? array_update_78557 : array_update_78546[3];
  assign array_update_78559[4] = add_77421 == 32'h0000_0004 ? array_update_78557 : array_update_78546[4];
  assign array_update_78559[5] = add_77421 == 32'h0000_0005 ? array_update_78557 : array_update_78546[5];
  assign array_update_78559[6] = add_77421 == 32'h0000_0006 ? array_update_78557 : array_update_78546[6];
  assign array_update_78559[7] = add_77421 == 32'h0000_0007 ? array_update_78557 : array_update_78546[7];
  assign array_update_78559[8] = add_77421 == 32'h0000_0008 ? array_update_78557 : array_update_78546[8];
  assign array_update_78559[9] = add_77421 == 32'h0000_0009 ? array_update_78557 : array_update_78546[9];
  assign array_index_78561 = array_update_72021[add_78558 > 32'h0000_0009 ? 4'h9 : add_78558[3:0]];
  assign array_index_78562 = array_update_78559[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_78566 = smul32b_32b_x_32b(array_index_77428[add_78558 > 32'h0000_0009 ? 4'h9 : add_78558[3:0]], array_index_78561[add_78504 > 32'h0000_0009 ? 4'h9 : add_78504[3:0]]);
  assign add_78568 = array_index_78562[add_78504 > 32'h0000_0009 ? 4'h9 : add_78504[3:0]] + smul_78566;
  assign array_update_78570[0] = add_78504 == 32'h0000_0000 ? add_78568 : array_index_78562[0];
  assign array_update_78570[1] = add_78504 == 32'h0000_0001 ? add_78568 : array_index_78562[1];
  assign array_update_78570[2] = add_78504 == 32'h0000_0002 ? add_78568 : array_index_78562[2];
  assign array_update_78570[3] = add_78504 == 32'h0000_0003 ? add_78568 : array_index_78562[3];
  assign array_update_78570[4] = add_78504 == 32'h0000_0004 ? add_78568 : array_index_78562[4];
  assign array_update_78570[5] = add_78504 == 32'h0000_0005 ? add_78568 : array_index_78562[5];
  assign array_update_78570[6] = add_78504 == 32'h0000_0006 ? add_78568 : array_index_78562[6];
  assign array_update_78570[7] = add_78504 == 32'h0000_0007 ? add_78568 : array_index_78562[7];
  assign array_update_78570[8] = add_78504 == 32'h0000_0008 ? add_78568 : array_index_78562[8];
  assign array_update_78570[9] = add_78504 == 32'h0000_0009 ? add_78568 : array_index_78562[9];
  assign add_78571 = add_78558 + 32'h0000_0001;
  assign array_update_78572[0] = add_77421 == 32'h0000_0000 ? array_update_78570 : array_update_78559[0];
  assign array_update_78572[1] = add_77421 == 32'h0000_0001 ? array_update_78570 : array_update_78559[1];
  assign array_update_78572[2] = add_77421 == 32'h0000_0002 ? array_update_78570 : array_update_78559[2];
  assign array_update_78572[3] = add_77421 == 32'h0000_0003 ? array_update_78570 : array_update_78559[3];
  assign array_update_78572[4] = add_77421 == 32'h0000_0004 ? array_update_78570 : array_update_78559[4];
  assign array_update_78572[5] = add_77421 == 32'h0000_0005 ? array_update_78570 : array_update_78559[5];
  assign array_update_78572[6] = add_77421 == 32'h0000_0006 ? array_update_78570 : array_update_78559[6];
  assign array_update_78572[7] = add_77421 == 32'h0000_0007 ? array_update_78570 : array_update_78559[7];
  assign array_update_78572[8] = add_77421 == 32'h0000_0008 ? array_update_78570 : array_update_78559[8];
  assign array_update_78572[9] = add_77421 == 32'h0000_0009 ? array_update_78570 : array_update_78559[9];
  assign array_index_78574 = array_update_72021[add_78571 > 32'h0000_0009 ? 4'h9 : add_78571[3:0]];
  assign array_index_78575 = array_update_78572[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_78579 = smul32b_32b_x_32b(array_index_77428[add_78571 > 32'h0000_0009 ? 4'h9 : add_78571[3:0]], array_index_78574[add_78504 > 32'h0000_0009 ? 4'h9 : add_78504[3:0]]);
  assign add_78581 = array_index_78575[add_78504 > 32'h0000_0009 ? 4'h9 : add_78504[3:0]] + smul_78579;
  assign array_update_78583[0] = add_78504 == 32'h0000_0000 ? add_78581 : array_index_78575[0];
  assign array_update_78583[1] = add_78504 == 32'h0000_0001 ? add_78581 : array_index_78575[1];
  assign array_update_78583[2] = add_78504 == 32'h0000_0002 ? add_78581 : array_index_78575[2];
  assign array_update_78583[3] = add_78504 == 32'h0000_0003 ? add_78581 : array_index_78575[3];
  assign array_update_78583[4] = add_78504 == 32'h0000_0004 ? add_78581 : array_index_78575[4];
  assign array_update_78583[5] = add_78504 == 32'h0000_0005 ? add_78581 : array_index_78575[5];
  assign array_update_78583[6] = add_78504 == 32'h0000_0006 ? add_78581 : array_index_78575[6];
  assign array_update_78583[7] = add_78504 == 32'h0000_0007 ? add_78581 : array_index_78575[7];
  assign array_update_78583[8] = add_78504 == 32'h0000_0008 ? add_78581 : array_index_78575[8];
  assign array_update_78583[9] = add_78504 == 32'h0000_0009 ? add_78581 : array_index_78575[9];
  assign add_78584 = add_78571 + 32'h0000_0001;
  assign array_update_78585[0] = add_77421 == 32'h0000_0000 ? array_update_78583 : array_update_78572[0];
  assign array_update_78585[1] = add_77421 == 32'h0000_0001 ? array_update_78583 : array_update_78572[1];
  assign array_update_78585[2] = add_77421 == 32'h0000_0002 ? array_update_78583 : array_update_78572[2];
  assign array_update_78585[3] = add_77421 == 32'h0000_0003 ? array_update_78583 : array_update_78572[3];
  assign array_update_78585[4] = add_77421 == 32'h0000_0004 ? array_update_78583 : array_update_78572[4];
  assign array_update_78585[5] = add_77421 == 32'h0000_0005 ? array_update_78583 : array_update_78572[5];
  assign array_update_78585[6] = add_77421 == 32'h0000_0006 ? array_update_78583 : array_update_78572[6];
  assign array_update_78585[7] = add_77421 == 32'h0000_0007 ? array_update_78583 : array_update_78572[7];
  assign array_update_78585[8] = add_77421 == 32'h0000_0008 ? array_update_78583 : array_update_78572[8];
  assign array_update_78585[9] = add_77421 == 32'h0000_0009 ? array_update_78583 : array_update_78572[9];
  assign array_index_78587 = array_update_72021[add_78584 > 32'h0000_0009 ? 4'h9 : add_78584[3:0]];
  assign array_index_78588 = array_update_78585[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_78592 = smul32b_32b_x_32b(array_index_77428[add_78584 > 32'h0000_0009 ? 4'h9 : add_78584[3:0]], array_index_78587[add_78504 > 32'h0000_0009 ? 4'h9 : add_78504[3:0]]);
  assign add_78594 = array_index_78588[add_78504 > 32'h0000_0009 ? 4'h9 : add_78504[3:0]] + smul_78592;
  assign array_update_78596[0] = add_78504 == 32'h0000_0000 ? add_78594 : array_index_78588[0];
  assign array_update_78596[1] = add_78504 == 32'h0000_0001 ? add_78594 : array_index_78588[1];
  assign array_update_78596[2] = add_78504 == 32'h0000_0002 ? add_78594 : array_index_78588[2];
  assign array_update_78596[3] = add_78504 == 32'h0000_0003 ? add_78594 : array_index_78588[3];
  assign array_update_78596[4] = add_78504 == 32'h0000_0004 ? add_78594 : array_index_78588[4];
  assign array_update_78596[5] = add_78504 == 32'h0000_0005 ? add_78594 : array_index_78588[5];
  assign array_update_78596[6] = add_78504 == 32'h0000_0006 ? add_78594 : array_index_78588[6];
  assign array_update_78596[7] = add_78504 == 32'h0000_0007 ? add_78594 : array_index_78588[7];
  assign array_update_78596[8] = add_78504 == 32'h0000_0008 ? add_78594 : array_index_78588[8];
  assign array_update_78596[9] = add_78504 == 32'h0000_0009 ? add_78594 : array_index_78588[9];
  assign add_78597 = add_78584 + 32'h0000_0001;
  assign array_update_78598[0] = add_77421 == 32'h0000_0000 ? array_update_78596 : array_update_78585[0];
  assign array_update_78598[1] = add_77421 == 32'h0000_0001 ? array_update_78596 : array_update_78585[1];
  assign array_update_78598[2] = add_77421 == 32'h0000_0002 ? array_update_78596 : array_update_78585[2];
  assign array_update_78598[3] = add_77421 == 32'h0000_0003 ? array_update_78596 : array_update_78585[3];
  assign array_update_78598[4] = add_77421 == 32'h0000_0004 ? array_update_78596 : array_update_78585[4];
  assign array_update_78598[5] = add_77421 == 32'h0000_0005 ? array_update_78596 : array_update_78585[5];
  assign array_update_78598[6] = add_77421 == 32'h0000_0006 ? array_update_78596 : array_update_78585[6];
  assign array_update_78598[7] = add_77421 == 32'h0000_0007 ? array_update_78596 : array_update_78585[7];
  assign array_update_78598[8] = add_77421 == 32'h0000_0008 ? array_update_78596 : array_update_78585[8];
  assign array_update_78598[9] = add_77421 == 32'h0000_0009 ? array_update_78596 : array_update_78585[9];
  assign array_index_78600 = array_update_72021[add_78597 > 32'h0000_0009 ? 4'h9 : add_78597[3:0]];
  assign array_index_78601 = array_update_78598[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_78605 = smul32b_32b_x_32b(array_index_77428[add_78597 > 32'h0000_0009 ? 4'h9 : add_78597[3:0]], array_index_78600[add_78504 > 32'h0000_0009 ? 4'h9 : add_78504[3:0]]);
  assign add_78607 = array_index_78601[add_78504 > 32'h0000_0009 ? 4'h9 : add_78504[3:0]] + smul_78605;
  assign array_update_78609[0] = add_78504 == 32'h0000_0000 ? add_78607 : array_index_78601[0];
  assign array_update_78609[1] = add_78504 == 32'h0000_0001 ? add_78607 : array_index_78601[1];
  assign array_update_78609[2] = add_78504 == 32'h0000_0002 ? add_78607 : array_index_78601[2];
  assign array_update_78609[3] = add_78504 == 32'h0000_0003 ? add_78607 : array_index_78601[3];
  assign array_update_78609[4] = add_78504 == 32'h0000_0004 ? add_78607 : array_index_78601[4];
  assign array_update_78609[5] = add_78504 == 32'h0000_0005 ? add_78607 : array_index_78601[5];
  assign array_update_78609[6] = add_78504 == 32'h0000_0006 ? add_78607 : array_index_78601[6];
  assign array_update_78609[7] = add_78504 == 32'h0000_0007 ? add_78607 : array_index_78601[7];
  assign array_update_78609[8] = add_78504 == 32'h0000_0008 ? add_78607 : array_index_78601[8];
  assign array_update_78609[9] = add_78504 == 32'h0000_0009 ? add_78607 : array_index_78601[9];
  assign add_78610 = add_78597 + 32'h0000_0001;
  assign array_update_78611[0] = add_77421 == 32'h0000_0000 ? array_update_78609 : array_update_78598[0];
  assign array_update_78611[1] = add_77421 == 32'h0000_0001 ? array_update_78609 : array_update_78598[1];
  assign array_update_78611[2] = add_77421 == 32'h0000_0002 ? array_update_78609 : array_update_78598[2];
  assign array_update_78611[3] = add_77421 == 32'h0000_0003 ? array_update_78609 : array_update_78598[3];
  assign array_update_78611[4] = add_77421 == 32'h0000_0004 ? array_update_78609 : array_update_78598[4];
  assign array_update_78611[5] = add_77421 == 32'h0000_0005 ? array_update_78609 : array_update_78598[5];
  assign array_update_78611[6] = add_77421 == 32'h0000_0006 ? array_update_78609 : array_update_78598[6];
  assign array_update_78611[7] = add_77421 == 32'h0000_0007 ? array_update_78609 : array_update_78598[7];
  assign array_update_78611[8] = add_77421 == 32'h0000_0008 ? array_update_78609 : array_update_78598[8];
  assign array_update_78611[9] = add_77421 == 32'h0000_0009 ? array_update_78609 : array_update_78598[9];
  assign array_index_78613 = array_update_72021[add_78610 > 32'h0000_0009 ? 4'h9 : add_78610[3:0]];
  assign array_index_78614 = array_update_78611[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_78618 = smul32b_32b_x_32b(array_index_77428[add_78610 > 32'h0000_0009 ? 4'h9 : add_78610[3:0]], array_index_78613[add_78504 > 32'h0000_0009 ? 4'h9 : add_78504[3:0]]);
  assign add_78620 = array_index_78614[add_78504 > 32'h0000_0009 ? 4'h9 : add_78504[3:0]] + smul_78618;
  assign array_update_78622[0] = add_78504 == 32'h0000_0000 ? add_78620 : array_index_78614[0];
  assign array_update_78622[1] = add_78504 == 32'h0000_0001 ? add_78620 : array_index_78614[1];
  assign array_update_78622[2] = add_78504 == 32'h0000_0002 ? add_78620 : array_index_78614[2];
  assign array_update_78622[3] = add_78504 == 32'h0000_0003 ? add_78620 : array_index_78614[3];
  assign array_update_78622[4] = add_78504 == 32'h0000_0004 ? add_78620 : array_index_78614[4];
  assign array_update_78622[5] = add_78504 == 32'h0000_0005 ? add_78620 : array_index_78614[5];
  assign array_update_78622[6] = add_78504 == 32'h0000_0006 ? add_78620 : array_index_78614[6];
  assign array_update_78622[7] = add_78504 == 32'h0000_0007 ? add_78620 : array_index_78614[7];
  assign array_update_78622[8] = add_78504 == 32'h0000_0008 ? add_78620 : array_index_78614[8];
  assign array_update_78622[9] = add_78504 == 32'h0000_0009 ? add_78620 : array_index_78614[9];
  assign add_78623 = add_78610 + 32'h0000_0001;
  assign array_update_78624[0] = add_77421 == 32'h0000_0000 ? array_update_78622 : array_update_78611[0];
  assign array_update_78624[1] = add_77421 == 32'h0000_0001 ? array_update_78622 : array_update_78611[1];
  assign array_update_78624[2] = add_77421 == 32'h0000_0002 ? array_update_78622 : array_update_78611[2];
  assign array_update_78624[3] = add_77421 == 32'h0000_0003 ? array_update_78622 : array_update_78611[3];
  assign array_update_78624[4] = add_77421 == 32'h0000_0004 ? array_update_78622 : array_update_78611[4];
  assign array_update_78624[5] = add_77421 == 32'h0000_0005 ? array_update_78622 : array_update_78611[5];
  assign array_update_78624[6] = add_77421 == 32'h0000_0006 ? array_update_78622 : array_update_78611[6];
  assign array_update_78624[7] = add_77421 == 32'h0000_0007 ? array_update_78622 : array_update_78611[7];
  assign array_update_78624[8] = add_77421 == 32'h0000_0008 ? array_update_78622 : array_update_78611[8];
  assign array_update_78624[9] = add_77421 == 32'h0000_0009 ? array_update_78622 : array_update_78611[9];
  assign array_index_78626 = array_update_72021[add_78623 > 32'h0000_0009 ? 4'h9 : add_78623[3:0]];
  assign array_index_78627 = array_update_78624[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_78631 = smul32b_32b_x_32b(array_index_77428[add_78623 > 32'h0000_0009 ? 4'h9 : add_78623[3:0]], array_index_78626[add_78504 > 32'h0000_0009 ? 4'h9 : add_78504[3:0]]);
  assign add_78633 = array_index_78627[add_78504 > 32'h0000_0009 ? 4'h9 : add_78504[3:0]] + smul_78631;
  assign array_update_78634[0] = add_78504 == 32'h0000_0000 ? add_78633 : array_index_78627[0];
  assign array_update_78634[1] = add_78504 == 32'h0000_0001 ? add_78633 : array_index_78627[1];
  assign array_update_78634[2] = add_78504 == 32'h0000_0002 ? add_78633 : array_index_78627[2];
  assign array_update_78634[3] = add_78504 == 32'h0000_0003 ? add_78633 : array_index_78627[3];
  assign array_update_78634[4] = add_78504 == 32'h0000_0004 ? add_78633 : array_index_78627[4];
  assign array_update_78634[5] = add_78504 == 32'h0000_0005 ? add_78633 : array_index_78627[5];
  assign array_update_78634[6] = add_78504 == 32'h0000_0006 ? add_78633 : array_index_78627[6];
  assign array_update_78634[7] = add_78504 == 32'h0000_0007 ? add_78633 : array_index_78627[7];
  assign array_update_78634[8] = add_78504 == 32'h0000_0008 ? add_78633 : array_index_78627[8];
  assign array_update_78634[9] = add_78504 == 32'h0000_0009 ? add_78633 : array_index_78627[9];
  assign array_update_78635[0] = add_77421 == 32'h0000_0000 ? array_update_78634 : array_update_78624[0];
  assign array_update_78635[1] = add_77421 == 32'h0000_0001 ? array_update_78634 : array_update_78624[1];
  assign array_update_78635[2] = add_77421 == 32'h0000_0002 ? array_update_78634 : array_update_78624[2];
  assign array_update_78635[3] = add_77421 == 32'h0000_0003 ? array_update_78634 : array_update_78624[3];
  assign array_update_78635[4] = add_77421 == 32'h0000_0004 ? array_update_78634 : array_update_78624[4];
  assign array_update_78635[5] = add_77421 == 32'h0000_0005 ? array_update_78634 : array_update_78624[5];
  assign array_update_78635[6] = add_77421 == 32'h0000_0006 ? array_update_78634 : array_update_78624[6];
  assign array_update_78635[7] = add_77421 == 32'h0000_0007 ? array_update_78634 : array_update_78624[7];
  assign array_update_78635[8] = add_77421 == 32'h0000_0008 ? array_update_78634 : array_update_78624[8];
  assign array_update_78635[9] = add_77421 == 32'h0000_0009 ? array_update_78634 : array_update_78624[9];
  assign array_index_78637 = array_update_78635[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign add_78639 = add_78504 + 32'h0000_0001;
  assign array_update_78640[0] = add_78639 == 32'h0000_0000 ? 32'h0000_0000 : array_index_78637[0];
  assign array_update_78640[1] = add_78639 == 32'h0000_0001 ? 32'h0000_0000 : array_index_78637[1];
  assign array_update_78640[2] = add_78639 == 32'h0000_0002 ? 32'h0000_0000 : array_index_78637[2];
  assign array_update_78640[3] = add_78639 == 32'h0000_0003 ? 32'h0000_0000 : array_index_78637[3];
  assign array_update_78640[4] = add_78639 == 32'h0000_0004 ? 32'h0000_0000 : array_index_78637[4];
  assign array_update_78640[5] = add_78639 == 32'h0000_0005 ? 32'h0000_0000 : array_index_78637[5];
  assign array_update_78640[6] = add_78639 == 32'h0000_0006 ? 32'h0000_0000 : array_index_78637[6];
  assign array_update_78640[7] = add_78639 == 32'h0000_0007 ? 32'h0000_0000 : array_index_78637[7];
  assign array_update_78640[8] = add_78639 == 32'h0000_0008 ? 32'h0000_0000 : array_index_78637[8];
  assign array_update_78640[9] = add_78639 == 32'h0000_0009 ? 32'h0000_0000 : array_index_78637[9];
  assign literal_78641 = 32'h0000_0000;
  assign array_update_78642[0] = add_77421 == 32'h0000_0000 ? array_update_78640 : array_update_78635[0];
  assign array_update_78642[1] = add_77421 == 32'h0000_0001 ? array_update_78640 : array_update_78635[1];
  assign array_update_78642[2] = add_77421 == 32'h0000_0002 ? array_update_78640 : array_update_78635[2];
  assign array_update_78642[3] = add_77421 == 32'h0000_0003 ? array_update_78640 : array_update_78635[3];
  assign array_update_78642[4] = add_77421 == 32'h0000_0004 ? array_update_78640 : array_update_78635[4];
  assign array_update_78642[5] = add_77421 == 32'h0000_0005 ? array_update_78640 : array_update_78635[5];
  assign array_update_78642[6] = add_77421 == 32'h0000_0006 ? array_update_78640 : array_update_78635[6];
  assign array_update_78642[7] = add_77421 == 32'h0000_0007 ? array_update_78640 : array_update_78635[7];
  assign array_update_78642[8] = add_77421 == 32'h0000_0008 ? array_update_78640 : array_update_78635[8];
  assign array_update_78642[9] = add_77421 == 32'h0000_0009 ? array_update_78640 : array_update_78635[9];
  assign array_index_78644 = array_update_72021[literal_78641 > 32'h0000_0009 ? 4'h9 : literal_78641[3:0]];
  assign array_index_78645 = array_update_78642[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_78649 = smul32b_32b_x_32b(array_index_77428[literal_78641 > 32'h0000_0009 ? 4'h9 : literal_78641[3:0]], array_index_78644[add_78639 > 32'h0000_0009 ? 4'h9 : add_78639[3:0]]);
  assign add_78651 = array_index_78645[add_78639 > 32'h0000_0009 ? 4'h9 : add_78639[3:0]] + smul_78649;
  assign array_update_78653[0] = add_78639 == 32'h0000_0000 ? add_78651 : array_index_78645[0];
  assign array_update_78653[1] = add_78639 == 32'h0000_0001 ? add_78651 : array_index_78645[1];
  assign array_update_78653[2] = add_78639 == 32'h0000_0002 ? add_78651 : array_index_78645[2];
  assign array_update_78653[3] = add_78639 == 32'h0000_0003 ? add_78651 : array_index_78645[3];
  assign array_update_78653[4] = add_78639 == 32'h0000_0004 ? add_78651 : array_index_78645[4];
  assign array_update_78653[5] = add_78639 == 32'h0000_0005 ? add_78651 : array_index_78645[5];
  assign array_update_78653[6] = add_78639 == 32'h0000_0006 ? add_78651 : array_index_78645[6];
  assign array_update_78653[7] = add_78639 == 32'h0000_0007 ? add_78651 : array_index_78645[7];
  assign array_update_78653[8] = add_78639 == 32'h0000_0008 ? add_78651 : array_index_78645[8];
  assign array_update_78653[9] = add_78639 == 32'h0000_0009 ? add_78651 : array_index_78645[9];
  assign add_78654 = literal_78641 + 32'h0000_0001;
  assign array_update_78655[0] = add_77421 == 32'h0000_0000 ? array_update_78653 : array_update_78642[0];
  assign array_update_78655[1] = add_77421 == 32'h0000_0001 ? array_update_78653 : array_update_78642[1];
  assign array_update_78655[2] = add_77421 == 32'h0000_0002 ? array_update_78653 : array_update_78642[2];
  assign array_update_78655[3] = add_77421 == 32'h0000_0003 ? array_update_78653 : array_update_78642[3];
  assign array_update_78655[4] = add_77421 == 32'h0000_0004 ? array_update_78653 : array_update_78642[4];
  assign array_update_78655[5] = add_77421 == 32'h0000_0005 ? array_update_78653 : array_update_78642[5];
  assign array_update_78655[6] = add_77421 == 32'h0000_0006 ? array_update_78653 : array_update_78642[6];
  assign array_update_78655[7] = add_77421 == 32'h0000_0007 ? array_update_78653 : array_update_78642[7];
  assign array_update_78655[8] = add_77421 == 32'h0000_0008 ? array_update_78653 : array_update_78642[8];
  assign array_update_78655[9] = add_77421 == 32'h0000_0009 ? array_update_78653 : array_update_78642[9];
  assign array_index_78657 = array_update_72021[add_78654 > 32'h0000_0009 ? 4'h9 : add_78654[3:0]];
  assign array_index_78658 = array_update_78655[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_78662 = smul32b_32b_x_32b(array_index_77428[add_78654 > 32'h0000_0009 ? 4'h9 : add_78654[3:0]], array_index_78657[add_78639 > 32'h0000_0009 ? 4'h9 : add_78639[3:0]]);
  assign add_78664 = array_index_78658[add_78639 > 32'h0000_0009 ? 4'h9 : add_78639[3:0]] + smul_78662;
  assign array_update_78666[0] = add_78639 == 32'h0000_0000 ? add_78664 : array_index_78658[0];
  assign array_update_78666[1] = add_78639 == 32'h0000_0001 ? add_78664 : array_index_78658[1];
  assign array_update_78666[2] = add_78639 == 32'h0000_0002 ? add_78664 : array_index_78658[2];
  assign array_update_78666[3] = add_78639 == 32'h0000_0003 ? add_78664 : array_index_78658[3];
  assign array_update_78666[4] = add_78639 == 32'h0000_0004 ? add_78664 : array_index_78658[4];
  assign array_update_78666[5] = add_78639 == 32'h0000_0005 ? add_78664 : array_index_78658[5];
  assign array_update_78666[6] = add_78639 == 32'h0000_0006 ? add_78664 : array_index_78658[6];
  assign array_update_78666[7] = add_78639 == 32'h0000_0007 ? add_78664 : array_index_78658[7];
  assign array_update_78666[8] = add_78639 == 32'h0000_0008 ? add_78664 : array_index_78658[8];
  assign array_update_78666[9] = add_78639 == 32'h0000_0009 ? add_78664 : array_index_78658[9];
  assign add_78667 = add_78654 + 32'h0000_0001;
  assign array_update_78668[0] = add_77421 == 32'h0000_0000 ? array_update_78666 : array_update_78655[0];
  assign array_update_78668[1] = add_77421 == 32'h0000_0001 ? array_update_78666 : array_update_78655[1];
  assign array_update_78668[2] = add_77421 == 32'h0000_0002 ? array_update_78666 : array_update_78655[2];
  assign array_update_78668[3] = add_77421 == 32'h0000_0003 ? array_update_78666 : array_update_78655[3];
  assign array_update_78668[4] = add_77421 == 32'h0000_0004 ? array_update_78666 : array_update_78655[4];
  assign array_update_78668[5] = add_77421 == 32'h0000_0005 ? array_update_78666 : array_update_78655[5];
  assign array_update_78668[6] = add_77421 == 32'h0000_0006 ? array_update_78666 : array_update_78655[6];
  assign array_update_78668[7] = add_77421 == 32'h0000_0007 ? array_update_78666 : array_update_78655[7];
  assign array_update_78668[8] = add_77421 == 32'h0000_0008 ? array_update_78666 : array_update_78655[8];
  assign array_update_78668[9] = add_77421 == 32'h0000_0009 ? array_update_78666 : array_update_78655[9];
  assign array_index_78670 = array_update_72021[add_78667 > 32'h0000_0009 ? 4'h9 : add_78667[3:0]];
  assign array_index_78671 = array_update_78668[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_78675 = smul32b_32b_x_32b(array_index_77428[add_78667 > 32'h0000_0009 ? 4'h9 : add_78667[3:0]], array_index_78670[add_78639 > 32'h0000_0009 ? 4'h9 : add_78639[3:0]]);
  assign add_78677 = array_index_78671[add_78639 > 32'h0000_0009 ? 4'h9 : add_78639[3:0]] + smul_78675;
  assign array_update_78679[0] = add_78639 == 32'h0000_0000 ? add_78677 : array_index_78671[0];
  assign array_update_78679[1] = add_78639 == 32'h0000_0001 ? add_78677 : array_index_78671[1];
  assign array_update_78679[2] = add_78639 == 32'h0000_0002 ? add_78677 : array_index_78671[2];
  assign array_update_78679[3] = add_78639 == 32'h0000_0003 ? add_78677 : array_index_78671[3];
  assign array_update_78679[4] = add_78639 == 32'h0000_0004 ? add_78677 : array_index_78671[4];
  assign array_update_78679[5] = add_78639 == 32'h0000_0005 ? add_78677 : array_index_78671[5];
  assign array_update_78679[6] = add_78639 == 32'h0000_0006 ? add_78677 : array_index_78671[6];
  assign array_update_78679[7] = add_78639 == 32'h0000_0007 ? add_78677 : array_index_78671[7];
  assign array_update_78679[8] = add_78639 == 32'h0000_0008 ? add_78677 : array_index_78671[8];
  assign array_update_78679[9] = add_78639 == 32'h0000_0009 ? add_78677 : array_index_78671[9];
  assign add_78680 = add_78667 + 32'h0000_0001;
  assign array_update_78681[0] = add_77421 == 32'h0000_0000 ? array_update_78679 : array_update_78668[0];
  assign array_update_78681[1] = add_77421 == 32'h0000_0001 ? array_update_78679 : array_update_78668[1];
  assign array_update_78681[2] = add_77421 == 32'h0000_0002 ? array_update_78679 : array_update_78668[2];
  assign array_update_78681[3] = add_77421 == 32'h0000_0003 ? array_update_78679 : array_update_78668[3];
  assign array_update_78681[4] = add_77421 == 32'h0000_0004 ? array_update_78679 : array_update_78668[4];
  assign array_update_78681[5] = add_77421 == 32'h0000_0005 ? array_update_78679 : array_update_78668[5];
  assign array_update_78681[6] = add_77421 == 32'h0000_0006 ? array_update_78679 : array_update_78668[6];
  assign array_update_78681[7] = add_77421 == 32'h0000_0007 ? array_update_78679 : array_update_78668[7];
  assign array_update_78681[8] = add_77421 == 32'h0000_0008 ? array_update_78679 : array_update_78668[8];
  assign array_update_78681[9] = add_77421 == 32'h0000_0009 ? array_update_78679 : array_update_78668[9];
  assign array_index_78683 = array_update_72021[add_78680 > 32'h0000_0009 ? 4'h9 : add_78680[3:0]];
  assign array_index_78684 = array_update_78681[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_78688 = smul32b_32b_x_32b(array_index_77428[add_78680 > 32'h0000_0009 ? 4'h9 : add_78680[3:0]], array_index_78683[add_78639 > 32'h0000_0009 ? 4'h9 : add_78639[3:0]]);
  assign add_78690 = array_index_78684[add_78639 > 32'h0000_0009 ? 4'h9 : add_78639[3:0]] + smul_78688;
  assign array_update_78692[0] = add_78639 == 32'h0000_0000 ? add_78690 : array_index_78684[0];
  assign array_update_78692[1] = add_78639 == 32'h0000_0001 ? add_78690 : array_index_78684[1];
  assign array_update_78692[2] = add_78639 == 32'h0000_0002 ? add_78690 : array_index_78684[2];
  assign array_update_78692[3] = add_78639 == 32'h0000_0003 ? add_78690 : array_index_78684[3];
  assign array_update_78692[4] = add_78639 == 32'h0000_0004 ? add_78690 : array_index_78684[4];
  assign array_update_78692[5] = add_78639 == 32'h0000_0005 ? add_78690 : array_index_78684[5];
  assign array_update_78692[6] = add_78639 == 32'h0000_0006 ? add_78690 : array_index_78684[6];
  assign array_update_78692[7] = add_78639 == 32'h0000_0007 ? add_78690 : array_index_78684[7];
  assign array_update_78692[8] = add_78639 == 32'h0000_0008 ? add_78690 : array_index_78684[8];
  assign array_update_78692[9] = add_78639 == 32'h0000_0009 ? add_78690 : array_index_78684[9];
  assign add_78693 = add_78680 + 32'h0000_0001;
  assign array_update_78694[0] = add_77421 == 32'h0000_0000 ? array_update_78692 : array_update_78681[0];
  assign array_update_78694[1] = add_77421 == 32'h0000_0001 ? array_update_78692 : array_update_78681[1];
  assign array_update_78694[2] = add_77421 == 32'h0000_0002 ? array_update_78692 : array_update_78681[2];
  assign array_update_78694[3] = add_77421 == 32'h0000_0003 ? array_update_78692 : array_update_78681[3];
  assign array_update_78694[4] = add_77421 == 32'h0000_0004 ? array_update_78692 : array_update_78681[4];
  assign array_update_78694[5] = add_77421 == 32'h0000_0005 ? array_update_78692 : array_update_78681[5];
  assign array_update_78694[6] = add_77421 == 32'h0000_0006 ? array_update_78692 : array_update_78681[6];
  assign array_update_78694[7] = add_77421 == 32'h0000_0007 ? array_update_78692 : array_update_78681[7];
  assign array_update_78694[8] = add_77421 == 32'h0000_0008 ? array_update_78692 : array_update_78681[8];
  assign array_update_78694[9] = add_77421 == 32'h0000_0009 ? array_update_78692 : array_update_78681[9];
  assign array_index_78696 = array_update_72021[add_78693 > 32'h0000_0009 ? 4'h9 : add_78693[3:0]];
  assign array_index_78697 = array_update_78694[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_78701 = smul32b_32b_x_32b(array_index_77428[add_78693 > 32'h0000_0009 ? 4'h9 : add_78693[3:0]], array_index_78696[add_78639 > 32'h0000_0009 ? 4'h9 : add_78639[3:0]]);
  assign add_78703 = array_index_78697[add_78639 > 32'h0000_0009 ? 4'h9 : add_78639[3:0]] + smul_78701;
  assign array_update_78705[0] = add_78639 == 32'h0000_0000 ? add_78703 : array_index_78697[0];
  assign array_update_78705[1] = add_78639 == 32'h0000_0001 ? add_78703 : array_index_78697[1];
  assign array_update_78705[2] = add_78639 == 32'h0000_0002 ? add_78703 : array_index_78697[2];
  assign array_update_78705[3] = add_78639 == 32'h0000_0003 ? add_78703 : array_index_78697[3];
  assign array_update_78705[4] = add_78639 == 32'h0000_0004 ? add_78703 : array_index_78697[4];
  assign array_update_78705[5] = add_78639 == 32'h0000_0005 ? add_78703 : array_index_78697[5];
  assign array_update_78705[6] = add_78639 == 32'h0000_0006 ? add_78703 : array_index_78697[6];
  assign array_update_78705[7] = add_78639 == 32'h0000_0007 ? add_78703 : array_index_78697[7];
  assign array_update_78705[8] = add_78639 == 32'h0000_0008 ? add_78703 : array_index_78697[8];
  assign array_update_78705[9] = add_78639 == 32'h0000_0009 ? add_78703 : array_index_78697[9];
  assign add_78706 = add_78693 + 32'h0000_0001;
  assign array_update_78707[0] = add_77421 == 32'h0000_0000 ? array_update_78705 : array_update_78694[0];
  assign array_update_78707[1] = add_77421 == 32'h0000_0001 ? array_update_78705 : array_update_78694[1];
  assign array_update_78707[2] = add_77421 == 32'h0000_0002 ? array_update_78705 : array_update_78694[2];
  assign array_update_78707[3] = add_77421 == 32'h0000_0003 ? array_update_78705 : array_update_78694[3];
  assign array_update_78707[4] = add_77421 == 32'h0000_0004 ? array_update_78705 : array_update_78694[4];
  assign array_update_78707[5] = add_77421 == 32'h0000_0005 ? array_update_78705 : array_update_78694[5];
  assign array_update_78707[6] = add_77421 == 32'h0000_0006 ? array_update_78705 : array_update_78694[6];
  assign array_update_78707[7] = add_77421 == 32'h0000_0007 ? array_update_78705 : array_update_78694[7];
  assign array_update_78707[8] = add_77421 == 32'h0000_0008 ? array_update_78705 : array_update_78694[8];
  assign array_update_78707[9] = add_77421 == 32'h0000_0009 ? array_update_78705 : array_update_78694[9];
  assign array_index_78709 = array_update_72021[add_78706 > 32'h0000_0009 ? 4'h9 : add_78706[3:0]];
  assign array_index_78710 = array_update_78707[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_78714 = smul32b_32b_x_32b(array_index_77428[add_78706 > 32'h0000_0009 ? 4'h9 : add_78706[3:0]], array_index_78709[add_78639 > 32'h0000_0009 ? 4'h9 : add_78639[3:0]]);
  assign add_78716 = array_index_78710[add_78639 > 32'h0000_0009 ? 4'h9 : add_78639[3:0]] + smul_78714;
  assign array_update_78718[0] = add_78639 == 32'h0000_0000 ? add_78716 : array_index_78710[0];
  assign array_update_78718[1] = add_78639 == 32'h0000_0001 ? add_78716 : array_index_78710[1];
  assign array_update_78718[2] = add_78639 == 32'h0000_0002 ? add_78716 : array_index_78710[2];
  assign array_update_78718[3] = add_78639 == 32'h0000_0003 ? add_78716 : array_index_78710[3];
  assign array_update_78718[4] = add_78639 == 32'h0000_0004 ? add_78716 : array_index_78710[4];
  assign array_update_78718[5] = add_78639 == 32'h0000_0005 ? add_78716 : array_index_78710[5];
  assign array_update_78718[6] = add_78639 == 32'h0000_0006 ? add_78716 : array_index_78710[6];
  assign array_update_78718[7] = add_78639 == 32'h0000_0007 ? add_78716 : array_index_78710[7];
  assign array_update_78718[8] = add_78639 == 32'h0000_0008 ? add_78716 : array_index_78710[8];
  assign array_update_78718[9] = add_78639 == 32'h0000_0009 ? add_78716 : array_index_78710[9];
  assign add_78719 = add_78706 + 32'h0000_0001;
  assign array_update_78720[0] = add_77421 == 32'h0000_0000 ? array_update_78718 : array_update_78707[0];
  assign array_update_78720[1] = add_77421 == 32'h0000_0001 ? array_update_78718 : array_update_78707[1];
  assign array_update_78720[2] = add_77421 == 32'h0000_0002 ? array_update_78718 : array_update_78707[2];
  assign array_update_78720[3] = add_77421 == 32'h0000_0003 ? array_update_78718 : array_update_78707[3];
  assign array_update_78720[4] = add_77421 == 32'h0000_0004 ? array_update_78718 : array_update_78707[4];
  assign array_update_78720[5] = add_77421 == 32'h0000_0005 ? array_update_78718 : array_update_78707[5];
  assign array_update_78720[6] = add_77421 == 32'h0000_0006 ? array_update_78718 : array_update_78707[6];
  assign array_update_78720[7] = add_77421 == 32'h0000_0007 ? array_update_78718 : array_update_78707[7];
  assign array_update_78720[8] = add_77421 == 32'h0000_0008 ? array_update_78718 : array_update_78707[8];
  assign array_update_78720[9] = add_77421 == 32'h0000_0009 ? array_update_78718 : array_update_78707[9];
  assign array_index_78722 = array_update_72021[add_78719 > 32'h0000_0009 ? 4'h9 : add_78719[3:0]];
  assign array_index_78723 = array_update_78720[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_78727 = smul32b_32b_x_32b(array_index_77428[add_78719 > 32'h0000_0009 ? 4'h9 : add_78719[3:0]], array_index_78722[add_78639 > 32'h0000_0009 ? 4'h9 : add_78639[3:0]]);
  assign add_78729 = array_index_78723[add_78639 > 32'h0000_0009 ? 4'h9 : add_78639[3:0]] + smul_78727;
  assign array_update_78731[0] = add_78639 == 32'h0000_0000 ? add_78729 : array_index_78723[0];
  assign array_update_78731[1] = add_78639 == 32'h0000_0001 ? add_78729 : array_index_78723[1];
  assign array_update_78731[2] = add_78639 == 32'h0000_0002 ? add_78729 : array_index_78723[2];
  assign array_update_78731[3] = add_78639 == 32'h0000_0003 ? add_78729 : array_index_78723[3];
  assign array_update_78731[4] = add_78639 == 32'h0000_0004 ? add_78729 : array_index_78723[4];
  assign array_update_78731[5] = add_78639 == 32'h0000_0005 ? add_78729 : array_index_78723[5];
  assign array_update_78731[6] = add_78639 == 32'h0000_0006 ? add_78729 : array_index_78723[6];
  assign array_update_78731[7] = add_78639 == 32'h0000_0007 ? add_78729 : array_index_78723[7];
  assign array_update_78731[8] = add_78639 == 32'h0000_0008 ? add_78729 : array_index_78723[8];
  assign array_update_78731[9] = add_78639 == 32'h0000_0009 ? add_78729 : array_index_78723[9];
  assign add_78732 = add_78719 + 32'h0000_0001;
  assign array_update_78733[0] = add_77421 == 32'h0000_0000 ? array_update_78731 : array_update_78720[0];
  assign array_update_78733[1] = add_77421 == 32'h0000_0001 ? array_update_78731 : array_update_78720[1];
  assign array_update_78733[2] = add_77421 == 32'h0000_0002 ? array_update_78731 : array_update_78720[2];
  assign array_update_78733[3] = add_77421 == 32'h0000_0003 ? array_update_78731 : array_update_78720[3];
  assign array_update_78733[4] = add_77421 == 32'h0000_0004 ? array_update_78731 : array_update_78720[4];
  assign array_update_78733[5] = add_77421 == 32'h0000_0005 ? array_update_78731 : array_update_78720[5];
  assign array_update_78733[6] = add_77421 == 32'h0000_0006 ? array_update_78731 : array_update_78720[6];
  assign array_update_78733[7] = add_77421 == 32'h0000_0007 ? array_update_78731 : array_update_78720[7];
  assign array_update_78733[8] = add_77421 == 32'h0000_0008 ? array_update_78731 : array_update_78720[8];
  assign array_update_78733[9] = add_77421 == 32'h0000_0009 ? array_update_78731 : array_update_78720[9];
  assign array_index_78735 = array_update_72021[add_78732 > 32'h0000_0009 ? 4'h9 : add_78732[3:0]];
  assign array_index_78736 = array_update_78733[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_78740 = smul32b_32b_x_32b(array_index_77428[add_78732 > 32'h0000_0009 ? 4'h9 : add_78732[3:0]], array_index_78735[add_78639 > 32'h0000_0009 ? 4'h9 : add_78639[3:0]]);
  assign add_78742 = array_index_78736[add_78639 > 32'h0000_0009 ? 4'h9 : add_78639[3:0]] + smul_78740;
  assign array_update_78744[0] = add_78639 == 32'h0000_0000 ? add_78742 : array_index_78736[0];
  assign array_update_78744[1] = add_78639 == 32'h0000_0001 ? add_78742 : array_index_78736[1];
  assign array_update_78744[2] = add_78639 == 32'h0000_0002 ? add_78742 : array_index_78736[2];
  assign array_update_78744[3] = add_78639 == 32'h0000_0003 ? add_78742 : array_index_78736[3];
  assign array_update_78744[4] = add_78639 == 32'h0000_0004 ? add_78742 : array_index_78736[4];
  assign array_update_78744[5] = add_78639 == 32'h0000_0005 ? add_78742 : array_index_78736[5];
  assign array_update_78744[6] = add_78639 == 32'h0000_0006 ? add_78742 : array_index_78736[6];
  assign array_update_78744[7] = add_78639 == 32'h0000_0007 ? add_78742 : array_index_78736[7];
  assign array_update_78744[8] = add_78639 == 32'h0000_0008 ? add_78742 : array_index_78736[8];
  assign array_update_78744[9] = add_78639 == 32'h0000_0009 ? add_78742 : array_index_78736[9];
  assign add_78745 = add_78732 + 32'h0000_0001;
  assign array_update_78746[0] = add_77421 == 32'h0000_0000 ? array_update_78744 : array_update_78733[0];
  assign array_update_78746[1] = add_77421 == 32'h0000_0001 ? array_update_78744 : array_update_78733[1];
  assign array_update_78746[2] = add_77421 == 32'h0000_0002 ? array_update_78744 : array_update_78733[2];
  assign array_update_78746[3] = add_77421 == 32'h0000_0003 ? array_update_78744 : array_update_78733[3];
  assign array_update_78746[4] = add_77421 == 32'h0000_0004 ? array_update_78744 : array_update_78733[4];
  assign array_update_78746[5] = add_77421 == 32'h0000_0005 ? array_update_78744 : array_update_78733[5];
  assign array_update_78746[6] = add_77421 == 32'h0000_0006 ? array_update_78744 : array_update_78733[6];
  assign array_update_78746[7] = add_77421 == 32'h0000_0007 ? array_update_78744 : array_update_78733[7];
  assign array_update_78746[8] = add_77421 == 32'h0000_0008 ? array_update_78744 : array_update_78733[8];
  assign array_update_78746[9] = add_77421 == 32'h0000_0009 ? array_update_78744 : array_update_78733[9];
  assign array_index_78748 = array_update_72021[add_78745 > 32'h0000_0009 ? 4'h9 : add_78745[3:0]];
  assign array_index_78749 = array_update_78746[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_78753 = smul32b_32b_x_32b(array_index_77428[add_78745 > 32'h0000_0009 ? 4'h9 : add_78745[3:0]], array_index_78748[add_78639 > 32'h0000_0009 ? 4'h9 : add_78639[3:0]]);
  assign add_78755 = array_index_78749[add_78639 > 32'h0000_0009 ? 4'h9 : add_78639[3:0]] + smul_78753;
  assign array_update_78757[0] = add_78639 == 32'h0000_0000 ? add_78755 : array_index_78749[0];
  assign array_update_78757[1] = add_78639 == 32'h0000_0001 ? add_78755 : array_index_78749[1];
  assign array_update_78757[2] = add_78639 == 32'h0000_0002 ? add_78755 : array_index_78749[2];
  assign array_update_78757[3] = add_78639 == 32'h0000_0003 ? add_78755 : array_index_78749[3];
  assign array_update_78757[4] = add_78639 == 32'h0000_0004 ? add_78755 : array_index_78749[4];
  assign array_update_78757[5] = add_78639 == 32'h0000_0005 ? add_78755 : array_index_78749[5];
  assign array_update_78757[6] = add_78639 == 32'h0000_0006 ? add_78755 : array_index_78749[6];
  assign array_update_78757[7] = add_78639 == 32'h0000_0007 ? add_78755 : array_index_78749[7];
  assign array_update_78757[8] = add_78639 == 32'h0000_0008 ? add_78755 : array_index_78749[8];
  assign array_update_78757[9] = add_78639 == 32'h0000_0009 ? add_78755 : array_index_78749[9];
  assign add_78758 = add_78745 + 32'h0000_0001;
  assign array_update_78759[0] = add_77421 == 32'h0000_0000 ? array_update_78757 : array_update_78746[0];
  assign array_update_78759[1] = add_77421 == 32'h0000_0001 ? array_update_78757 : array_update_78746[1];
  assign array_update_78759[2] = add_77421 == 32'h0000_0002 ? array_update_78757 : array_update_78746[2];
  assign array_update_78759[3] = add_77421 == 32'h0000_0003 ? array_update_78757 : array_update_78746[3];
  assign array_update_78759[4] = add_77421 == 32'h0000_0004 ? array_update_78757 : array_update_78746[4];
  assign array_update_78759[5] = add_77421 == 32'h0000_0005 ? array_update_78757 : array_update_78746[5];
  assign array_update_78759[6] = add_77421 == 32'h0000_0006 ? array_update_78757 : array_update_78746[6];
  assign array_update_78759[7] = add_77421 == 32'h0000_0007 ? array_update_78757 : array_update_78746[7];
  assign array_update_78759[8] = add_77421 == 32'h0000_0008 ? array_update_78757 : array_update_78746[8];
  assign array_update_78759[9] = add_77421 == 32'h0000_0009 ? array_update_78757 : array_update_78746[9];
  assign array_index_78761 = array_update_72021[add_78758 > 32'h0000_0009 ? 4'h9 : add_78758[3:0]];
  assign array_index_78762 = array_update_78759[add_77421 > 32'h0000_0009 ? 4'h9 : add_77421[3:0]];
  assign smul_78766 = smul32b_32b_x_32b(array_index_77428[add_78758 > 32'h0000_0009 ? 4'h9 : add_78758[3:0]], array_index_78761[add_78639 > 32'h0000_0009 ? 4'h9 : add_78639[3:0]]);
  assign add_78768 = array_index_78762[add_78639 > 32'h0000_0009 ? 4'h9 : add_78639[3:0]] + smul_78766;
  assign array_update_78769[0] = add_78639 == 32'h0000_0000 ? add_78768 : array_index_78762[0];
  assign array_update_78769[1] = add_78639 == 32'h0000_0001 ? add_78768 : array_index_78762[1];
  assign array_update_78769[2] = add_78639 == 32'h0000_0002 ? add_78768 : array_index_78762[2];
  assign array_update_78769[3] = add_78639 == 32'h0000_0003 ? add_78768 : array_index_78762[3];
  assign array_update_78769[4] = add_78639 == 32'h0000_0004 ? add_78768 : array_index_78762[4];
  assign array_update_78769[5] = add_78639 == 32'h0000_0005 ? add_78768 : array_index_78762[5];
  assign array_update_78769[6] = add_78639 == 32'h0000_0006 ? add_78768 : array_index_78762[6];
  assign array_update_78769[7] = add_78639 == 32'h0000_0007 ? add_78768 : array_index_78762[7];
  assign array_update_78769[8] = add_78639 == 32'h0000_0008 ? add_78768 : array_index_78762[8];
  assign array_update_78769[9] = add_78639 == 32'h0000_0009 ? add_78768 : array_index_78762[9];
  assign array_update_78771[0] = add_77421 == 32'h0000_0000 ? array_update_78769 : array_update_78759[0];
  assign array_update_78771[1] = add_77421 == 32'h0000_0001 ? array_update_78769 : array_update_78759[1];
  assign array_update_78771[2] = add_77421 == 32'h0000_0002 ? array_update_78769 : array_update_78759[2];
  assign array_update_78771[3] = add_77421 == 32'h0000_0003 ? array_update_78769 : array_update_78759[3];
  assign array_update_78771[4] = add_77421 == 32'h0000_0004 ? array_update_78769 : array_update_78759[4];
  assign array_update_78771[5] = add_77421 == 32'h0000_0005 ? array_update_78769 : array_update_78759[5];
  assign array_update_78771[6] = add_77421 == 32'h0000_0006 ? array_update_78769 : array_update_78759[6];
  assign array_update_78771[7] = add_77421 == 32'h0000_0007 ? array_update_78769 : array_update_78759[7];
  assign array_update_78771[8] = add_77421 == 32'h0000_0008 ? array_update_78769 : array_update_78759[8];
  assign array_update_78771[9] = add_77421 == 32'h0000_0009 ? array_update_78769 : array_update_78759[9];
  assign add_78772 = add_77421 + 32'h0000_0001;
  assign array_index_78773 = array_update_78771[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign literal_78775 = 32'h0000_0000;
  assign array_update_78776[0] = literal_78775 == 32'h0000_0000 ? 32'h0000_0000 : array_index_78773[0];
  assign array_update_78776[1] = literal_78775 == 32'h0000_0001 ? 32'h0000_0000 : array_index_78773[1];
  assign array_update_78776[2] = literal_78775 == 32'h0000_0002 ? 32'h0000_0000 : array_index_78773[2];
  assign array_update_78776[3] = literal_78775 == 32'h0000_0003 ? 32'h0000_0000 : array_index_78773[3];
  assign array_update_78776[4] = literal_78775 == 32'h0000_0004 ? 32'h0000_0000 : array_index_78773[4];
  assign array_update_78776[5] = literal_78775 == 32'h0000_0005 ? 32'h0000_0000 : array_index_78773[5];
  assign array_update_78776[6] = literal_78775 == 32'h0000_0006 ? 32'h0000_0000 : array_index_78773[6];
  assign array_update_78776[7] = literal_78775 == 32'h0000_0007 ? 32'h0000_0000 : array_index_78773[7];
  assign array_update_78776[8] = literal_78775 == 32'h0000_0008 ? 32'h0000_0000 : array_index_78773[8];
  assign array_update_78776[9] = literal_78775 == 32'h0000_0009 ? 32'h0000_0000 : array_index_78773[9];
  assign literal_78777 = 32'h0000_0000;
  assign array_update_78778[0] = add_78772 == 32'h0000_0000 ? array_update_78776 : array_update_78771[0];
  assign array_update_78778[1] = add_78772 == 32'h0000_0001 ? array_update_78776 : array_update_78771[1];
  assign array_update_78778[2] = add_78772 == 32'h0000_0002 ? array_update_78776 : array_update_78771[2];
  assign array_update_78778[3] = add_78772 == 32'h0000_0003 ? array_update_78776 : array_update_78771[3];
  assign array_update_78778[4] = add_78772 == 32'h0000_0004 ? array_update_78776 : array_update_78771[4];
  assign array_update_78778[5] = add_78772 == 32'h0000_0005 ? array_update_78776 : array_update_78771[5];
  assign array_update_78778[6] = add_78772 == 32'h0000_0006 ? array_update_78776 : array_update_78771[6];
  assign array_update_78778[7] = add_78772 == 32'h0000_0007 ? array_update_78776 : array_update_78771[7];
  assign array_update_78778[8] = add_78772 == 32'h0000_0008 ? array_update_78776 : array_update_78771[8];
  assign array_update_78778[9] = add_78772 == 32'h0000_0009 ? array_update_78776 : array_update_78771[9];
  assign array_index_78779 = array_update_72020[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign array_index_78780 = array_update_72021[literal_78777 > 32'h0000_0009 ? 4'h9 : literal_78777[3:0]];
  assign array_index_78781 = array_update_78778[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_78785 = smul32b_32b_x_32b(array_index_78779[literal_78777 > 32'h0000_0009 ? 4'h9 : literal_78777[3:0]], array_index_78780[literal_78775 > 32'h0000_0009 ? 4'h9 : literal_78775[3:0]]);
  assign add_78787 = array_index_78781[literal_78775 > 32'h0000_0009 ? 4'h9 : literal_78775[3:0]] + smul_78785;
  assign array_update_78789[0] = literal_78775 == 32'h0000_0000 ? add_78787 : array_index_78781[0];
  assign array_update_78789[1] = literal_78775 == 32'h0000_0001 ? add_78787 : array_index_78781[1];
  assign array_update_78789[2] = literal_78775 == 32'h0000_0002 ? add_78787 : array_index_78781[2];
  assign array_update_78789[3] = literal_78775 == 32'h0000_0003 ? add_78787 : array_index_78781[3];
  assign array_update_78789[4] = literal_78775 == 32'h0000_0004 ? add_78787 : array_index_78781[4];
  assign array_update_78789[5] = literal_78775 == 32'h0000_0005 ? add_78787 : array_index_78781[5];
  assign array_update_78789[6] = literal_78775 == 32'h0000_0006 ? add_78787 : array_index_78781[6];
  assign array_update_78789[7] = literal_78775 == 32'h0000_0007 ? add_78787 : array_index_78781[7];
  assign array_update_78789[8] = literal_78775 == 32'h0000_0008 ? add_78787 : array_index_78781[8];
  assign array_update_78789[9] = literal_78775 == 32'h0000_0009 ? add_78787 : array_index_78781[9];
  assign add_78790 = literal_78777 + 32'h0000_0001;
  assign array_update_78791[0] = add_78772 == 32'h0000_0000 ? array_update_78789 : array_update_78778[0];
  assign array_update_78791[1] = add_78772 == 32'h0000_0001 ? array_update_78789 : array_update_78778[1];
  assign array_update_78791[2] = add_78772 == 32'h0000_0002 ? array_update_78789 : array_update_78778[2];
  assign array_update_78791[3] = add_78772 == 32'h0000_0003 ? array_update_78789 : array_update_78778[3];
  assign array_update_78791[4] = add_78772 == 32'h0000_0004 ? array_update_78789 : array_update_78778[4];
  assign array_update_78791[5] = add_78772 == 32'h0000_0005 ? array_update_78789 : array_update_78778[5];
  assign array_update_78791[6] = add_78772 == 32'h0000_0006 ? array_update_78789 : array_update_78778[6];
  assign array_update_78791[7] = add_78772 == 32'h0000_0007 ? array_update_78789 : array_update_78778[7];
  assign array_update_78791[8] = add_78772 == 32'h0000_0008 ? array_update_78789 : array_update_78778[8];
  assign array_update_78791[9] = add_78772 == 32'h0000_0009 ? array_update_78789 : array_update_78778[9];
  assign array_index_78793 = array_update_72021[add_78790 > 32'h0000_0009 ? 4'h9 : add_78790[3:0]];
  assign array_index_78794 = array_update_78791[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_78798 = smul32b_32b_x_32b(array_index_78779[add_78790 > 32'h0000_0009 ? 4'h9 : add_78790[3:0]], array_index_78793[literal_78775 > 32'h0000_0009 ? 4'h9 : literal_78775[3:0]]);
  assign add_78800 = array_index_78794[literal_78775 > 32'h0000_0009 ? 4'h9 : literal_78775[3:0]] + smul_78798;
  assign array_update_78802[0] = literal_78775 == 32'h0000_0000 ? add_78800 : array_index_78794[0];
  assign array_update_78802[1] = literal_78775 == 32'h0000_0001 ? add_78800 : array_index_78794[1];
  assign array_update_78802[2] = literal_78775 == 32'h0000_0002 ? add_78800 : array_index_78794[2];
  assign array_update_78802[3] = literal_78775 == 32'h0000_0003 ? add_78800 : array_index_78794[3];
  assign array_update_78802[4] = literal_78775 == 32'h0000_0004 ? add_78800 : array_index_78794[4];
  assign array_update_78802[5] = literal_78775 == 32'h0000_0005 ? add_78800 : array_index_78794[5];
  assign array_update_78802[6] = literal_78775 == 32'h0000_0006 ? add_78800 : array_index_78794[6];
  assign array_update_78802[7] = literal_78775 == 32'h0000_0007 ? add_78800 : array_index_78794[7];
  assign array_update_78802[8] = literal_78775 == 32'h0000_0008 ? add_78800 : array_index_78794[8];
  assign array_update_78802[9] = literal_78775 == 32'h0000_0009 ? add_78800 : array_index_78794[9];
  assign add_78803 = add_78790 + 32'h0000_0001;
  assign array_update_78804[0] = add_78772 == 32'h0000_0000 ? array_update_78802 : array_update_78791[0];
  assign array_update_78804[1] = add_78772 == 32'h0000_0001 ? array_update_78802 : array_update_78791[1];
  assign array_update_78804[2] = add_78772 == 32'h0000_0002 ? array_update_78802 : array_update_78791[2];
  assign array_update_78804[3] = add_78772 == 32'h0000_0003 ? array_update_78802 : array_update_78791[3];
  assign array_update_78804[4] = add_78772 == 32'h0000_0004 ? array_update_78802 : array_update_78791[4];
  assign array_update_78804[5] = add_78772 == 32'h0000_0005 ? array_update_78802 : array_update_78791[5];
  assign array_update_78804[6] = add_78772 == 32'h0000_0006 ? array_update_78802 : array_update_78791[6];
  assign array_update_78804[7] = add_78772 == 32'h0000_0007 ? array_update_78802 : array_update_78791[7];
  assign array_update_78804[8] = add_78772 == 32'h0000_0008 ? array_update_78802 : array_update_78791[8];
  assign array_update_78804[9] = add_78772 == 32'h0000_0009 ? array_update_78802 : array_update_78791[9];
  assign array_index_78806 = array_update_72021[add_78803 > 32'h0000_0009 ? 4'h9 : add_78803[3:0]];
  assign array_index_78807 = array_update_78804[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_78811 = smul32b_32b_x_32b(array_index_78779[add_78803 > 32'h0000_0009 ? 4'h9 : add_78803[3:0]], array_index_78806[literal_78775 > 32'h0000_0009 ? 4'h9 : literal_78775[3:0]]);
  assign add_78813 = array_index_78807[literal_78775 > 32'h0000_0009 ? 4'h9 : literal_78775[3:0]] + smul_78811;
  assign array_update_78815[0] = literal_78775 == 32'h0000_0000 ? add_78813 : array_index_78807[0];
  assign array_update_78815[1] = literal_78775 == 32'h0000_0001 ? add_78813 : array_index_78807[1];
  assign array_update_78815[2] = literal_78775 == 32'h0000_0002 ? add_78813 : array_index_78807[2];
  assign array_update_78815[3] = literal_78775 == 32'h0000_0003 ? add_78813 : array_index_78807[3];
  assign array_update_78815[4] = literal_78775 == 32'h0000_0004 ? add_78813 : array_index_78807[4];
  assign array_update_78815[5] = literal_78775 == 32'h0000_0005 ? add_78813 : array_index_78807[5];
  assign array_update_78815[6] = literal_78775 == 32'h0000_0006 ? add_78813 : array_index_78807[6];
  assign array_update_78815[7] = literal_78775 == 32'h0000_0007 ? add_78813 : array_index_78807[7];
  assign array_update_78815[8] = literal_78775 == 32'h0000_0008 ? add_78813 : array_index_78807[8];
  assign array_update_78815[9] = literal_78775 == 32'h0000_0009 ? add_78813 : array_index_78807[9];
  assign add_78816 = add_78803 + 32'h0000_0001;
  assign array_update_78817[0] = add_78772 == 32'h0000_0000 ? array_update_78815 : array_update_78804[0];
  assign array_update_78817[1] = add_78772 == 32'h0000_0001 ? array_update_78815 : array_update_78804[1];
  assign array_update_78817[2] = add_78772 == 32'h0000_0002 ? array_update_78815 : array_update_78804[2];
  assign array_update_78817[3] = add_78772 == 32'h0000_0003 ? array_update_78815 : array_update_78804[3];
  assign array_update_78817[4] = add_78772 == 32'h0000_0004 ? array_update_78815 : array_update_78804[4];
  assign array_update_78817[5] = add_78772 == 32'h0000_0005 ? array_update_78815 : array_update_78804[5];
  assign array_update_78817[6] = add_78772 == 32'h0000_0006 ? array_update_78815 : array_update_78804[6];
  assign array_update_78817[7] = add_78772 == 32'h0000_0007 ? array_update_78815 : array_update_78804[7];
  assign array_update_78817[8] = add_78772 == 32'h0000_0008 ? array_update_78815 : array_update_78804[8];
  assign array_update_78817[9] = add_78772 == 32'h0000_0009 ? array_update_78815 : array_update_78804[9];
  assign array_index_78819 = array_update_72021[add_78816 > 32'h0000_0009 ? 4'h9 : add_78816[3:0]];
  assign array_index_78820 = array_update_78817[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_78824 = smul32b_32b_x_32b(array_index_78779[add_78816 > 32'h0000_0009 ? 4'h9 : add_78816[3:0]], array_index_78819[literal_78775 > 32'h0000_0009 ? 4'h9 : literal_78775[3:0]]);
  assign add_78826 = array_index_78820[literal_78775 > 32'h0000_0009 ? 4'h9 : literal_78775[3:0]] + smul_78824;
  assign array_update_78828[0] = literal_78775 == 32'h0000_0000 ? add_78826 : array_index_78820[0];
  assign array_update_78828[1] = literal_78775 == 32'h0000_0001 ? add_78826 : array_index_78820[1];
  assign array_update_78828[2] = literal_78775 == 32'h0000_0002 ? add_78826 : array_index_78820[2];
  assign array_update_78828[3] = literal_78775 == 32'h0000_0003 ? add_78826 : array_index_78820[3];
  assign array_update_78828[4] = literal_78775 == 32'h0000_0004 ? add_78826 : array_index_78820[4];
  assign array_update_78828[5] = literal_78775 == 32'h0000_0005 ? add_78826 : array_index_78820[5];
  assign array_update_78828[6] = literal_78775 == 32'h0000_0006 ? add_78826 : array_index_78820[6];
  assign array_update_78828[7] = literal_78775 == 32'h0000_0007 ? add_78826 : array_index_78820[7];
  assign array_update_78828[8] = literal_78775 == 32'h0000_0008 ? add_78826 : array_index_78820[8];
  assign array_update_78828[9] = literal_78775 == 32'h0000_0009 ? add_78826 : array_index_78820[9];
  assign add_78829 = add_78816 + 32'h0000_0001;
  assign array_update_78830[0] = add_78772 == 32'h0000_0000 ? array_update_78828 : array_update_78817[0];
  assign array_update_78830[1] = add_78772 == 32'h0000_0001 ? array_update_78828 : array_update_78817[1];
  assign array_update_78830[2] = add_78772 == 32'h0000_0002 ? array_update_78828 : array_update_78817[2];
  assign array_update_78830[3] = add_78772 == 32'h0000_0003 ? array_update_78828 : array_update_78817[3];
  assign array_update_78830[4] = add_78772 == 32'h0000_0004 ? array_update_78828 : array_update_78817[4];
  assign array_update_78830[5] = add_78772 == 32'h0000_0005 ? array_update_78828 : array_update_78817[5];
  assign array_update_78830[6] = add_78772 == 32'h0000_0006 ? array_update_78828 : array_update_78817[6];
  assign array_update_78830[7] = add_78772 == 32'h0000_0007 ? array_update_78828 : array_update_78817[7];
  assign array_update_78830[8] = add_78772 == 32'h0000_0008 ? array_update_78828 : array_update_78817[8];
  assign array_update_78830[9] = add_78772 == 32'h0000_0009 ? array_update_78828 : array_update_78817[9];
  assign array_index_78832 = array_update_72021[add_78829 > 32'h0000_0009 ? 4'h9 : add_78829[3:0]];
  assign array_index_78833 = array_update_78830[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_78837 = smul32b_32b_x_32b(array_index_78779[add_78829 > 32'h0000_0009 ? 4'h9 : add_78829[3:0]], array_index_78832[literal_78775 > 32'h0000_0009 ? 4'h9 : literal_78775[3:0]]);
  assign add_78839 = array_index_78833[literal_78775 > 32'h0000_0009 ? 4'h9 : literal_78775[3:0]] + smul_78837;
  assign array_update_78841[0] = literal_78775 == 32'h0000_0000 ? add_78839 : array_index_78833[0];
  assign array_update_78841[1] = literal_78775 == 32'h0000_0001 ? add_78839 : array_index_78833[1];
  assign array_update_78841[2] = literal_78775 == 32'h0000_0002 ? add_78839 : array_index_78833[2];
  assign array_update_78841[3] = literal_78775 == 32'h0000_0003 ? add_78839 : array_index_78833[3];
  assign array_update_78841[4] = literal_78775 == 32'h0000_0004 ? add_78839 : array_index_78833[4];
  assign array_update_78841[5] = literal_78775 == 32'h0000_0005 ? add_78839 : array_index_78833[5];
  assign array_update_78841[6] = literal_78775 == 32'h0000_0006 ? add_78839 : array_index_78833[6];
  assign array_update_78841[7] = literal_78775 == 32'h0000_0007 ? add_78839 : array_index_78833[7];
  assign array_update_78841[8] = literal_78775 == 32'h0000_0008 ? add_78839 : array_index_78833[8];
  assign array_update_78841[9] = literal_78775 == 32'h0000_0009 ? add_78839 : array_index_78833[9];
  assign add_78842 = add_78829 + 32'h0000_0001;
  assign array_update_78843[0] = add_78772 == 32'h0000_0000 ? array_update_78841 : array_update_78830[0];
  assign array_update_78843[1] = add_78772 == 32'h0000_0001 ? array_update_78841 : array_update_78830[1];
  assign array_update_78843[2] = add_78772 == 32'h0000_0002 ? array_update_78841 : array_update_78830[2];
  assign array_update_78843[3] = add_78772 == 32'h0000_0003 ? array_update_78841 : array_update_78830[3];
  assign array_update_78843[4] = add_78772 == 32'h0000_0004 ? array_update_78841 : array_update_78830[4];
  assign array_update_78843[5] = add_78772 == 32'h0000_0005 ? array_update_78841 : array_update_78830[5];
  assign array_update_78843[6] = add_78772 == 32'h0000_0006 ? array_update_78841 : array_update_78830[6];
  assign array_update_78843[7] = add_78772 == 32'h0000_0007 ? array_update_78841 : array_update_78830[7];
  assign array_update_78843[8] = add_78772 == 32'h0000_0008 ? array_update_78841 : array_update_78830[8];
  assign array_update_78843[9] = add_78772 == 32'h0000_0009 ? array_update_78841 : array_update_78830[9];
  assign array_index_78845 = array_update_72021[add_78842 > 32'h0000_0009 ? 4'h9 : add_78842[3:0]];
  assign array_index_78846 = array_update_78843[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_78850 = smul32b_32b_x_32b(array_index_78779[add_78842 > 32'h0000_0009 ? 4'h9 : add_78842[3:0]], array_index_78845[literal_78775 > 32'h0000_0009 ? 4'h9 : literal_78775[3:0]]);
  assign add_78852 = array_index_78846[literal_78775 > 32'h0000_0009 ? 4'h9 : literal_78775[3:0]] + smul_78850;
  assign array_update_78854[0] = literal_78775 == 32'h0000_0000 ? add_78852 : array_index_78846[0];
  assign array_update_78854[1] = literal_78775 == 32'h0000_0001 ? add_78852 : array_index_78846[1];
  assign array_update_78854[2] = literal_78775 == 32'h0000_0002 ? add_78852 : array_index_78846[2];
  assign array_update_78854[3] = literal_78775 == 32'h0000_0003 ? add_78852 : array_index_78846[3];
  assign array_update_78854[4] = literal_78775 == 32'h0000_0004 ? add_78852 : array_index_78846[4];
  assign array_update_78854[5] = literal_78775 == 32'h0000_0005 ? add_78852 : array_index_78846[5];
  assign array_update_78854[6] = literal_78775 == 32'h0000_0006 ? add_78852 : array_index_78846[6];
  assign array_update_78854[7] = literal_78775 == 32'h0000_0007 ? add_78852 : array_index_78846[7];
  assign array_update_78854[8] = literal_78775 == 32'h0000_0008 ? add_78852 : array_index_78846[8];
  assign array_update_78854[9] = literal_78775 == 32'h0000_0009 ? add_78852 : array_index_78846[9];
  assign add_78855 = add_78842 + 32'h0000_0001;
  assign array_update_78856[0] = add_78772 == 32'h0000_0000 ? array_update_78854 : array_update_78843[0];
  assign array_update_78856[1] = add_78772 == 32'h0000_0001 ? array_update_78854 : array_update_78843[1];
  assign array_update_78856[2] = add_78772 == 32'h0000_0002 ? array_update_78854 : array_update_78843[2];
  assign array_update_78856[3] = add_78772 == 32'h0000_0003 ? array_update_78854 : array_update_78843[3];
  assign array_update_78856[4] = add_78772 == 32'h0000_0004 ? array_update_78854 : array_update_78843[4];
  assign array_update_78856[5] = add_78772 == 32'h0000_0005 ? array_update_78854 : array_update_78843[5];
  assign array_update_78856[6] = add_78772 == 32'h0000_0006 ? array_update_78854 : array_update_78843[6];
  assign array_update_78856[7] = add_78772 == 32'h0000_0007 ? array_update_78854 : array_update_78843[7];
  assign array_update_78856[8] = add_78772 == 32'h0000_0008 ? array_update_78854 : array_update_78843[8];
  assign array_update_78856[9] = add_78772 == 32'h0000_0009 ? array_update_78854 : array_update_78843[9];
  assign array_index_78858 = array_update_72021[add_78855 > 32'h0000_0009 ? 4'h9 : add_78855[3:0]];
  assign array_index_78859 = array_update_78856[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_78863 = smul32b_32b_x_32b(array_index_78779[add_78855 > 32'h0000_0009 ? 4'h9 : add_78855[3:0]], array_index_78858[literal_78775 > 32'h0000_0009 ? 4'h9 : literal_78775[3:0]]);
  assign add_78865 = array_index_78859[literal_78775 > 32'h0000_0009 ? 4'h9 : literal_78775[3:0]] + smul_78863;
  assign array_update_78867[0] = literal_78775 == 32'h0000_0000 ? add_78865 : array_index_78859[0];
  assign array_update_78867[1] = literal_78775 == 32'h0000_0001 ? add_78865 : array_index_78859[1];
  assign array_update_78867[2] = literal_78775 == 32'h0000_0002 ? add_78865 : array_index_78859[2];
  assign array_update_78867[3] = literal_78775 == 32'h0000_0003 ? add_78865 : array_index_78859[3];
  assign array_update_78867[4] = literal_78775 == 32'h0000_0004 ? add_78865 : array_index_78859[4];
  assign array_update_78867[5] = literal_78775 == 32'h0000_0005 ? add_78865 : array_index_78859[5];
  assign array_update_78867[6] = literal_78775 == 32'h0000_0006 ? add_78865 : array_index_78859[6];
  assign array_update_78867[7] = literal_78775 == 32'h0000_0007 ? add_78865 : array_index_78859[7];
  assign array_update_78867[8] = literal_78775 == 32'h0000_0008 ? add_78865 : array_index_78859[8];
  assign array_update_78867[9] = literal_78775 == 32'h0000_0009 ? add_78865 : array_index_78859[9];
  assign add_78868 = add_78855 + 32'h0000_0001;
  assign array_update_78869[0] = add_78772 == 32'h0000_0000 ? array_update_78867 : array_update_78856[0];
  assign array_update_78869[1] = add_78772 == 32'h0000_0001 ? array_update_78867 : array_update_78856[1];
  assign array_update_78869[2] = add_78772 == 32'h0000_0002 ? array_update_78867 : array_update_78856[2];
  assign array_update_78869[3] = add_78772 == 32'h0000_0003 ? array_update_78867 : array_update_78856[3];
  assign array_update_78869[4] = add_78772 == 32'h0000_0004 ? array_update_78867 : array_update_78856[4];
  assign array_update_78869[5] = add_78772 == 32'h0000_0005 ? array_update_78867 : array_update_78856[5];
  assign array_update_78869[6] = add_78772 == 32'h0000_0006 ? array_update_78867 : array_update_78856[6];
  assign array_update_78869[7] = add_78772 == 32'h0000_0007 ? array_update_78867 : array_update_78856[7];
  assign array_update_78869[8] = add_78772 == 32'h0000_0008 ? array_update_78867 : array_update_78856[8];
  assign array_update_78869[9] = add_78772 == 32'h0000_0009 ? array_update_78867 : array_update_78856[9];
  assign array_index_78871 = array_update_72021[add_78868 > 32'h0000_0009 ? 4'h9 : add_78868[3:0]];
  assign array_index_78872 = array_update_78869[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_78876 = smul32b_32b_x_32b(array_index_78779[add_78868 > 32'h0000_0009 ? 4'h9 : add_78868[3:0]], array_index_78871[literal_78775 > 32'h0000_0009 ? 4'h9 : literal_78775[3:0]]);
  assign add_78878 = array_index_78872[literal_78775 > 32'h0000_0009 ? 4'h9 : literal_78775[3:0]] + smul_78876;
  assign array_update_78880[0] = literal_78775 == 32'h0000_0000 ? add_78878 : array_index_78872[0];
  assign array_update_78880[1] = literal_78775 == 32'h0000_0001 ? add_78878 : array_index_78872[1];
  assign array_update_78880[2] = literal_78775 == 32'h0000_0002 ? add_78878 : array_index_78872[2];
  assign array_update_78880[3] = literal_78775 == 32'h0000_0003 ? add_78878 : array_index_78872[3];
  assign array_update_78880[4] = literal_78775 == 32'h0000_0004 ? add_78878 : array_index_78872[4];
  assign array_update_78880[5] = literal_78775 == 32'h0000_0005 ? add_78878 : array_index_78872[5];
  assign array_update_78880[6] = literal_78775 == 32'h0000_0006 ? add_78878 : array_index_78872[6];
  assign array_update_78880[7] = literal_78775 == 32'h0000_0007 ? add_78878 : array_index_78872[7];
  assign array_update_78880[8] = literal_78775 == 32'h0000_0008 ? add_78878 : array_index_78872[8];
  assign array_update_78880[9] = literal_78775 == 32'h0000_0009 ? add_78878 : array_index_78872[9];
  assign add_78881 = add_78868 + 32'h0000_0001;
  assign array_update_78882[0] = add_78772 == 32'h0000_0000 ? array_update_78880 : array_update_78869[0];
  assign array_update_78882[1] = add_78772 == 32'h0000_0001 ? array_update_78880 : array_update_78869[1];
  assign array_update_78882[2] = add_78772 == 32'h0000_0002 ? array_update_78880 : array_update_78869[2];
  assign array_update_78882[3] = add_78772 == 32'h0000_0003 ? array_update_78880 : array_update_78869[3];
  assign array_update_78882[4] = add_78772 == 32'h0000_0004 ? array_update_78880 : array_update_78869[4];
  assign array_update_78882[5] = add_78772 == 32'h0000_0005 ? array_update_78880 : array_update_78869[5];
  assign array_update_78882[6] = add_78772 == 32'h0000_0006 ? array_update_78880 : array_update_78869[6];
  assign array_update_78882[7] = add_78772 == 32'h0000_0007 ? array_update_78880 : array_update_78869[7];
  assign array_update_78882[8] = add_78772 == 32'h0000_0008 ? array_update_78880 : array_update_78869[8];
  assign array_update_78882[9] = add_78772 == 32'h0000_0009 ? array_update_78880 : array_update_78869[9];
  assign array_index_78884 = array_update_72021[add_78881 > 32'h0000_0009 ? 4'h9 : add_78881[3:0]];
  assign array_index_78885 = array_update_78882[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_78889 = smul32b_32b_x_32b(array_index_78779[add_78881 > 32'h0000_0009 ? 4'h9 : add_78881[3:0]], array_index_78884[literal_78775 > 32'h0000_0009 ? 4'h9 : literal_78775[3:0]]);
  assign add_78891 = array_index_78885[literal_78775 > 32'h0000_0009 ? 4'h9 : literal_78775[3:0]] + smul_78889;
  assign array_update_78893[0] = literal_78775 == 32'h0000_0000 ? add_78891 : array_index_78885[0];
  assign array_update_78893[1] = literal_78775 == 32'h0000_0001 ? add_78891 : array_index_78885[1];
  assign array_update_78893[2] = literal_78775 == 32'h0000_0002 ? add_78891 : array_index_78885[2];
  assign array_update_78893[3] = literal_78775 == 32'h0000_0003 ? add_78891 : array_index_78885[3];
  assign array_update_78893[4] = literal_78775 == 32'h0000_0004 ? add_78891 : array_index_78885[4];
  assign array_update_78893[5] = literal_78775 == 32'h0000_0005 ? add_78891 : array_index_78885[5];
  assign array_update_78893[6] = literal_78775 == 32'h0000_0006 ? add_78891 : array_index_78885[6];
  assign array_update_78893[7] = literal_78775 == 32'h0000_0007 ? add_78891 : array_index_78885[7];
  assign array_update_78893[8] = literal_78775 == 32'h0000_0008 ? add_78891 : array_index_78885[8];
  assign array_update_78893[9] = literal_78775 == 32'h0000_0009 ? add_78891 : array_index_78885[9];
  assign add_78894 = add_78881 + 32'h0000_0001;
  assign array_update_78895[0] = add_78772 == 32'h0000_0000 ? array_update_78893 : array_update_78882[0];
  assign array_update_78895[1] = add_78772 == 32'h0000_0001 ? array_update_78893 : array_update_78882[1];
  assign array_update_78895[2] = add_78772 == 32'h0000_0002 ? array_update_78893 : array_update_78882[2];
  assign array_update_78895[3] = add_78772 == 32'h0000_0003 ? array_update_78893 : array_update_78882[3];
  assign array_update_78895[4] = add_78772 == 32'h0000_0004 ? array_update_78893 : array_update_78882[4];
  assign array_update_78895[5] = add_78772 == 32'h0000_0005 ? array_update_78893 : array_update_78882[5];
  assign array_update_78895[6] = add_78772 == 32'h0000_0006 ? array_update_78893 : array_update_78882[6];
  assign array_update_78895[7] = add_78772 == 32'h0000_0007 ? array_update_78893 : array_update_78882[7];
  assign array_update_78895[8] = add_78772 == 32'h0000_0008 ? array_update_78893 : array_update_78882[8];
  assign array_update_78895[9] = add_78772 == 32'h0000_0009 ? array_update_78893 : array_update_78882[9];
  assign array_index_78897 = array_update_72021[add_78894 > 32'h0000_0009 ? 4'h9 : add_78894[3:0]];
  assign array_index_78898 = array_update_78895[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_78902 = smul32b_32b_x_32b(array_index_78779[add_78894 > 32'h0000_0009 ? 4'h9 : add_78894[3:0]], array_index_78897[literal_78775 > 32'h0000_0009 ? 4'h9 : literal_78775[3:0]]);
  assign add_78904 = array_index_78898[literal_78775 > 32'h0000_0009 ? 4'h9 : literal_78775[3:0]] + smul_78902;
  assign array_update_78905[0] = literal_78775 == 32'h0000_0000 ? add_78904 : array_index_78898[0];
  assign array_update_78905[1] = literal_78775 == 32'h0000_0001 ? add_78904 : array_index_78898[1];
  assign array_update_78905[2] = literal_78775 == 32'h0000_0002 ? add_78904 : array_index_78898[2];
  assign array_update_78905[3] = literal_78775 == 32'h0000_0003 ? add_78904 : array_index_78898[3];
  assign array_update_78905[4] = literal_78775 == 32'h0000_0004 ? add_78904 : array_index_78898[4];
  assign array_update_78905[5] = literal_78775 == 32'h0000_0005 ? add_78904 : array_index_78898[5];
  assign array_update_78905[6] = literal_78775 == 32'h0000_0006 ? add_78904 : array_index_78898[6];
  assign array_update_78905[7] = literal_78775 == 32'h0000_0007 ? add_78904 : array_index_78898[7];
  assign array_update_78905[8] = literal_78775 == 32'h0000_0008 ? add_78904 : array_index_78898[8];
  assign array_update_78905[9] = literal_78775 == 32'h0000_0009 ? add_78904 : array_index_78898[9];
  assign array_update_78906[0] = add_78772 == 32'h0000_0000 ? array_update_78905 : array_update_78895[0];
  assign array_update_78906[1] = add_78772 == 32'h0000_0001 ? array_update_78905 : array_update_78895[1];
  assign array_update_78906[2] = add_78772 == 32'h0000_0002 ? array_update_78905 : array_update_78895[2];
  assign array_update_78906[3] = add_78772 == 32'h0000_0003 ? array_update_78905 : array_update_78895[3];
  assign array_update_78906[4] = add_78772 == 32'h0000_0004 ? array_update_78905 : array_update_78895[4];
  assign array_update_78906[5] = add_78772 == 32'h0000_0005 ? array_update_78905 : array_update_78895[5];
  assign array_update_78906[6] = add_78772 == 32'h0000_0006 ? array_update_78905 : array_update_78895[6];
  assign array_update_78906[7] = add_78772 == 32'h0000_0007 ? array_update_78905 : array_update_78895[7];
  assign array_update_78906[8] = add_78772 == 32'h0000_0008 ? array_update_78905 : array_update_78895[8];
  assign array_update_78906[9] = add_78772 == 32'h0000_0009 ? array_update_78905 : array_update_78895[9];
  assign array_index_78908 = array_update_78906[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign add_78910 = literal_78775 + 32'h0000_0001;
  assign array_update_78911[0] = add_78910 == 32'h0000_0000 ? 32'h0000_0000 : array_index_78908[0];
  assign array_update_78911[1] = add_78910 == 32'h0000_0001 ? 32'h0000_0000 : array_index_78908[1];
  assign array_update_78911[2] = add_78910 == 32'h0000_0002 ? 32'h0000_0000 : array_index_78908[2];
  assign array_update_78911[3] = add_78910 == 32'h0000_0003 ? 32'h0000_0000 : array_index_78908[3];
  assign array_update_78911[4] = add_78910 == 32'h0000_0004 ? 32'h0000_0000 : array_index_78908[4];
  assign array_update_78911[5] = add_78910 == 32'h0000_0005 ? 32'h0000_0000 : array_index_78908[5];
  assign array_update_78911[6] = add_78910 == 32'h0000_0006 ? 32'h0000_0000 : array_index_78908[6];
  assign array_update_78911[7] = add_78910 == 32'h0000_0007 ? 32'h0000_0000 : array_index_78908[7];
  assign array_update_78911[8] = add_78910 == 32'h0000_0008 ? 32'h0000_0000 : array_index_78908[8];
  assign array_update_78911[9] = add_78910 == 32'h0000_0009 ? 32'h0000_0000 : array_index_78908[9];
  assign literal_78912 = 32'h0000_0000;
  assign array_update_78913[0] = add_78772 == 32'h0000_0000 ? array_update_78911 : array_update_78906[0];
  assign array_update_78913[1] = add_78772 == 32'h0000_0001 ? array_update_78911 : array_update_78906[1];
  assign array_update_78913[2] = add_78772 == 32'h0000_0002 ? array_update_78911 : array_update_78906[2];
  assign array_update_78913[3] = add_78772 == 32'h0000_0003 ? array_update_78911 : array_update_78906[3];
  assign array_update_78913[4] = add_78772 == 32'h0000_0004 ? array_update_78911 : array_update_78906[4];
  assign array_update_78913[5] = add_78772 == 32'h0000_0005 ? array_update_78911 : array_update_78906[5];
  assign array_update_78913[6] = add_78772 == 32'h0000_0006 ? array_update_78911 : array_update_78906[6];
  assign array_update_78913[7] = add_78772 == 32'h0000_0007 ? array_update_78911 : array_update_78906[7];
  assign array_update_78913[8] = add_78772 == 32'h0000_0008 ? array_update_78911 : array_update_78906[8];
  assign array_update_78913[9] = add_78772 == 32'h0000_0009 ? array_update_78911 : array_update_78906[9];
  assign array_index_78915 = array_update_72021[literal_78912 > 32'h0000_0009 ? 4'h9 : literal_78912[3:0]];
  assign array_index_78916 = array_update_78913[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_78920 = smul32b_32b_x_32b(array_index_78779[literal_78912 > 32'h0000_0009 ? 4'h9 : literal_78912[3:0]], array_index_78915[add_78910 > 32'h0000_0009 ? 4'h9 : add_78910[3:0]]);
  assign add_78922 = array_index_78916[add_78910 > 32'h0000_0009 ? 4'h9 : add_78910[3:0]] + smul_78920;
  assign array_update_78924[0] = add_78910 == 32'h0000_0000 ? add_78922 : array_index_78916[0];
  assign array_update_78924[1] = add_78910 == 32'h0000_0001 ? add_78922 : array_index_78916[1];
  assign array_update_78924[2] = add_78910 == 32'h0000_0002 ? add_78922 : array_index_78916[2];
  assign array_update_78924[3] = add_78910 == 32'h0000_0003 ? add_78922 : array_index_78916[3];
  assign array_update_78924[4] = add_78910 == 32'h0000_0004 ? add_78922 : array_index_78916[4];
  assign array_update_78924[5] = add_78910 == 32'h0000_0005 ? add_78922 : array_index_78916[5];
  assign array_update_78924[6] = add_78910 == 32'h0000_0006 ? add_78922 : array_index_78916[6];
  assign array_update_78924[7] = add_78910 == 32'h0000_0007 ? add_78922 : array_index_78916[7];
  assign array_update_78924[8] = add_78910 == 32'h0000_0008 ? add_78922 : array_index_78916[8];
  assign array_update_78924[9] = add_78910 == 32'h0000_0009 ? add_78922 : array_index_78916[9];
  assign add_78925 = literal_78912 + 32'h0000_0001;
  assign array_update_78926[0] = add_78772 == 32'h0000_0000 ? array_update_78924 : array_update_78913[0];
  assign array_update_78926[1] = add_78772 == 32'h0000_0001 ? array_update_78924 : array_update_78913[1];
  assign array_update_78926[2] = add_78772 == 32'h0000_0002 ? array_update_78924 : array_update_78913[2];
  assign array_update_78926[3] = add_78772 == 32'h0000_0003 ? array_update_78924 : array_update_78913[3];
  assign array_update_78926[4] = add_78772 == 32'h0000_0004 ? array_update_78924 : array_update_78913[4];
  assign array_update_78926[5] = add_78772 == 32'h0000_0005 ? array_update_78924 : array_update_78913[5];
  assign array_update_78926[6] = add_78772 == 32'h0000_0006 ? array_update_78924 : array_update_78913[6];
  assign array_update_78926[7] = add_78772 == 32'h0000_0007 ? array_update_78924 : array_update_78913[7];
  assign array_update_78926[8] = add_78772 == 32'h0000_0008 ? array_update_78924 : array_update_78913[8];
  assign array_update_78926[9] = add_78772 == 32'h0000_0009 ? array_update_78924 : array_update_78913[9];
  assign array_index_78928 = array_update_72021[add_78925 > 32'h0000_0009 ? 4'h9 : add_78925[3:0]];
  assign array_index_78929 = array_update_78926[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_78933 = smul32b_32b_x_32b(array_index_78779[add_78925 > 32'h0000_0009 ? 4'h9 : add_78925[3:0]], array_index_78928[add_78910 > 32'h0000_0009 ? 4'h9 : add_78910[3:0]]);
  assign add_78935 = array_index_78929[add_78910 > 32'h0000_0009 ? 4'h9 : add_78910[3:0]] + smul_78933;
  assign array_update_78937[0] = add_78910 == 32'h0000_0000 ? add_78935 : array_index_78929[0];
  assign array_update_78937[1] = add_78910 == 32'h0000_0001 ? add_78935 : array_index_78929[1];
  assign array_update_78937[2] = add_78910 == 32'h0000_0002 ? add_78935 : array_index_78929[2];
  assign array_update_78937[3] = add_78910 == 32'h0000_0003 ? add_78935 : array_index_78929[3];
  assign array_update_78937[4] = add_78910 == 32'h0000_0004 ? add_78935 : array_index_78929[4];
  assign array_update_78937[5] = add_78910 == 32'h0000_0005 ? add_78935 : array_index_78929[5];
  assign array_update_78937[6] = add_78910 == 32'h0000_0006 ? add_78935 : array_index_78929[6];
  assign array_update_78937[7] = add_78910 == 32'h0000_0007 ? add_78935 : array_index_78929[7];
  assign array_update_78937[8] = add_78910 == 32'h0000_0008 ? add_78935 : array_index_78929[8];
  assign array_update_78937[9] = add_78910 == 32'h0000_0009 ? add_78935 : array_index_78929[9];
  assign add_78938 = add_78925 + 32'h0000_0001;
  assign array_update_78939[0] = add_78772 == 32'h0000_0000 ? array_update_78937 : array_update_78926[0];
  assign array_update_78939[1] = add_78772 == 32'h0000_0001 ? array_update_78937 : array_update_78926[1];
  assign array_update_78939[2] = add_78772 == 32'h0000_0002 ? array_update_78937 : array_update_78926[2];
  assign array_update_78939[3] = add_78772 == 32'h0000_0003 ? array_update_78937 : array_update_78926[3];
  assign array_update_78939[4] = add_78772 == 32'h0000_0004 ? array_update_78937 : array_update_78926[4];
  assign array_update_78939[5] = add_78772 == 32'h0000_0005 ? array_update_78937 : array_update_78926[5];
  assign array_update_78939[6] = add_78772 == 32'h0000_0006 ? array_update_78937 : array_update_78926[6];
  assign array_update_78939[7] = add_78772 == 32'h0000_0007 ? array_update_78937 : array_update_78926[7];
  assign array_update_78939[8] = add_78772 == 32'h0000_0008 ? array_update_78937 : array_update_78926[8];
  assign array_update_78939[9] = add_78772 == 32'h0000_0009 ? array_update_78937 : array_update_78926[9];
  assign array_index_78941 = array_update_72021[add_78938 > 32'h0000_0009 ? 4'h9 : add_78938[3:0]];
  assign array_index_78942 = array_update_78939[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_78946 = smul32b_32b_x_32b(array_index_78779[add_78938 > 32'h0000_0009 ? 4'h9 : add_78938[3:0]], array_index_78941[add_78910 > 32'h0000_0009 ? 4'h9 : add_78910[3:0]]);
  assign add_78948 = array_index_78942[add_78910 > 32'h0000_0009 ? 4'h9 : add_78910[3:0]] + smul_78946;
  assign array_update_78950[0] = add_78910 == 32'h0000_0000 ? add_78948 : array_index_78942[0];
  assign array_update_78950[1] = add_78910 == 32'h0000_0001 ? add_78948 : array_index_78942[1];
  assign array_update_78950[2] = add_78910 == 32'h0000_0002 ? add_78948 : array_index_78942[2];
  assign array_update_78950[3] = add_78910 == 32'h0000_0003 ? add_78948 : array_index_78942[3];
  assign array_update_78950[4] = add_78910 == 32'h0000_0004 ? add_78948 : array_index_78942[4];
  assign array_update_78950[5] = add_78910 == 32'h0000_0005 ? add_78948 : array_index_78942[5];
  assign array_update_78950[6] = add_78910 == 32'h0000_0006 ? add_78948 : array_index_78942[6];
  assign array_update_78950[7] = add_78910 == 32'h0000_0007 ? add_78948 : array_index_78942[7];
  assign array_update_78950[8] = add_78910 == 32'h0000_0008 ? add_78948 : array_index_78942[8];
  assign array_update_78950[9] = add_78910 == 32'h0000_0009 ? add_78948 : array_index_78942[9];
  assign add_78951 = add_78938 + 32'h0000_0001;
  assign array_update_78952[0] = add_78772 == 32'h0000_0000 ? array_update_78950 : array_update_78939[0];
  assign array_update_78952[1] = add_78772 == 32'h0000_0001 ? array_update_78950 : array_update_78939[1];
  assign array_update_78952[2] = add_78772 == 32'h0000_0002 ? array_update_78950 : array_update_78939[2];
  assign array_update_78952[3] = add_78772 == 32'h0000_0003 ? array_update_78950 : array_update_78939[3];
  assign array_update_78952[4] = add_78772 == 32'h0000_0004 ? array_update_78950 : array_update_78939[4];
  assign array_update_78952[5] = add_78772 == 32'h0000_0005 ? array_update_78950 : array_update_78939[5];
  assign array_update_78952[6] = add_78772 == 32'h0000_0006 ? array_update_78950 : array_update_78939[6];
  assign array_update_78952[7] = add_78772 == 32'h0000_0007 ? array_update_78950 : array_update_78939[7];
  assign array_update_78952[8] = add_78772 == 32'h0000_0008 ? array_update_78950 : array_update_78939[8];
  assign array_update_78952[9] = add_78772 == 32'h0000_0009 ? array_update_78950 : array_update_78939[9];
  assign array_index_78954 = array_update_72021[add_78951 > 32'h0000_0009 ? 4'h9 : add_78951[3:0]];
  assign array_index_78955 = array_update_78952[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_78959 = smul32b_32b_x_32b(array_index_78779[add_78951 > 32'h0000_0009 ? 4'h9 : add_78951[3:0]], array_index_78954[add_78910 > 32'h0000_0009 ? 4'h9 : add_78910[3:0]]);
  assign add_78961 = array_index_78955[add_78910 > 32'h0000_0009 ? 4'h9 : add_78910[3:0]] + smul_78959;
  assign array_update_78963[0] = add_78910 == 32'h0000_0000 ? add_78961 : array_index_78955[0];
  assign array_update_78963[1] = add_78910 == 32'h0000_0001 ? add_78961 : array_index_78955[1];
  assign array_update_78963[2] = add_78910 == 32'h0000_0002 ? add_78961 : array_index_78955[2];
  assign array_update_78963[3] = add_78910 == 32'h0000_0003 ? add_78961 : array_index_78955[3];
  assign array_update_78963[4] = add_78910 == 32'h0000_0004 ? add_78961 : array_index_78955[4];
  assign array_update_78963[5] = add_78910 == 32'h0000_0005 ? add_78961 : array_index_78955[5];
  assign array_update_78963[6] = add_78910 == 32'h0000_0006 ? add_78961 : array_index_78955[6];
  assign array_update_78963[7] = add_78910 == 32'h0000_0007 ? add_78961 : array_index_78955[7];
  assign array_update_78963[8] = add_78910 == 32'h0000_0008 ? add_78961 : array_index_78955[8];
  assign array_update_78963[9] = add_78910 == 32'h0000_0009 ? add_78961 : array_index_78955[9];
  assign add_78964 = add_78951 + 32'h0000_0001;
  assign array_update_78965[0] = add_78772 == 32'h0000_0000 ? array_update_78963 : array_update_78952[0];
  assign array_update_78965[1] = add_78772 == 32'h0000_0001 ? array_update_78963 : array_update_78952[1];
  assign array_update_78965[2] = add_78772 == 32'h0000_0002 ? array_update_78963 : array_update_78952[2];
  assign array_update_78965[3] = add_78772 == 32'h0000_0003 ? array_update_78963 : array_update_78952[3];
  assign array_update_78965[4] = add_78772 == 32'h0000_0004 ? array_update_78963 : array_update_78952[4];
  assign array_update_78965[5] = add_78772 == 32'h0000_0005 ? array_update_78963 : array_update_78952[5];
  assign array_update_78965[6] = add_78772 == 32'h0000_0006 ? array_update_78963 : array_update_78952[6];
  assign array_update_78965[7] = add_78772 == 32'h0000_0007 ? array_update_78963 : array_update_78952[7];
  assign array_update_78965[8] = add_78772 == 32'h0000_0008 ? array_update_78963 : array_update_78952[8];
  assign array_update_78965[9] = add_78772 == 32'h0000_0009 ? array_update_78963 : array_update_78952[9];
  assign array_index_78967 = array_update_72021[add_78964 > 32'h0000_0009 ? 4'h9 : add_78964[3:0]];
  assign array_index_78968 = array_update_78965[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_78972 = smul32b_32b_x_32b(array_index_78779[add_78964 > 32'h0000_0009 ? 4'h9 : add_78964[3:0]], array_index_78967[add_78910 > 32'h0000_0009 ? 4'h9 : add_78910[3:0]]);
  assign add_78974 = array_index_78968[add_78910 > 32'h0000_0009 ? 4'h9 : add_78910[3:0]] + smul_78972;
  assign array_update_78976[0] = add_78910 == 32'h0000_0000 ? add_78974 : array_index_78968[0];
  assign array_update_78976[1] = add_78910 == 32'h0000_0001 ? add_78974 : array_index_78968[1];
  assign array_update_78976[2] = add_78910 == 32'h0000_0002 ? add_78974 : array_index_78968[2];
  assign array_update_78976[3] = add_78910 == 32'h0000_0003 ? add_78974 : array_index_78968[3];
  assign array_update_78976[4] = add_78910 == 32'h0000_0004 ? add_78974 : array_index_78968[4];
  assign array_update_78976[5] = add_78910 == 32'h0000_0005 ? add_78974 : array_index_78968[5];
  assign array_update_78976[6] = add_78910 == 32'h0000_0006 ? add_78974 : array_index_78968[6];
  assign array_update_78976[7] = add_78910 == 32'h0000_0007 ? add_78974 : array_index_78968[7];
  assign array_update_78976[8] = add_78910 == 32'h0000_0008 ? add_78974 : array_index_78968[8];
  assign array_update_78976[9] = add_78910 == 32'h0000_0009 ? add_78974 : array_index_78968[9];
  assign add_78977 = add_78964 + 32'h0000_0001;
  assign array_update_78978[0] = add_78772 == 32'h0000_0000 ? array_update_78976 : array_update_78965[0];
  assign array_update_78978[1] = add_78772 == 32'h0000_0001 ? array_update_78976 : array_update_78965[1];
  assign array_update_78978[2] = add_78772 == 32'h0000_0002 ? array_update_78976 : array_update_78965[2];
  assign array_update_78978[3] = add_78772 == 32'h0000_0003 ? array_update_78976 : array_update_78965[3];
  assign array_update_78978[4] = add_78772 == 32'h0000_0004 ? array_update_78976 : array_update_78965[4];
  assign array_update_78978[5] = add_78772 == 32'h0000_0005 ? array_update_78976 : array_update_78965[5];
  assign array_update_78978[6] = add_78772 == 32'h0000_0006 ? array_update_78976 : array_update_78965[6];
  assign array_update_78978[7] = add_78772 == 32'h0000_0007 ? array_update_78976 : array_update_78965[7];
  assign array_update_78978[8] = add_78772 == 32'h0000_0008 ? array_update_78976 : array_update_78965[8];
  assign array_update_78978[9] = add_78772 == 32'h0000_0009 ? array_update_78976 : array_update_78965[9];
  assign array_index_78980 = array_update_72021[add_78977 > 32'h0000_0009 ? 4'h9 : add_78977[3:0]];
  assign array_index_78981 = array_update_78978[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_78985 = smul32b_32b_x_32b(array_index_78779[add_78977 > 32'h0000_0009 ? 4'h9 : add_78977[3:0]], array_index_78980[add_78910 > 32'h0000_0009 ? 4'h9 : add_78910[3:0]]);
  assign add_78987 = array_index_78981[add_78910 > 32'h0000_0009 ? 4'h9 : add_78910[3:0]] + smul_78985;
  assign array_update_78989[0] = add_78910 == 32'h0000_0000 ? add_78987 : array_index_78981[0];
  assign array_update_78989[1] = add_78910 == 32'h0000_0001 ? add_78987 : array_index_78981[1];
  assign array_update_78989[2] = add_78910 == 32'h0000_0002 ? add_78987 : array_index_78981[2];
  assign array_update_78989[3] = add_78910 == 32'h0000_0003 ? add_78987 : array_index_78981[3];
  assign array_update_78989[4] = add_78910 == 32'h0000_0004 ? add_78987 : array_index_78981[4];
  assign array_update_78989[5] = add_78910 == 32'h0000_0005 ? add_78987 : array_index_78981[5];
  assign array_update_78989[6] = add_78910 == 32'h0000_0006 ? add_78987 : array_index_78981[6];
  assign array_update_78989[7] = add_78910 == 32'h0000_0007 ? add_78987 : array_index_78981[7];
  assign array_update_78989[8] = add_78910 == 32'h0000_0008 ? add_78987 : array_index_78981[8];
  assign array_update_78989[9] = add_78910 == 32'h0000_0009 ? add_78987 : array_index_78981[9];
  assign add_78990 = add_78977 + 32'h0000_0001;
  assign array_update_78991[0] = add_78772 == 32'h0000_0000 ? array_update_78989 : array_update_78978[0];
  assign array_update_78991[1] = add_78772 == 32'h0000_0001 ? array_update_78989 : array_update_78978[1];
  assign array_update_78991[2] = add_78772 == 32'h0000_0002 ? array_update_78989 : array_update_78978[2];
  assign array_update_78991[3] = add_78772 == 32'h0000_0003 ? array_update_78989 : array_update_78978[3];
  assign array_update_78991[4] = add_78772 == 32'h0000_0004 ? array_update_78989 : array_update_78978[4];
  assign array_update_78991[5] = add_78772 == 32'h0000_0005 ? array_update_78989 : array_update_78978[5];
  assign array_update_78991[6] = add_78772 == 32'h0000_0006 ? array_update_78989 : array_update_78978[6];
  assign array_update_78991[7] = add_78772 == 32'h0000_0007 ? array_update_78989 : array_update_78978[7];
  assign array_update_78991[8] = add_78772 == 32'h0000_0008 ? array_update_78989 : array_update_78978[8];
  assign array_update_78991[9] = add_78772 == 32'h0000_0009 ? array_update_78989 : array_update_78978[9];
  assign array_index_78993 = array_update_72021[add_78990 > 32'h0000_0009 ? 4'h9 : add_78990[3:0]];
  assign array_index_78994 = array_update_78991[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_78998 = smul32b_32b_x_32b(array_index_78779[add_78990 > 32'h0000_0009 ? 4'h9 : add_78990[3:0]], array_index_78993[add_78910 > 32'h0000_0009 ? 4'h9 : add_78910[3:0]]);
  assign add_79000 = array_index_78994[add_78910 > 32'h0000_0009 ? 4'h9 : add_78910[3:0]] + smul_78998;
  assign array_update_79002[0] = add_78910 == 32'h0000_0000 ? add_79000 : array_index_78994[0];
  assign array_update_79002[1] = add_78910 == 32'h0000_0001 ? add_79000 : array_index_78994[1];
  assign array_update_79002[2] = add_78910 == 32'h0000_0002 ? add_79000 : array_index_78994[2];
  assign array_update_79002[3] = add_78910 == 32'h0000_0003 ? add_79000 : array_index_78994[3];
  assign array_update_79002[4] = add_78910 == 32'h0000_0004 ? add_79000 : array_index_78994[4];
  assign array_update_79002[5] = add_78910 == 32'h0000_0005 ? add_79000 : array_index_78994[5];
  assign array_update_79002[6] = add_78910 == 32'h0000_0006 ? add_79000 : array_index_78994[6];
  assign array_update_79002[7] = add_78910 == 32'h0000_0007 ? add_79000 : array_index_78994[7];
  assign array_update_79002[8] = add_78910 == 32'h0000_0008 ? add_79000 : array_index_78994[8];
  assign array_update_79002[9] = add_78910 == 32'h0000_0009 ? add_79000 : array_index_78994[9];
  assign add_79003 = add_78990 + 32'h0000_0001;
  assign array_update_79004[0] = add_78772 == 32'h0000_0000 ? array_update_79002 : array_update_78991[0];
  assign array_update_79004[1] = add_78772 == 32'h0000_0001 ? array_update_79002 : array_update_78991[1];
  assign array_update_79004[2] = add_78772 == 32'h0000_0002 ? array_update_79002 : array_update_78991[2];
  assign array_update_79004[3] = add_78772 == 32'h0000_0003 ? array_update_79002 : array_update_78991[3];
  assign array_update_79004[4] = add_78772 == 32'h0000_0004 ? array_update_79002 : array_update_78991[4];
  assign array_update_79004[5] = add_78772 == 32'h0000_0005 ? array_update_79002 : array_update_78991[5];
  assign array_update_79004[6] = add_78772 == 32'h0000_0006 ? array_update_79002 : array_update_78991[6];
  assign array_update_79004[7] = add_78772 == 32'h0000_0007 ? array_update_79002 : array_update_78991[7];
  assign array_update_79004[8] = add_78772 == 32'h0000_0008 ? array_update_79002 : array_update_78991[8];
  assign array_update_79004[9] = add_78772 == 32'h0000_0009 ? array_update_79002 : array_update_78991[9];
  assign array_index_79006 = array_update_72021[add_79003 > 32'h0000_0009 ? 4'h9 : add_79003[3:0]];
  assign array_index_79007 = array_update_79004[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_79011 = smul32b_32b_x_32b(array_index_78779[add_79003 > 32'h0000_0009 ? 4'h9 : add_79003[3:0]], array_index_79006[add_78910 > 32'h0000_0009 ? 4'h9 : add_78910[3:0]]);
  assign add_79013 = array_index_79007[add_78910 > 32'h0000_0009 ? 4'h9 : add_78910[3:0]] + smul_79011;
  assign array_update_79015[0] = add_78910 == 32'h0000_0000 ? add_79013 : array_index_79007[0];
  assign array_update_79015[1] = add_78910 == 32'h0000_0001 ? add_79013 : array_index_79007[1];
  assign array_update_79015[2] = add_78910 == 32'h0000_0002 ? add_79013 : array_index_79007[2];
  assign array_update_79015[3] = add_78910 == 32'h0000_0003 ? add_79013 : array_index_79007[3];
  assign array_update_79015[4] = add_78910 == 32'h0000_0004 ? add_79013 : array_index_79007[4];
  assign array_update_79015[5] = add_78910 == 32'h0000_0005 ? add_79013 : array_index_79007[5];
  assign array_update_79015[6] = add_78910 == 32'h0000_0006 ? add_79013 : array_index_79007[6];
  assign array_update_79015[7] = add_78910 == 32'h0000_0007 ? add_79013 : array_index_79007[7];
  assign array_update_79015[8] = add_78910 == 32'h0000_0008 ? add_79013 : array_index_79007[8];
  assign array_update_79015[9] = add_78910 == 32'h0000_0009 ? add_79013 : array_index_79007[9];
  assign add_79016 = add_79003 + 32'h0000_0001;
  assign array_update_79017[0] = add_78772 == 32'h0000_0000 ? array_update_79015 : array_update_79004[0];
  assign array_update_79017[1] = add_78772 == 32'h0000_0001 ? array_update_79015 : array_update_79004[1];
  assign array_update_79017[2] = add_78772 == 32'h0000_0002 ? array_update_79015 : array_update_79004[2];
  assign array_update_79017[3] = add_78772 == 32'h0000_0003 ? array_update_79015 : array_update_79004[3];
  assign array_update_79017[4] = add_78772 == 32'h0000_0004 ? array_update_79015 : array_update_79004[4];
  assign array_update_79017[5] = add_78772 == 32'h0000_0005 ? array_update_79015 : array_update_79004[5];
  assign array_update_79017[6] = add_78772 == 32'h0000_0006 ? array_update_79015 : array_update_79004[6];
  assign array_update_79017[7] = add_78772 == 32'h0000_0007 ? array_update_79015 : array_update_79004[7];
  assign array_update_79017[8] = add_78772 == 32'h0000_0008 ? array_update_79015 : array_update_79004[8];
  assign array_update_79017[9] = add_78772 == 32'h0000_0009 ? array_update_79015 : array_update_79004[9];
  assign array_index_79019 = array_update_72021[add_79016 > 32'h0000_0009 ? 4'h9 : add_79016[3:0]];
  assign array_index_79020 = array_update_79017[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_79024 = smul32b_32b_x_32b(array_index_78779[add_79016 > 32'h0000_0009 ? 4'h9 : add_79016[3:0]], array_index_79019[add_78910 > 32'h0000_0009 ? 4'h9 : add_78910[3:0]]);
  assign add_79026 = array_index_79020[add_78910 > 32'h0000_0009 ? 4'h9 : add_78910[3:0]] + smul_79024;
  assign array_update_79028[0] = add_78910 == 32'h0000_0000 ? add_79026 : array_index_79020[0];
  assign array_update_79028[1] = add_78910 == 32'h0000_0001 ? add_79026 : array_index_79020[1];
  assign array_update_79028[2] = add_78910 == 32'h0000_0002 ? add_79026 : array_index_79020[2];
  assign array_update_79028[3] = add_78910 == 32'h0000_0003 ? add_79026 : array_index_79020[3];
  assign array_update_79028[4] = add_78910 == 32'h0000_0004 ? add_79026 : array_index_79020[4];
  assign array_update_79028[5] = add_78910 == 32'h0000_0005 ? add_79026 : array_index_79020[5];
  assign array_update_79028[6] = add_78910 == 32'h0000_0006 ? add_79026 : array_index_79020[6];
  assign array_update_79028[7] = add_78910 == 32'h0000_0007 ? add_79026 : array_index_79020[7];
  assign array_update_79028[8] = add_78910 == 32'h0000_0008 ? add_79026 : array_index_79020[8];
  assign array_update_79028[9] = add_78910 == 32'h0000_0009 ? add_79026 : array_index_79020[9];
  assign add_79029 = add_79016 + 32'h0000_0001;
  assign array_update_79030[0] = add_78772 == 32'h0000_0000 ? array_update_79028 : array_update_79017[0];
  assign array_update_79030[1] = add_78772 == 32'h0000_0001 ? array_update_79028 : array_update_79017[1];
  assign array_update_79030[2] = add_78772 == 32'h0000_0002 ? array_update_79028 : array_update_79017[2];
  assign array_update_79030[3] = add_78772 == 32'h0000_0003 ? array_update_79028 : array_update_79017[3];
  assign array_update_79030[4] = add_78772 == 32'h0000_0004 ? array_update_79028 : array_update_79017[4];
  assign array_update_79030[5] = add_78772 == 32'h0000_0005 ? array_update_79028 : array_update_79017[5];
  assign array_update_79030[6] = add_78772 == 32'h0000_0006 ? array_update_79028 : array_update_79017[6];
  assign array_update_79030[7] = add_78772 == 32'h0000_0007 ? array_update_79028 : array_update_79017[7];
  assign array_update_79030[8] = add_78772 == 32'h0000_0008 ? array_update_79028 : array_update_79017[8];
  assign array_update_79030[9] = add_78772 == 32'h0000_0009 ? array_update_79028 : array_update_79017[9];
  assign array_index_79032 = array_update_72021[add_79029 > 32'h0000_0009 ? 4'h9 : add_79029[3:0]];
  assign array_index_79033 = array_update_79030[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_79037 = smul32b_32b_x_32b(array_index_78779[add_79029 > 32'h0000_0009 ? 4'h9 : add_79029[3:0]], array_index_79032[add_78910 > 32'h0000_0009 ? 4'h9 : add_78910[3:0]]);
  assign add_79039 = array_index_79033[add_78910 > 32'h0000_0009 ? 4'h9 : add_78910[3:0]] + smul_79037;
  assign array_update_79040[0] = add_78910 == 32'h0000_0000 ? add_79039 : array_index_79033[0];
  assign array_update_79040[1] = add_78910 == 32'h0000_0001 ? add_79039 : array_index_79033[1];
  assign array_update_79040[2] = add_78910 == 32'h0000_0002 ? add_79039 : array_index_79033[2];
  assign array_update_79040[3] = add_78910 == 32'h0000_0003 ? add_79039 : array_index_79033[3];
  assign array_update_79040[4] = add_78910 == 32'h0000_0004 ? add_79039 : array_index_79033[4];
  assign array_update_79040[5] = add_78910 == 32'h0000_0005 ? add_79039 : array_index_79033[5];
  assign array_update_79040[6] = add_78910 == 32'h0000_0006 ? add_79039 : array_index_79033[6];
  assign array_update_79040[7] = add_78910 == 32'h0000_0007 ? add_79039 : array_index_79033[7];
  assign array_update_79040[8] = add_78910 == 32'h0000_0008 ? add_79039 : array_index_79033[8];
  assign array_update_79040[9] = add_78910 == 32'h0000_0009 ? add_79039 : array_index_79033[9];
  assign array_update_79041[0] = add_78772 == 32'h0000_0000 ? array_update_79040 : array_update_79030[0];
  assign array_update_79041[1] = add_78772 == 32'h0000_0001 ? array_update_79040 : array_update_79030[1];
  assign array_update_79041[2] = add_78772 == 32'h0000_0002 ? array_update_79040 : array_update_79030[2];
  assign array_update_79041[3] = add_78772 == 32'h0000_0003 ? array_update_79040 : array_update_79030[3];
  assign array_update_79041[4] = add_78772 == 32'h0000_0004 ? array_update_79040 : array_update_79030[4];
  assign array_update_79041[5] = add_78772 == 32'h0000_0005 ? array_update_79040 : array_update_79030[5];
  assign array_update_79041[6] = add_78772 == 32'h0000_0006 ? array_update_79040 : array_update_79030[6];
  assign array_update_79041[7] = add_78772 == 32'h0000_0007 ? array_update_79040 : array_update_79030[7];
  assign array_update_79041[8] = add_78772 == 32'h0000_0008 ? array_update_79040 : array_update_79030[8];
  assign array_update_79041[9] = add_78772 == 32'h0000_0009 ? array_update_79040 : array_update_79030[9];
  assign array_index_79043 = array_update_79041[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign add_79045 = add_78910 + 32'h0000_0001;
  assign array_update_79046[0] = add_79045 == 32'h0000_0000 ? 32'h0000_0000 : array_index_79043[0];
  assign array_update_79046[1] = add_79045 == 32'h0000_0001 ? 32'h0000_0000 : array_index_79043[1];
  assign array_update_79046[2] = add_79045 == 32'h0000_0002 ? 32'h0000_0000 : array_index_79043[2];
  assign array_update_79046[3] = add_79045 == 32'h0000_0003 ? 32'h0000_0000 : array_index_79043[3];
  assign array_update_79046[4] = add_79045 == 32'h0000_0004 ? 32'h0000_0000 : array_index_79043[4];
  assign array_update_79046[5] = add_79045 == 32'h0000_0005 ? 32'h0000_0000 : array_index_79043[5];
  assign array_update_79046[6] = add_79045 == 32'h0000_0006 ? 32'h0000_0000 : array_index_79043[6];
  assign array_update_79046[7] = add_79045 == 32'h0000_0007 ? 32'h0000_0000 : array_index_79043[7];
  assign array_update_79046[8] = add_79045 == 32'h0000_0008 ? 32'h0000_0000 : array_index_79043[8];
  assign array_update_79046[9] = add_79045 == 32'h0000_0009 ? 32'h0000_0000 : array_index_79043[9];
  assign literal_79047 = 32'h0000_0000;
  assign array_update_79048[0] = add_78772 == 32'h0000_0000 ? array_update_79046 : array_update_79041[0];
  assign array_update_79048[1] = add_78772 == 32'h0000_0001 ? array_update_79046 : array_update_79041[1];
  assign array_update_79048[2] = add_78772 == 32'h0000_0002 ? array_update_79046 : array_update_79041[2];
  assign array_update_79048[3] = add_78772 == 32'h0000_0003 ? array_update_79046 : array_update_79041[3];
  assign array_update_79048[4] = add_78772 == 32'h0000_0004 ? array_update_79046 : array_update_79041[4];
  assign array_update_79048[5] = add_78772 == 32'h0000_0005 ? array_update_79046 : array_update_79041[5];
  assign array_update_79048[6] = add_78772 == 32'h0000_0006 ? array_update_79046 : array_update_79041[6];
  assign array_update_79048[7] = add_78772 == 32'h0000_0007 ? array_update_79046 : array_update_79041[7];
  assign array_update_79048[8] = add_78772 == 32'h0000_0008 ? array_update_79046 : array_update_79041[8];
  assign array_update_79048[9] = add_78772 == 32'h0000_0009 ? array_update_79046 : array_update_79041[9];
  assign array_index_79050 = array_update_72021[literal_79047 > 32'h0000_0009 ? 4'h9 : literal_79047[3:0]];
  assign array_index_79051 = array_update_79048[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_79055 = smul32b_32b_x_32b(array_index_78779[literal_79047 > 32'h0000_0009 ? 4'h9 : literal_79047[3:0]], array_index_79050[add_79045 > 32'h0000_0009 ? 4'h9 : add_79045[3:0]]);
  assign add_79057 = array_index_79051[add_79045 > 32'h0000_0009 ? 4'h9 : add_79045[3:0]] + smul_79055;
  assign array_update_79059[0] = add_79045 == 32'h0000_0000 ? add_79057 : array_index_79051[0];
  assign array_update_79059[1] = add_79045 == 32'h0000_0001 ? add_79057 : array_index_79051[1];
  assign array_update_79059[2] = add_79045 == 32'h0000_0002 ? add_79057 : array_index_79051[2];
  assign array_update_79059[3] = add_79045 == 32'h0000_0003 ? add_79057 : array_index_79051[3];
  assign array_update_79059[4] = add_79045 == 32'h0000_0004 ? add_79057 : array_index_79051[4];
  assign array_update_79059[5] = add_79045 == 32'h0000_0005 ? add_79057 : array_index_79051[5];
  assign array_update_79059[6] = add_79045 == 32'h0000_0006 ? add_79057 : array_index_79051[6];
  assign array_update_79059[7] = add_79045 == 32'h0000_0007 ? add_79057 : array_index_79051[7];
  assign array_update_79059[8] = add_79045 == 32'h0000_0008 ? add_79057 : array_index_79051[8];
  assign array_update_79059[9] = add_79045 == 32'h0000_0009 ? add_79057 : array_index_79051[9];
  assign add_79060 = literal_79047 + 32'h0000_0001;
  assign array_update_79061[0] = add_78772 == 32'h0000_0000 ? array_update_79059 : array_update_79048[0];
  assign array_update_79061[1] = add_78772 == 32'h0000_0001 ? array_update_79059 : array_update_79048[1];
  assign array_update_79061[2] = add_78772 == 32'h0000_0002 ? array_update_79059 : array_update_79048[2];
  assign array_update_79061[3] = add_78772 == 32'h0000_0003 ? array_update_79059 : array_update_79048[3];
  assign array_update_79061[4] = add_78772 == 32'h0000_0004 ? array_update_79059 : array_update_79048[4];
  assign array_update_79061[5] = add_78772 == 32'h0000_0005 ? array_update_79059 : array_update_79048[5];
  assign array_update_79061[6] = add_78772 == 32'h0000_0006 ? array_update_79059 : array_update_79048[6];
  assign array_update_79061[7] = add_78772 == 32'h0000_0007 ? array_update_79059 : array_update_79048[7];
  assign array_update_79061[8] = add_78772 == 32'h0000_0008 ? array_update_79059 : array_update_79048[8];
  assign array_update_79061[9] = add_78772 == 32'h0000_0009 ? array_update_79059 : array_update_79048[9];
  assign array_index_79063 = array_update_72021[add_79060 > 32'h0000_0009 ? 4'h9 : add_79060[3:0]];
  assign array_index_79064 = array_update_79061[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_79068 = smul32b_32b_x_32b(array_index_78779[add_79060 > 32'h0000_0009 ? 4'h9 : add_79060[3:0]], array_index_79063[add_79045 > 32'h0000_0009 ? 4'h9 : add_79045[3:0]]);
  assign add_79070 = array_index_79064[add_79045 > 32'h0000_0009 ? 4'h9 : add_79045[3:0]] + smul_79068;
  assign array_update_79072[0] = add_79045 == 32'h0000_0000 ? add_79070 : array_index_79064[0];
  assign array_update_79072[1] = add_79045 == 32'h0000_0001 ? add_79070 : array_index_79064[1];
  assign array_update_79072[2] = add_79045 == 32'h0000_0002 ? add_79070 : array_index_79064[2];
  assign array_update_79072[3] = add_79045 == 32'h0000_0003 ? add_79070 : array_index_79064[3];
  assign array_update_79072[4] = add_79045 == 32'h0000_0004 ? add_79070 : array_index_79064[4];
  assign array_update_79072[5] = add_79045 == 32'h0000_0005 ? add_79070 : array_index_79064[5];
  assign array_update_79072[6] = add_79045 == 32'h0000_0006 ? add_79070 : array_index_79064[6];
  assign array_update_79072[7] = add_79045 == 32'h0000_0007 ? add_79070 : array_index_79064[7];
  assign array_update_79072[8] = add_79045 == 32'h0000_0008 ? add_79070 : array_index_79064[8];
  assign array_update_79072[9] = add_79045 == 32'h0000_0009 ? add_79070 : array_index_79064[9];
  assign add_79073 = add_79060 + 32'h0000_0001;
  assign array_update_79074[0] = add_78772 == 32'h0000_0000 ? array_update_79072 : array_update_79061[0];
  assign array_update_79074[1] = add_78772 == 32'h0000_0001 ? array_update_79072 : array_update_79061[1];
  assign array_update_79074[2] = add_78772 == 32'h0000_0002 ? array_update_79072 : array_update_79061[2];
  assign array_update_79074[3] = add_78772 == 32'h0000_0003 ? array_update_79072 : array_update_79061[3];
  assign array_update_79074[4] = add_78772 == 32'h0000_0004 ? array_update_79072 : array_update_79061[4];
  assign array_update_79074[5] = add_78772 == 32'h0000_0005 ? array_update_79072 : array_update_79061[5];
  assign array_update_79074[6] = add_78772 == 32'h0000_0006 ? array_update_79072 : array_update_79061[6];
  assign array_update_79074[7] = add_78772 == 32'h0000_0007 ? array_update_79072 : array_update_79061[7];
  assign array_update_79074[8] = add_78772 == 32'h0000_0008 ? array_update_79072 : array_update_79061[8];
  assign array_update_79074[9] = add_78772 == 32'h0000_0009 ? array_update_79072 : array_update_79061[9];
  assign array_index_79076 = array_update_72021[add_79073 > 32'h0000_0009 ? 4'h9 : add_79073[3:0]];
  assign array_index_79077 = array_update_79074[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_79081 = smul32b_32b_x_32b(array_index_78779[add_79073 > 32'h0000_0009 ? 4'h9 : add_79073[3:0]], array_index_79076[add_79045 > 32'h0000_0009 ? 4'h9 : add_79045[3:0]]);
  assign add_79083 = array_index_79077[add_79045 > 32'h0000_0009 ? 4'h9 : add_79045[3:0]] + smul_79081;
  assign array_update_79085[0] = add_79045 == 32'h0000_0000 ? add_79083 : array_index_79077[0];
  assign array_update_79085[1] = add_79045 == 32'h0000_0001 ? add_79083 : array_index_79077[1];
  assign array_update_79085[2] = add_79045 == 32'h0000_0002 ? add_79083 : array_index_79077[2];
  assign array_update_79085[3] = add_79045 == 32'h0000_0003 ? add_79083 : array_index_79077[3];
  assign array_update_79085[4] = add_79045 == 32'h0000_0004 ? add_79083 : array_index_79077[4];
  assign array_update_79085[5] = add_79045 == 32'h0000_0005 ? add_79083 : array_index_79077[5];
  assign array_update_79085[6] = add_79045 == 32'h0000_0006 ? add_79083 : array_index_79077[6];
  assign array_update_79085[7] = add_79045 == 32'h0000_0007 ? add_79083 : array_index_79077[7];
  assign array_update_79085[8] = add_79045 == 32'h0000_0008 ? add_79083 : array_index_79077[8];
  assign array_update_79085[9] = add_79045 == 32'h0000_0009 ? add_79083 : array_index_79077[9];
  assign add_79086 = add_79073 + 32'h0000_0001;
  assign array_update_79087[0] = add_78772 == 32'h0000_0000 ? array_update_79085 : array_update_79074[0];
  assign array_update_79087[1] = add_78772 == 32'h0000_0001 ? array_update_79085 : array_update_79074[1];
  assign array_update_79087[2] = add_78772 == 32'h0000_0002 ? array_update_79085 : array_update_79074[2];
  assign array_update_79087[3] = add_78772 == 32'h0000_0003 ? array_update_79085 : array_update_79074[3];
  assign array_update_79087[4] = add_78772 == 32'h0000_0004 ? array_update_79085 : array_update_79074[4];
  assign array_update_79087[5] = add_78772 == 32'h0000_0005 ? array_update_79085 : array_update_79074[5];
  assign array_update_79087[6] = add_78772 == 32'h0000_0006 ? array_update_79085 : array_update_79074[6];
  assign array_update_79087[7] = add_78772 == 32'h0000_0007 ? array_update_79085 : array_update_79074[7];
  assign array_update_79087[8] = add_78772 == 32'h0000_0008 ? array_update_79085 : array_update_79074[8];
  assign array_update_79087[9] = add_78772 == 32'h0000_0009 ? array_update_79085 : array_update_79074[9];
  assign array_index_79089 = array_update_72021[add_79086 > 32'h0000_0009 ? 4'h9 : add_79086[3:0]];
  assign array_index_79090 = array_update_79087[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_79094 = smul32b_32b_x_32b(array_index_78779[add_79086 > 32'h0000_0009 ? 4'h9 : add_79086[3:0]], array_index_79089[add_79045 > 32'h0000_0009 ? 4'h9 : add_79045[3:0]]);
  assign add_79096 = array_index_79090[add_79045 > 32'h0000_0009 ? 4'h9 : add_79045[3:0]] + smul_79094;
  assign array_update_79098[0] = add_79045 == 32'h0000_0000 ? add_79096 : array_index_79090[0];
  assign array_update_79098[1] = add_79045 == 32'h0000_0001 ? add_79096 : array_index_79090[1];
  assign array_update_79098[2] = add_79045 == 32'h0000_0002 ? add_79096 : array_index_79090[2];
  assign array_update_79098[3] = add_79045 == 32'h0000_0003 ? add_79096 : array_index_79090[3];
  assign array_update_79098[4] = add_79045 == 32'h0000_0004 ? add_79096 : array_index_79090[4];
  assign array_update_79098[5] = add_79045 == 32'h0000_0005 ? add_79096 : array_index_79090[5];
  assign array_update_79098[6] = add_79045 == 32'h0000_0006 ? add_79096 : array_index_79090[6];
  assign array_update_79098[7] = add_79045 == 32'h0000_0007 ? add_79096 : array_index_79090[7];
  assign array_update_79098[8] = add_79045 == 32'h0000_0008 ? add_79096 : array_index_79090[8];
  assign array_update_79098[9] = add_79045 == 32'h0000_0009 ? add_79096 : array_index_79090[9];
  assign add_79099 = add_79086 + 32'h0000_0001;
  assign array_update_79100[0] = add_78772 == 32'h0000_0000 ? array_update_79098 : array_update_79087[0];
  assign array_update_79100[1] = add_78772 == 32'h0000_0001 ? array_update_79098 : array_update_79087[1];
  assign array_update_79100[2] = add_78772 == 32'h0000_0002 ? array_update_79098 : array_update_79087[2];
  assign array_update_79100[3] = add_78772 == 32'h0000_0003 ? array_update_79098 : array_update_79087[3];
  assign array_update_79100[4] = add_78772 == 32'h0000_0004 ? array_update_79098 : array_update_79087[4];
  assign array_update_79100[5] = add_78772 == 32'h0000_0005 ? array_update_79098 : array_update_79087[5];
  assign array_update_79100[6] = add_78772 == 32'h0000_0006 ? array_update_79098 : array_update_79087[6];
  assign array_update_79100[7] = add_78772 == 32'h0000_0007 ? array_update_79098 : array_update_79087[7];
  assign array_update_79100[8] = add_78772 == 32'h0000_0008 ? array_update_79098 : array_update_79087[8];
  assign array_update_79100[9] = add_78772 == 32'h0000_0009 ? array_update_79098 : array_update_79087[9];
  assign array_index_79102 = array_update_72021[add_79099 > 32'h0000_0009 ? 4'h9 : add_79099[3:0]];
  assign array_index_79103 = array_update_79100[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_79107 = smul32b_32b_x_32b(array_index_78779[add_79099 > 32'h0000_0009 ? 4'h9 : add_79099[3:0]], array_index_79102[add_79045 > 32'h0000_0009 ? 4'h9 : add_79045[3:0]]);
  assign add_79109 = array_index_79103[add_79045 > 32'h0000_0009 ? 4'h9 : add_79045[3:0]] + smul_79107;
  assign array_update_79111[0] = add_79045 == 32'h0000_0000 ? add_79109 : array_index_79103[0];
  assign array_update_79111[1] = add_79045 == 32'h0000_0001 ? add_79109 : array_index_79103[1];
  assign array_update_79111[2] = add_79045 == 32'h0000_0002 ? add_79109 : array_index_79103[2];
  assign array_update_79111[3] = add_79045 == 32'h0000_0003 ? add_79109 : array_index_79103[3];
  assign array_update_79111[4] = add_79045 == 32'h0000_0004 ? add_79109 : array_index_79103[4];
  assign array_update_79111[5] = add_79045 == 32'h0000_0005 ? add_79109 : array_index_79103[5];
  assign array_update_79111[6] = add_79045 == 32'h0000_0006 ? add_79109 : array_index_79103[6];
  assign array_update_79111[7] = add_79045 == 32'h0000_0007 ? add_79109 : array_index_79103[7];
  assign array_update_79111[8] = add_79045 == 32'h0000_0008 ? add_79109 : array_index_79103[8];
  assign array_update_79111[9] = add_79045 == 32'h0000_0009 ? add_79109 : array_index_79103[9];
  assign add_79112 = add_79099 + 32'h0000_0001;
  assign array_update_79113[0] = add_78772 == 32'h0000_0000 ? array_update_79111 : array_update_79100[0];
  assign array_update_79113[1] = add_78772 == 32'h0000_0001 ? array_update_79111 : array_update_79100[1];
  assign array_update_79113[2] = add_78772 == 32'h0000_0002 ? array_update_79111 : array_update_79100[2];
  assign array_update_79113[3] = add_78772 == 32'h0000_0003 ? array_update_79111 : array_update_79100[3];
  assign array_update_79113[4] = add_78772 == 32'h0000_0004 ? array_update_79111 : array_update_79100[4];
  assign array_update_79113[5] = add_78772 == 32'h0000_0005 ? array_update_79111 : array_update_79100[5];
  assign array_update_79113[6] = add_78772 == 32'h0000_0006 ? array_update_79111 : array_update_79100[6];
  assign array_update_79113[7] = add_78772 == 32'h0000_0007 ? array_update_79111 : array_update_79100[7];
  assign array_update_79113[8] = add_78772 == 32'h0000_0008 ? array_update_79111 : array_update_79100[8];
  assign array_update_79113[9] = add_78772 == 32'h0000_0009 ? array_update_79111 : array_update_79100[9];
  assign array_index_79115 = array_update_72021[add_79112 > 32'h0000_0009 ? 4'h9 : add_79112[3:0]];
  assign array_index_79116 = array_update_79113[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_79120 = smul32b_32b_x_32b(array_index_78779[add_79112 > 32'h0000_0009 ? 4'h9 : add_79112[3:0]], array_index_79115[add_79045 > 32'h0000_0009 ? 4'h9 : add_79045[3:0]]);
  assign add_79122 = array_index_79116[add_79045 > 32'h0000_0009 ? 4'h9 : add_79045[3:0]] + smul_79120;
  assign array_update_79124[0] = add_79045 == 32'h0000_0000 ? add_79122 : array_index_79116[0];
  assign array_update_79124[1] = add_79045 == 32'h0000_0001 ? add_79122 : array_index_79116[1];
  assign array_update_79124[2] = add_79045 == 32'h0000_0002 ? add_79122 : array_index_79116[2];
  assign array_update_79124[3] = add_79045 == 32'h0000_0003 ? add_79122 : array_index_79116[3];
  assign array_update_79124[4] = add_79045 == 32'h0000_0004 ? add_79122 : array_index_79116[4];
  assign array_update_79124[5] = add_79045 == 32'h0000_0005 ? add_79122 : array_index_79116[5];
  assign array_update_79124[6] = add_79045 == 32'h0000_0006 ? add_79122 : array_index_79116[6];
  assign array_update_79124[7] = add_79045 == 32'h0000_0007 ? add_79122 : array_index_79116[7];
  assign array_update_79124[8] = add_79045 == 32'h0000_0008 ? add_79122 : array_index_79116[8];
  assign array_update_79124[9] = add_79045 == 32'h0000_0009 ? add_79122 : array_index_79116[9];
  assign add_79125 = add_79112 + 32'h0000_0001;
  assign array_update_79126[0] = add_78772 == 32'h0000_0000 ? array_update_79124 : array_update_79113[0];
  assign array_update_79126[1] = add_78772 == 32'h0000_0001 ? array_update_79124 : array_update_79113[1];
  assign array_update_79126[2] = add_78772 == 32'h0000_0002 ? array_update_79124 : array_update_79113[2];
  assign array_update_79126[3] = add_78772 == 32'h0000_0003 ? array_update_79124 : array_update_79113[3];
  assign array_update_79126[4] = add_78772 == 32'h0000_0004 ? array_update_79124 : array_update_79113[4];
  assign array_update_79126[5] = add_78772 == 32'h0000_0005 ? array_update_79124 : array_update_79113[5];
  assign array_update_79126[6] = add_78772 == 32'h0000_0006 ? array_update_79124 : array_update_79113[6];
  assign array_update_79126[7] = add_78772 == 32'h0000_0007 ? array_update_79124 : array_update_79113[7];
  assign array_update_79126[8] = add_78772 == 32'h0000_0008 ? array_update_79124 : array_update_79113[8];
  assign array_update_79126[9] = add_78772 == 32'h0000_0009 ? array_update_79124 : array_update_79113[9];
  assign array_index_79128 = array_update_72021[add_79125 > 32'h0000_0009 ? 4'h9 : add_79125[3:0]];
  assign array_index_79129 = array_update_79126[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_79133 = smul32b_32b_x_32b(array_index_78779[add_79125 > 32'h0000_0009 ? 4'h9 : add_79125[3:0]], array_index_79128[add_79045 > 32'h0000_0009 ? 4'h9 : add_79045[3:0]]);
  assign add_79135 = array_index_79129[add_79045 > 32'h0000_0009 ? 4'h9 : add_79045[3:0]] + smul_79133;
  assign array_update_79137[0] = add_79045 == 32'h0000_0000 ? add_79135 : array_index_79129[0];
  assign array_update_79137[1] = add_79045 == 32'h0000_0001 ? add_79135 : array_index_79129[1];
  assign array_update_79137[2] = add_79045 == 32'h0000_0002 ? add_79135 : array_index_79129[2];
  assign array_update_79137[3] = add_79045 == 32'h0000_0003 ? add_79135 : array_index_79129[3];
  assign array_update_79137[4] = add_79045 == 32'h0000_0004 ? add_79135 : array_index_79129[4];
  assign array_update_79137[5] = add_79045 == 32'h0000_0005 ? add_79135 : array_index_79129[5];
  assign array_update_79137[6] = add_79045 == 32'h0000_0006 ? add_79135 : array_index_79129[6];
  assign array_update_79137[7] = add_79045 == 32'h0000_0007 ? add_79135 : array_index_79129[7];
  assign array_update_79137[8] = add_79045 == 32'h0000_0008 ? add_79135 : array_index_79129[8];
  assign array_update_79137[9] = add_79045 == 32'h0000_0009 ? add_79135 : array_index_79129[9];
  assign add_79138 = add_79125 + 32'h0000_0001;
  assign array_update_79139[0] = add_78772 == 32'h0000_0000 ? array_update_79137 : array_update_79126[0];
  assign array_update_79139[1] = add_78772 == 32'h0000_0001 ? array_update_79137 : array_update_79126[1];
  assign array_update_79139[2] = add_78772 == 32'h0000_0002 ? array_update_79137 : array_update_79126[2];
  assign array_update_79139[3] = add_78772 == 32'h0000_0003 ? array_update_79137 : array_update_79126[3];
  assign array_update_79139[4] = add_78772 == 32'h0000_0004 ? array_update_79137 : array_update_79126[4];
  assign array_update_79139[5] = add_78772 == 32'h0000_0005 ? array_update_79137 : array_update_79126[5];
  assign array_update_79139[6] = add_78772 == 32'h0000_0006 ? array_update_79137 : array_update_79126[6];
  assign array_update_79139[7] = add_78772 == 32'h0000_0007 ? array_update_79137 : array_update_79126[7];
  assign array_update_79139[8] = add_78772 == 32'h0000_0008 ? array_update_79137 : array_update_79126[8];
  assign array_update_79139[9] = add_78772 == 32'h0000_0009 ? array_update_79137 : array_update_79126[9];
  assign array_index_79141 = array_update_72021[add_79138 > 32'h0000_0009 ? 4'h9 : add_79138[3:0]];
  assign array_index_79142 = array_update_79139[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_79146 = smul32b_32b_x_32b(array_index_78779[add_79138 > 32'h0000_0009 ? 4'h9 : add_79138[3:0]], array_index_79141[add_79045 > 32'h0000_0009 ? 4'h9 : add_79045[3:0]]);
  assign add_79148 = array_index_79142[add_79045 > 32'h0000_0009 ? 4'h9 : add_79045[3:0]] + smul_79146;
  assign array_update_79150[0] = add_79045 == 32'h0000_0000 ? add_79148 : array_index_79142[0];
  assign array_update_79150[1] = add_79045 == 32'h0000_0001 ? add_79148 : array_index_79142[1];
  assign array_update_79150[2] = add_79045 == 32'h0000_0002 ? add_79148 : array_index_79142[2];
  assign array_update_79150[3] = add_79045 == 32'h0000_0003 ? add_79148 : array_index_79142[3];
  assign array_update_79150[4] = add_79045 == 32'h0000_0004 ? add_79148 : array_index_79142[4];
  assign array_update_79150[5] = add_79045 == 32'h0000_0005 ? add_79148 : array_index_79142[5];
  assign array_update_79150[6] = add_79045 == 32'h0000_0006 ? add_79148 : array_index_79142[6];
  assign array_update_79150[7] = add_79045 == 32'h0000_0007 ? add_79148 : array_index_79142[7];
  assign array_update_79150[8] = add_79045 == 32'h0000_0008 ? add_79148 : array_index_79142[8];
  assign array_update_79150[9] = add_79045 == 32'h0000_0009 ? add_79148 : array_index_79142[9];
  assign add_79151 = add_79138 + 32'h0000_0001;
  assign array_update_79152[0] = add_78772 == 32'h0000_0000 ? array_update_79150 : array_update_79139[0];
  assign array_update_79152[1] = add_78772 == 32'h0000_0001 ? array_update_79150 : array_update_79139[1];
  assign array_update_79152[2] = add_78772 == 32'h0000_0002 ? array_update_79150 : array_update_79139[2];
  assign array_update_79152[3] = add_78772 == 32'h0000_0003 ? array_update_79150 : array_update_79139[3];
  assign array_update_79152[4] = add_78772 == 32'h0000_0004 ? array_update_79150 : array_update_79139[4];
  assign array_update_79152[5] = add_78772 == 32'h0000_0005 ? array_update_79150 : array_update_79139[5];
  assign array_update_79152[6] = add_78772 == 32'h0000_0006 ? array_update_79150 : array_update_79139[6];
  assign array_update_79152[7] = add_78772 == 32'h0000_0007 ? array_update_79150 : array_update_79139[7];
  assign array_update_79152[8] = add_78772 == 32'h0000_0008 ? array_update_79150 : array_update_79139[8];
  assign array_update_79152[9] = add_78772 == 32'h0000_0009 ? array_update_79150 : array_update_79139[9];
  assign array_index_79154 = array_update_72021[add_79151 > 32'h0000_0009 ? 4'h9 : add_79151[3:0]];
  assign array_index_79155 = array_update_79152[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_79159 = smul32b_32b_x_32b(array_index_78779[add_79151 > 32'h0000_0009 ? 4'h9 : add_79151[3:0]], array_index_79154[add_79045 > 32'h0000_0009 ? 4'h9 : add_79045[3:0]]);
  assign add_79161 = array_index_79155[add_79045 > 32'h0000_0009 ? 4'h9 : add_79045[3:0]] + smul_79159;
  assign array_update_79163[0] = add_79045 == 32'h0000_0000 ? add_79161 : array_index_79155[0];
  assign array_update_79163[1] = add_79045 == 32'h0000_0001 ? add_79161 : array_index_79155[1];
  assign array_update_79163[2] = add_79045 == 32'h0000_0002 ? add_79161 : array_index_79155[2];
  assign array_update_79163[3] = add_79045 == 32'h0000_0003 ? add_79161 : array_index_79155[3];
  assign array_update_79163[4] = add_79045 == 32'h0000_0004 ? add_79161 : array_index_79155[4];
  assign array_update_79163[5] = add_79045 == 32'h0000_0005 ? add_79161 : array_index_79155[5];
  assign array_update_79163[6] = add_79045 == 32'h0000_0006 ? add_79161 : array_index_79155[6];
  assign array_update_79163[7] = add_79045 == 32'h0000_0007 ? add_79161 : array_index_79155[7];
  assign array_update_79163[8] = add_79045 == 32'h0000_0008 ? add_79161 : array_index_79155[8];
  assign array_update_79163[9] = add_79045 == 32'h0000_0009 ? add_79161 : array_index_79155[9];
  assign add_79164 = add_79151 + 32'h0000_0001;
  assign array_update_79165[0] = add_78772 == 32'h0000_0000 ? array_update_79163 : array_update_79152[0];
  assign array_update_79165[1] = add_78772 == 32'h0000_0001 ? array_update_79163 : array_update_79152[1];
  assign array_update_79165[2] = add_78772 == 32'h0000_0002 ? array_update_79163 : array_update_79152[2];
  assign array_update_79165[3] = add_78772 == 32'h0000_0003 ? array_update_79163 : array_update_79152[3];
  assign array_update_79165[4] = add_78772 == 32'h0000_0004 ? array_update_79163 : array_update_79152[4];
  assign array_update_79165[5] = add_78772 == 32'h0000_0005 ? array_update_79163 : array_update_79152[5];
  assign array_update_79165[6] = add_78772 == 32'h0000_0006 ? array_update_79163 : array_update_79152[6];
  assign array_update_79165[7] = add_78772 == 32'h0000_0007 ? array_update_79163 : array_update_79152[7];
  assign array_update_79165[8] = add_78772 == 32'h0000_0008 ? array_update_79163 : array_update_79152[8];
  assign array_update_79165[9] = add_78772 == 32'h0000_0009 ? array_update_79163 : array_update_79152[9];
  assign array_index_79167 = array_update_72021[add_79164 > 32'h0000_0009 ? 4'h9 : add_79164[3:0]];
  assign array_index_79168 = array_update_79165[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_79172 = smul32b_32b_x_32b(array_index_78779[add_79164 > 32'h0000_0009 ? 4'h9 : add_79164[3:0]], array_index_79167[add_79045 > 32'h0000_0009 ? 4'h9 : add_79045[3:0]]);
  assign add_79174 = array_index_79168[add_79045 > 32'h0000_0009 ? 4'h9 : add_79045[3:0]] + smul_79172;
  assign array_update_79175[0] = add_79045 == 32'h0000_0000 ? add_79174 : array_index_79168[0];
  assign array_update_79175[1] = add_79045 == 32'h0000_0001 ? add_79174 : array_index_79168[1];
  assign array_update_79175[2] = add_79045 == 32'h0000_0002 ? add_79174 : array_index_79168[2];
  assign array_update_79175[3] = add_79045 == 32'h0000_0003 ? add_79174 : array_index_79168[3];
  assign array_update_79175[4] = add_79045 == 32'h0000_0004 ? add_79174 : array_index_79168[4];
  assign array_update_79175[5] = add_79045 == 32'h0000_0005 ? add_79174 : array_index_79168[5];
  assign array_update_79175[6] = add_79045 == 32'h0000_0006 ? add_79174 : array_index_79168[6];
  assign array_update_79175[7] = add_79045 == 32'h0000_0007 ? add_79174 : array_index_79168[7];
  assign array_update_79175[8] = add_79045 == 32'h0000_0008 ? add_79174 : array_index_79168[8];
  assign array_update_79175[9] = add_79045 == 32'h0000_0009 ? add_79174 : array_index_79168[9];
  assign array_update_79176[0] = add_78772 == 32'h0000_0000 ? array_update_79175 : array_update_79165[0];
  assign array_update_79176[1] = add_78772 == 32'h0000_0001 ? array_update_79175 : array_update_79165[1];
  assign array_update_79176[2] = add_78772 == 32'h0000_0002 ? array_update_79175 : array_update_79165[2];
  assign array_update_79176[3] = add_78772 == 32'h0000_0003 ? array_update_79175 : array_update_79165[3];
  assign array_update_79176[4] = add_78772 == 32'h0000_0004 ? array_update_79175 : array_update_79165[4];
  assign array_update_79176[5] = add_78772 == 32'h0000_0005 ? array_update_79175 : array_update_79165[5];
  assign array_update_79176[6] = add_78772 == 32'h0000_0006 ? array_update_79175 : array_update_79165[6];
  assign array_update_79176[7] = add_78772 == 32'h0000_0007 ? array_update_79175 : array_update_79165[7];
  assign array_update_79176[8] = add_78772 == 32'h0000_0008 ? array_update_79175 : array_update_79165[8];
  assign array_update_79176[9] = add_78772 == 32'h0000_0009 ? array_update_79175 : array_update_79165[9];
  assign array_index_79178 = array_update_79176[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign add_79180 = add_79045 + 32'h0000_0001;
  assign array_update_79181[0] = add_79180 == 32'h0000_0000 ? 32'h0000_0000 : array_index_79178[0];
  assign array_update_79181[1] = add_79180 == 32'h0000_0001 ? 32'h0000_0000 : array_index_79178[1];
  assign array_update_79181[2] = add_79180 == 32'h0000_0002 ? 32'h0000_0000 : array_index_79178[2];
  assign array_update_79181[3] = add_79180 == 32'h0000_0003 ? 32'h0000_0000 : array_index_79178[3];
  assign array_update_79181[4] = add_79180 == 32'h0000_0004 ? 32'h0000_0000 : array_index_79178[4];
  assign array_update_79181[5] = add_79180 == 32'h0000_0005 ? 32'h0000_0000 : array_index_79178[5];
  assign array_update_79181[6] = add_79180 == 32'h0000_0006 ? 32'h0000_0000 : array_index_79178[6];
  assign array_update_79181[7] = add_79180 == 32'h0000_0007 ? 32'h0000_0000 : array_index_79178[7];
  assign array_update_79181[8] = add_79180 == 32'h0000_0008 ? 32'h0000_0000 : array_index_79178[8];
  assign array_update_79181[9] = add_79180 == 32'h0000_0009 ? 32'h0000_0000 : array_index_79178[9];
  assign literal_79182 = 32'h0000_0000;
  assign array_update_79183[0] = add_78772 == 32'h0000_0000 ? array_update_79181 : array_update_79176[0];
  assign array_update_79183[1] = add_78772 == 32'h0000_0001 ? array_update_79181 : array_update_79176[1];
  assign array_update_79183[2] = add_78772 == 32'h0000_0002 ? array_update_79181 : array_update_79176[2];
  assign array_update_79183[3] = add_78772 == 32'h0000_0003 ? array_update_79181 : array_update_79176[3];
  assign array_update_79183[4] = add_78772 == 32'h0000_0004 ? array_update_79181 : array_update_79176[4];
  assign array_update_79183[5] = add_78772 == 32'h0000_0005 ? array_update_79181 : array_update_79176[5];
  assign array_update_79183[6] = add_78772 == 32'h0000_0006 ? array_update_79181 : array_update_79176[6];
  assign array_update_79183[7] = add_78772 == 32'h0000_0007 ? array_update_79181 : array_update_79176[7];
  assign array_update_79183[8] = add_78772 == 32'h0000_0008 ? array_update_79181 : array_update_79176[8];
  assign array_update_79183[9] = add_78772 == 32'h0000_0009 ? array_update_79181 : array_update_79176[9];
  assign array_index_79185 = array_update_72021[literal_79182 > 32'h0000_0009 ? 4'h9 : literal_79182[3:0]];
  assign array_index_79186 = array_update_79183[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_79190 = smul32b_32b_x_32b(array_index_78779[literal_79182 > 32'h0000_0009 ? 4'h9 : literal_79182[3:0]], array_index_79185[add_79180 > 32'h0000_0009 ? 4'h9 : add_79180[3:0]]);
  assign add_79192 = array_index_79186[add_79180 > 32'h0000_0009 ? 4'h9 : add_79180[3:0]] + smul_79190;
  assign array_update_79194[0] = add_79180 == 32'h0000_0000 ? add_79192 : array_index_79186[0];
  assign array_update_79194[1] = add_79180 == 32'h0000_0001 ? add_79192 : array_index_79186[1];
  assign array_update_79194[2] = add_79180 == 32'h0000_0002 ? add_79192 : array_index_79186[2];
  assign array_update_79194[3] = add_79180 == 32'h0000_0003 ? add_79192 : array_index_79186[3];
  assign array_update_79194[4] = add_79180 == 32'h0000_0004 ? add_79192 : array_index_79186[4];
  assign array_update_79194[5] = add_79180 == 32'h0000_0005 ? add_79192 : array_index_79186[5];
  assign array_update_79194[6] = add_79180 == 32'h0000_0006 ? add_79192 : array_index_79186[6];
  assign array_update_79194[7] = add_79180 == 32'h0000_0007 ? add_79192 : array_index_79186[7];
  assign array_update_79194[8] = add_79180 == 32'h0000_0008 ? add_79192 : array_index_79186[8];
  assign array_update_79194[9] = add_79180 == 32'h0000_0009 ? add_79192 : array_index_79186[9];
  assign add_79195 = literal_79182 + 32'h0000_0001;
  assign array_update_79196[0] = add_78772 == 32'h0000_0000 ? array_update_79194 : array_update_79183[0];
  assign array_update_79196[1] = add_78772 == 32'h0000_0001 ? array_update_79194 : array_update_79183[1];
  assign array_update_79196[2] = add_78772 == 32'h0000_0002 ? array_update_79194 : array_update_79183[2];
  assign array_update_79196[3] = add_78772 == 32'h0000_0003 ? array_update_79194 : array_update_79183[3];
  assign array_update_79196[4] = add_78772 == 32'h0000_0004 ? array_update_79194 : array_update_79183[4];
  assign array_update_79196[5] = add_78772 == 32'h0000_0005 ? array_update_79194 : array_update_79183[5];
  assign array_update_79196[6] = add_78772 == 32'h0000_0006 ? array_update_79194 : array_update_79183[6];
  assign array_update_79196[7] = add_78772 == 32'h0000_0007 ? array_update_79194 : array_update_79183[7];
  assign array_update_79196[8] = add_78772 == 32'h0000_0008 ? array_update_79194 : array_update_79183[8];
  assign array_update_79196[9] = add_78772 == 32'h0000_0009 ? array_update_79194 : array_update_79183[9];
  assign array_index_79198 = array_update_72021[add_79195 > 32'h0000_0009 ? 4'h9 : add_79195[3:0]];
  assign array_index_79199 = array_update_79196[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_79203 = smul32b_32b_x_32b(array_index_78779[add_79195 > 32'h0000_0009 ? 4'h9 : add_79195[3:0]], array_index_79198[add_79180 > 32'h0000_0009 ? 4'h9 : add_79180[3:0]]);
  assign add_79205 = array_index_79199[add_79180 > 32'h0000_0009 ? 4'h9 : add_79180[3:0]] + smul_79203;
  assign array_update_79207[0] = add_79180 == 32'h0000_0000 ? add_79205 : array_index_79199[0];
  assign array_update_79207[1] = add_79180 == 32'h0000_0001 ? add_79205 : array_index_79199[1];
  assign array_update_79207[2] = add_79180 == 32'h0000_0002 ? add_79205 : array_index_79199[2];
  assign array_update_79207[3] = add_79180 == 32'h0000_0003 ? add_79205 : array_index_79199[3];
  assign array_update_79207[4] = add_79180 == 32'h0000_0004 ? add_79205 : array_index_79199[4];
  assign array_update_79207[5] = add_79180 == 32'h0000_0005 ? add_79205 : array_index_79199[5];
  assign array_update_79207[6] = add_79180 == 32'h0000_0006 ? add_79205 : array_index_79199[6];
  assign array_update_79207[7] = add_79180 == 32'h0000_0007 ? add_79205 : array_index_79199[7];
  assign array_update_79207[8] = add_79180 == 32'h0000_0008 ? add_79205 : array_index_79199[8];
  assign array_update_79207[9] = add_79180 == 32'h0000_0009 ? add_79205 : array_index_79199[9];
  assign add_79208 = add_79195 + 32'h0000_0001;
  assign array_update_79209[0] = add_78772 == 32'h0000_0000 ? array_update_79207 : array_update_79196[0];
  assign array_update_79209[1] = add_78772 == 32'h0000_0001 ? array_update_79207 : array_update_79196[1];
  assign array_update_79209[2] = add_78772 == 32'h0000_0002 ? array_update_79207 : array_update_79196[2];
  assign array_update_79209[3] = add_78772 == 32'h0000_0003 ? array_update_79207 : array_update_79196[3];
  assign array_update_79209[4] = add_78772 == 32'h0000_0004 ? array_update_79207 : array_update_79196[4];
  assign array_update_79209[5] = add_78772 == 32'h0000_0005 ? array_update_79207 : array_update_79196[5];
  assign array_update_79209[6] = add_78772 == 32'h0000_0006 ? array_update_79207 : array_update_79196[6];
  assign array_update_79209[7] = add_78772 == 32'h0000_0007 ? array_update_79207 : array_update_79196[7];
  assign array_update_79209[8] = add_78772 == 32'h0000_0008 ? array_update_79207 : array_update_79196[8];
  assign array_update_79209[9] = add_78772 == 32'h0000_0009 ? array_update_79207 : array_update_79196[9];
  assign array_index_79211 = array_update_72021[add_79208 > 32'h0000_0009 ? 4'h9 : add_79208[3:0]];
  assign array_index_79212 = array_update_79209[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_79216 = smul32b_32b_x_32b(array_index_78779[add_79208 > 32'h0000_0009 ? 4'h9 : add_79208[3:0]], array_index_79211[add_79180 > 32'h0000_0009 ? 4'h9 : add_79180[3:0]]);
  assign add_79218 = array_index_79212[add_79180 > 32'h0000_0009 ? 4'h9 : add_79180[3:0]] + smul_79216;
  assign array_update_79220[0] = add_79180 == 32'h0000_0000 ? add_79218 : array_index_79212[0];
  assign array_update_79220[1] = add_79180 == 32'h0000_0001 ? add_79218 : array_index_79212[1];
  assign array_update_79220[2] = add_79180 == 32'h0000_0002 ? add_79218 : array_index_79212[2];
  assign array_update_79220[3] = add_79180 == 32'h0000_0003 ? add_79218 : array_index_79212[3];
  assign array_update_79220[4] = add_79180 == 32'h0000_0004 ? add_79218 : array_index_79212[4];
  assign array_update_79220[5] = add_79180 == 32'h0000_0005 ? add_79218 : array_index_79212[5];
  assign array_update_79220[6] = add_79180 == 32'h0000_0006 ? add_79218 : array_index_79212[6];
  assign array_update_79220[7] = add_79180 == 32'h0000_0007 ? add_79218 : array_index_79212[7];
  assign array_update_79220[8] = add_79180 == 32'h0000_0008 ? add_79218 : array_index_79212[8];
  assign array_update_79220[9] = add_79180 == 32'h0000_0009 ? add_79218 : array_index_79212[9];
  assign add_79221 = add_79208 + 32'h0000_0001;
  assign array_update_79222[0] = add_78772 == 32'h0000_0000 ? array_update_79220 : array_update_79209[0];
  assign array_update_79222[1] = add_78772 == 32'h0000_0001 ? array_update_79220 : array_update_79209[1];
  assign array_update_79222[2] = add_78772 == 32'h0000_0002 ? array_update_79220 : array_update_79209[2];
  assign array_update_79222[3] = add_78772 == 32'h0000_0003 ? array_update_79220 : array_update_79209[3];
  assign array_update_79222[4] = add_78772 == 32'h0000_0004 ? array_update_79220 : array_update_79209[4];
  assign array_update_79222[5] = add_78772 == 32'h0000_0005 ? array_update_79220 : array_update_79209[5];
  assign array_update_79222[6] = add_78772 == 32'h0000_0006 ? array_update_79220 : array_update_79209[6];
  assign array_update_79222[7] = add_78772 == 32'h0000_0007 ? array_update_79220 : array_update_79209[7];
  assign array_update_79222[8] = add_78772 == 32'h0000_0008 ? array_update_79220 : array_update_79209[8];
  assign array_update_79222[9] = add_78772 == 32'h0000_0009 ? array_update_79220 : array_update_79209[9];
  assign array_index_79224 = array_update_72021[add_79221 > 32'h0000_0009 ? 4'h9 : add_79221[3:0]];
  assign array_index_79225 = array_update_79222[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_79229 = smul32b_32b_x_32b(array_index_78779[add_79221 > 32'h0000_0009 ? 4'h9 : add_79221[3:0]], array_index_79224[add_79180 > 32'h0000_0009 ? 4'h9 : add_79180[3:0]]);
  assign add_79231 = array_index_79225[add_79180 > 32'h0000_0009 ? 4'h9 : add_79180[3:0]] + smul_79229;
  assign array_update_79233[0] = add_79180 == 32'h0000_0000 ? add_79231 : array_index_79225[0];
  assign array_update_79233[1] = add_79180 == 32'h0000_0001 ? add_79231 : array_index_79225[1];
  assign array_update_79233[2] = add_79180 == 32'h0000_0002 ? add_79231 : array_index_79225[2];
  assign array_update_79233[3] = add_79180 == 32'h0000_0003 ? add_79231 : array_index_79225[3];
  assign array_update_79233[4] = add_79180 == 32'h0000_0004 ? add_79231 : array_index_79225[4];
  assign array_update_79233[5] = add_79180 == 32'h0000_0005 ? add_79231 : array_index_79225[5];
  assign array_update_79233[6] = add_79180 == 32'h0000_0006 ? add_79231 : array_index_79225[6];
  assign array_update_79233[7] = add_79180 == 32'h0000_0007 ? add_79231 : array_index_79225[7];
  assign array_update_79233[8] = add_79180 == 32'h0000_0008 ? add_79231 : array_index_79225[8];
  assign array_update_79233[9] = add_79180 == 32'h0000_0009 ? add_79231 : array_index_79225[9];
  assign add_79234 = add_79221 + 32'h0000_0001;
  assign array_update_79235[0] = add_78772 == 32'h0000_0000 ? array_update_79233 : array_update_79222[0];
  assign array_update_79235[1] = add_78772 == 32'h0000_0001 ? array_update_79233 : array_update_79222[1];
  assign array_update_79235[2] = add_78772 == 32'h0000_0002 ? array_update_79233 : array_update_79222[2];
  assign array_update_79235[3] = add_78772 == 32'h0000_0003 ? array_update_79233 : array_update_79222[3];
  assign array_update_79235[4] = add_78772 == 32'h0000_0004 ? array_update_79233 : array_update_79222[4];
  assign array_update_79235[5] = add_78772 == 32'h0000_0005 ? array_update_79233 : array_update_79222[5];
  assign array_update_79235[6] = add_78772 == 32'h0000_0006 ? array_update_79233 : array_update_79222[6];
  assign array_update_79235[7] = add_78772 == 32'h0000_0007 ? array_update_79233 : array_update_79222[7];
  assign array_update_79235[8] = add_78772 == 32'h0000_0008 ? array_update_79233 : array_update_79222[8];
  assign array_update_79235[9] = add_78772 == 32'h0000_0009 ? array_update_79233 : array_update_79222[9];
  assign array_index_79237 = array_update_72021[add_79234 > 32'h0000_0009 ? 4'h9 : add_79234[3:0]];
  assign array_index_79238 = array_update_79235[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_79242 = smul32b_32b_x_32b(array_index_78779[add_79234 > 32'h0000_0009 ? 4'h9 : add_79234[3:0]], array_index_79237[add_79180 > 32'h0000_0009 ? 4'h9 : add_79180[3:0]]);
  assign add_79244 = array_index_79238[add_79180 > 32'h0000_0009 ? 4'h9 : add_79180[3:0]] + smul_79242;
  assign array_update_79246[0] = add_79180 == 32'h0000_0000 ? add_79244 : array_index_79238[0];
  assign array_update_79246[1] = add_79180 == 32'h0000_0001 ? add_79244 : array_index_79238[1];
  assign array_update_79246[2] = add_79180 == 32'h0000_0002 ? add_79244 : array_index_79238[2];
  assign array_update_79246[3] = add_79180 == 32'h0000_0003 ? add_79244 : array_index_79238[3];
  assign array_update_79246[4] = add_79180 == 32'h0000_0004 ? add_79244 : array_index_79238[4];
  assign array_update_79246[5] = add_79180 == 32'h0000_0005 ? add_79244 : array_index_79238[5];
  assign array_update_79246[6] = add_79180 == 32'h0000_0006 ? add_79244 : array_index_79238[6];
  assign array_update_79246[7] = add_79180 == 32'h0000_0007 ? add_79244 : array_index_79238[7];
  assign array_update_79246[8] = add_79180 == 32'h0000_0008 ? add_79244 : array_index_79238[8];
  assign array_update_79246[9] = add_79180 == 32'h0000_0009 ? add_79244 : array_index_79238[9];
  assign add_79247 = add_79234 + 32'h0000_0001;
  assign array_update_79248[0] = add_78772 == 32'h0000_0000 ? array_update_79246 : array_update_79235[0];
  assign array_update_79248[1] = add_78772 == 32'h0000_0001 ? array_update_79246 : array_update_79235[1];
  assign array_update_79248[2] = add_78772 == 32'h0000_0002 ? array_update_79246 : array_update_79235[2];
  assign array_update_79248[3] = add_78772 == 32'h0000_0003 ? array_update_79246 : array_update_79235[3];
  assign array_update_79248[4] = add_78772 == 32'h0000_0004 ? array_update_79246 : array_update_79235[4];
  assign array_update_79248[5] = add_78772 == 32'h0000_0005 ? array_update_79246 : array_update_79235[5];
  assign array_update_79248[6] = add_78772 == 32'h0000_0006 ? array_update_79246 : array_update_79235[6];
  assign array_update_79248[7] = add_78772 == 32'h0000_0007 ? array_update_79246 : array_update_79235[7];
  assign array_update_79248[8] = add_78772 == 32'h0000_0008 ? array_update_79246 : array_update_79235[8];
  assign array_update_79248[9] = add_78772 == 32'h0000_0009 ? array_update_79246 : array_update_79235[9];
  assign array_index_79250 = array_update_72021[add_79247 > 32'h0000_0009 ? 4'h9 : add_79247[3:0]];
  assign array_index_79251 = array_update_79248[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_79255 = smul32b_32b_x_32b(array_index_78779[add_79247 > 32'h0000_0009 ? 4'h9 : add_79247[3:0]], array_index_79250[add_79180 > 32'h0000_0009 ? 4'h9 : add_79180[3:0]]);
  assign add_79257 = array_index_79251[add_79180 > 32'h0000_0009 ? 4'h9 : add_79180[3:0]] + smul_79255;
  assign array_update_79259[0] = add_79180 == 32'h0000_0000 ? add_79257 : array_index_79251[0];
  assign array_update_79259[1] = add_79180 == 32'h0000_0001 ? add_79257 : array_index_79251[1];
  assign array_update_79259[2] = add_79180 == 32'h0000_0002 ? add_79257 : array_index_79251[2];
  assign array_update_79259[3] = add_79180 == 32'h0000_0003 ? add_79257 : array_index_79251[3];
  assign array_update_79259[4] = add_79180 == 32'h0000_0004 ? add_79257 : array_index_79251[4];
  assign array_update_79259[5] = add_79180 == 32'h0000_0005 ? add_79257 : array_index_79251[5];
  assign array_update_79259[6] = add_79180 == 32'h0000_0006 ? add_79257 : array_index_79251[6];
  assign array_update_79259[7] = add_79180 == 32'h0000_0007 ? add_79257 : array_index_79251[7];
  assign array_update_79259[8] = add_79180 == 32'h0000_0008 ? add_79257 : array_index_79251[8];
  assign array_update_79259[9] = add_79180 == 32'h0000_0009 ? add_79257 : array_index_79251[9];
  assign add_79260 = add_79247 + 32'h0000_0001;
  assign array_update_79261[0] = add_78772 == 32'h0000_0000 ? array_update_79259 : array_update_79248[0];
  assign array_update_79261[1] = add_78772 == 32'h0000_0001 ? array_update_79259 : array_update_79248[1];
  assign array_update_79261[2] = add_78772 == 32'h0000_0002 ? array_update_79259 : array_update_79248[2];
  assign array_update_79261[3] = add_78772 == 32'h0000_0003 ? array_update_79259 : array_update_79248[3];
  assign array_update_79261[4] = add_78772 == 32'h0000_0004 ? array_update_79259 : array_update_79248[4];
  assign array_update_79261[5] = add_78772 == 32'h0000_0005 ? array_update_79259 : array_update_79248[5];
  assign array_update_79261[6] = add_78772 == 32'h0000_0006 ? array_update_79259 : array_update_79248[6];
  assign array_update_79261[7] = add_78772 == 32'h0000_0007 ? array_update_79259 : array_update_79248[7];
  assign array_update_79261[8] = add_78772 == 32'h0000_0008 ? array_update_79259 : array_update_79248[8];
  assign array_update_79261[9] = add_78772 == 32'h0000_0009 ? array_update_79259 : array_update_79248[9];
  assign array_index_79263 = array_update_72021[add_79260 > 32'h0000_0009 ? 4'h9 : add_79260[3:0]];
  assign array_index_79264 = array_update_79261[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_79268 = smul32b_32b_x_32b(array_index_78779[add_79260 > 32'h0000_0009 ? 4'h9 : add_79260[3:0]], array_index_79263[add_79180 > 32'h0000_0009 ? 4'h9 : add_79180[3:0]]);
  assign add_79270 = array_index_79264[add_79180 > 32'h0000_0009 ? 4'h9 : add_79180[3:0]] + smul_79268;
  assign array_update_79272[0] = add_79180 == 32'h0000_0000 ? add_79270 : array_index_79264[0];
  assign array_update_79272[1] = add_79180 == 32'h0000_0001 ? add_79270 : array_index_79264[1];
  assign array_update_79272[2] = add_79180 == 32'h0000_0002 ? add_79270 : array_index_79264[2];
  assign array_update_79272[3] = add_79180 == 32'h0000_0003 ? add_79270 : array_index_79264[3];
  assign array_update_79272[4] = add_79180 == 32'h0000_0004 ? add_79270 : array_index_79264[4];
  assign array_update_79272[5] = add_79180 == 32'h0000_0005 ? add_79270 : array_index_79264[5];
  assign array_update_79272[6] = add_79180 == 32'h0000_0006 ? add_79270 : array_index_79264[6];
  assign array_update_79272[7] = add_79180 == 32'h0000_0007 ? add_79270 : array_index_79264[7];
  assign array_update_79272[8] = add_79180 == 32'h0000_0008 ? add_79270 : array_index_79264[8];
  assign array_update_79272[9] = add_79180 == 32'h0000_0009 ? add_79270 : array_index_79264[9];
  assign add_79273 = add_79260 + 32'h0000_0001;
  assign array_update_79274[0] = add_78772 == 32'h0000_0000 ? array_update_79272 : array_update_79261[0];
  assign array_update_79274[1] = add_78772 == 32'h0000_0001 ? array_update_79272 : array_update_79261[1];
  assign array_update_79274[2] = add_78772 == 32'h0000_0002 ? array_update_79272 : array_update_79261[2];
  assign array_update_79274[3] = add_78772 == 32'h0000_0003 ? array_update_79272 : array_update_79261[3];
  assign array_update_79274[4] = add_78772 == 32'h0000_0004 ? array_update_79272 : array_update_79261[4];
  assign array_update_79274[5] = add_78772 == 32'h0000_0005 ? array_update_79272 : array_update_79261[5];
  assign array_update_79274[6] = add_78772 == 32'h0000_0006 ? array_update_79272 : array_update_79261[6];
  assign array_update_79274[7] = add_78772 == 32'h0000_0007 ? array_update_79272 : array_update_79261[7];
  assign array_update_79274[8] = add_78772 == 32'h0000_0008 ? array_update_79272 : array_update_79261[8];
  assign array_update_79274[9] = add_78772 == 32'h0000_0009 ? array_update_79272 : array_update_79261[9];
  assign array_index_79276 = array_update_72021[add_79273 > 32'h0000_0009 ? 4'h9 : add_79273[3:0]];
  assign array_index_79277 = array_update_79274[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_79281 = smul32b_32b_x_32b(array_index_78779[add_79273 > 32'h0000_0009 ? 4'h9 : add_79273[3:0]], array_index_79276[add_79180 > 32'h0000_0009 ? 4'h9 : add_79180[3:0]]);
  assign add_79283 = array_index_79277[add_79180 > 32'h0000_0009 ? 4'h9 : add_79180[3:0]] + smul_79281;
  assign array_update_79285[0] = add_79180 == 32'h0000_0000 ? add_79283 : array_index_79277[0];
  assign array_update_79285[1] = add_79180 == 32'h0000_0001 ? add_79283 : array_index_79277[1];
  assign array_update_79285[2] = add_79180 == 32'h0000_0002 ? add_79283 : array_index_79277[2];
  assign array_update_79285[3] = add_79180 == 32'h0000_0003 ? add_79283 : array_index_79277[3];
  assign array_update_79285[4] = add_79180 == 32'h0000_0004 ? add_79283 : array_index_79277[4];
  assign array_update_79285[5] = add_79180 == 32'h0000_0005 ? add_79283 : array_index_79277[5];
  assign array_update_79285[6] = add_79180 == 32'h0000_0006 ? add_79283 : array_index_79277[6];
  assign array_update_79285[7] = add_79180 == 32'h0000_0007 ? add_79283 : array_index_79277[7];
  assign array_update_79285[8] = add_79180 == 32'h0000_0008 ? add_79283 : array_index_79277[8];
  assign array_update_79285[9] = add_79180 == 32'h0000_0009 ? add_79283 : array_index_79277[9];
  assign add_79286 = add_79273 + 32'h0000_0001;
  assign array_update_79287[0] = add_78772 == 32'h0000_0000 ? array_update_79285 : array_update_79274[0];
  assign array_update_79287[1] = add_78772 == 32'h0000_0001 ? array_update_79285 : array_update_79274[1];
  assign array_update_79287[2] = add_78772 == 32'h0000_0002 ? array_update_79285 : array_update_79274[2];
  assign array_update_79287[3] = add_78772 == 32'h0000_0003 ? array_update_79285 : array_update_79274[3];
  assign array_update_79287[4] = add_78772 == 32'h0000_0004 ? array_update_79285 : array_update_79274[4];
  assign array_update_79287[5] = add_78772 == 32'h0000_0005 ? array_update_79285 : array_update_79274[5];
  assign array_update_79287[6] = add_78772 == 32'h0000_0006 ? array_update_79285 : array_update_79274[6];
  assign array_update_79287[7] = add_78772 == 32'h0000_0007 ? array_update_79285 : array_update_79274[7];
  assign array_update_79287[8] = add_78772 == 32'h0000_0008 ? array_update_79285 : array_update_79274[8];
  assign array_update_79287[9] = add_78772 == 32'h0000_0009 ? array_update_79285 : array_update_79274[9];
  assign array_index_79289 = array_update_72021[add_79286 > 32'h0000_0009 ? 4'h9 : add_79286[3:0]];
  assign array_index_79290 = array_update_79287[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_79294 = smul32b_32b_x_32b(array_index_78779[add_79286 > 32'h0000_0009 ? 4'h9 : add_79286[3:0]], array_index_79289[add_79180 > 32'h0000_0009 ? 4'h9 : add_79180[3:0]]);
  assign add_79296 = array_index_79290[add_79180 > 32'h0000_0009 ? 4'h9 : add_79180[3:0]] + smul_79294;
  assign array_update_79298[0] = add_79180 == 32'h0000_0000 ? add_79296 : array_index_79290[0];
  assign array_update_79298[1] = add_79180 == 32'h0000_0001 ? add_79296 : array_index_79290[1];
  assign array_update_79298[2] = add_79180 == 32'h0000_0002 ? add_79296 : array_index_79290[2];
  assign array_update_79298[3] = add_79180 == 32'h0000_0003 ? add_79296 : array_index_79290[3];
  assign array_update_79298[4] = add_79180 == 32'h0000_0004 ? add_79296 : array_index_79290[4];
  assign array_update_79298[5] = add_79180 == 32'h0000_0005 ? add_79296 : array_index_79290[5];
  assign array_update_79298[6] = add_79180 == 32'h0000_0006 ? add_79296 : array_index_79290[6];
  assign array_update_79298[7] = add_79180 == 32'h0000_0007 ? add_79296 : array_index_79290[7];
  assign array_update_79298[8] = add_79180 == 32'h0000_0008 ? add_79296 : array_index_79290[8];
  assign array_update_79298[9] = add_79180 == 32'h0000_0009 ? add_79296 : array_index_79290[9];
  assign add_79299 = add_79286 + 32'h0000_0001;
  assign array_update_79300[0] = add_78772 == 32'h0000_0000 ? array_update_79298 : array_update_79287[0];
  assign array_update_79300[1] = add_78772 == 32'h0000_0001 ? array_update_79298 : array_update_79287[1];
  assign array_update_79300[2] = add_78772 == 32'h0000_0002 ? array_update_79298 : array_update_79287[2];
  assign array_update_79300[3] = add_78772 == 32'h0000_0003 ? array_update_79298 : array_update_79287[3];
  assign array_update_79300[4] = add_78772 == 32'h0000_0004 ? array_update_79298 : array_update_79287[4];
  assign array_update_79300[5] = add_78772 == 32'h0000_0005 ? array_update_79298 : array_update_79287[5];
  assign array_update_79300[6] = add_78772 == 32'h0000_0006 ? array_update_79298 : array_update_79287[6];
  assign array_update_79300[7] = add_78772 == 32'h0000_0007 ? array_update_79298 : array_update_79287[7];
  assign array_update_79300[8] = add_78772 == 32'h0000_0008 ? array_update_79298 : array_update_79287[8];
  assign array_update_79300[9] = add_78772 == 32'h0000_0009 ? array_update_79298 : array_update_79287[9];
  assign array_index_79302 = array_update_72021[add_79299 > 32'h0000_0009 ? 4'h9 : add_79299[3:0]];
  assign array_index_79303 = array_update_79300[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_79307 = smul32b_32b_x_32b(array_index_78779[add_79299 > 32'h0000_0009 ? 4'h9 : add_79299[3:0]], array_index_79302[add_79180 > 32'h0000_0009 ? 4'h9 : add_79180[3:0]]);
  assign add_79309 = array_index_79303[add_79180 > 32'h0000_0009 ? 4'h9 : add_79180[3:0]] + smul_79307;
  assign array_update_79310[0] = add_79180 == 32'h0000_0000 ? add_79309 : array_index_79303[0];
  assign array_update_79310[1] = add_79180 == 32'h0000_0001 ? add_79309 : array_index_79303[1];
  assign array_update_79310[2] = add_79180 == 32'h0000_0002 ? add_79309 : array_index_79303[2];
  assign array_update_79310[3] = add_79180 == 32'h0000_0003 ? add_79309 : array_index_79303[3];
  assign array_update_79310[4] = add_79180 == 32'h0000_0004 ? add_79309 : array_index_79303[4];
  assign array_update_79310[5] = add_79180 == 32'h0000_0005 ? add_79309 : array_index_79303[5];
  assign array_update_79310[6] = add_79180 == 32'h0000_0006 ? add_79309 : array_index_79303[6];
  assign array_update_79310[7] = add_79180 == 32'h0000_0007 ? add_79309 : array_index_79303[7];
  assign array_update_79310[8] = add_79180 == 32'h0000_0008 ? add_79309 : array_index_79303[8];
  assign array_update_79310[9] = add_79180 == 32'h0000_0009 ? add_79309 : array_index_79303[9];
  assign array_update_79311[0] = add_78772 == 32'h0000_0000 ? array_update_79310 : array_update_79300[0];
  assign array_update_79311[1] = add_78772 == 32'h0000_0001 ? array_update_79310 : array_update_79300[1];
  assign array_update_79311[2] = add_78772 == 32'h0000_0002 ? array_update_79310 : array_update_79300[2];
  assign array_update_79311[3] = add_78772 == 32'h0000_0003 ? array_update_79310 : array_update_79300[3];
  assign array_update_79311[4] = add_78772 == 32'h0000_0004 ? array_update_79310 : array_update_79300[4];
  assign array_update_79311[5] = add_78772 == 32'h0000_0005 ? array_update_79310 : array_update_79300[5];
  assign array_update_79311[6] = add_78772 == 32'h0000_0006 ? array_update_79310 : array_update_79300[6];
  assign array_update_79311[7] = add_78772 == 32'h0000_0007 ? array_update_79310 : array_update_79300[7];
  assign array_update_79311[8] = add_78772 == 32'h0000_0008 ? array_update_79310 : array_update_79300[8];
  assign array_update_79311[9] = add_78772 == 32'h0000_0009 ? array_update_79310 : array_update_79300[9];
  assign array_index_79313 = array_update_79311[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign add_79315 = add_79180 + 32'h0000_0001;
  assign array_update_79316[0] = add_79315 == 32'h0000_0000 ? 32'h0000_0000 : array_index_79313[0];
  assign array_update_79316[1] = add_79315 == 32'h0000_0001 ? 32'h0000_0000 : array_index_79313[1];
  assign array_update_79316[2] = add_79315 == 32'h0000_0002 ? 32'h0000_0000 : array_index_79313[2];
  assign array_update_79316[3] = add_79315 == 32'h0000_0003 ? 32'h0000_0000 : array_index_79313[3];
  assign array_update_79316[4] = add_79315 == 32'h0000_0004 ? 32'h0000_0000 : array_index_79313[4];
  assign array_update_79316[5] = add_79315 == 32'h0000_0005 ? 32'h0000_0000 : array_index_79313[5];
  assign array_update_79316[6] = add_79315 == 32'h0000_0006 ? 32'h0000_0000 : array_index_79313[6];
  assign array_update_79316[7] = add_79315 == 32'h0000_0007 ? 32'h0000_0000 : array_index_79313[7];
  assign array_update_79316[8] = add_79315 == 32'h0000_0008 ? 32'h0000_0000 : array_index_79313[8];
  assign array_update_79316[9] = add_79315 == 32'h0000_0009 ? 32'h0000_0000 : array_index_79313[9];
  assign literal_79317 = 32'h0000_0000;
  assign array_update_79318[0] = add_78772 == 32'h0000_0000 ? array_update_79316 : array_update_79311[0];
  assign array_update_79318[1] = add_78772 == 32'h0000_0001 ? array_update_79316 : array_update_79311[1];
  assign array_update_79318[2] = add_78772 == 32'h0000_0002 ? array_update_79316 : array_update_79311[2];
  assign array_update_79318[3] = add_78772 == 32'h0000_0003 ? array_update_79316 : array_update_79311[3];
  assign array_update_79318[4] = add_78772 == 32'h0000_0004 ? array_update_79316 : array_update_79311[4];
  assign array_update_79318[5] = add_78772 == 32'h0000_0005 ? array_update_79316 : array_update_79311[5];
  assign array_update_79318[6] = add_78772 == 32'h0000_0006 ? array_update_79316 : array_update_79311[6];
  assign array_update_79318[7] = add_78772 == 32'h0000_0007 ? array_update_79316 : array_update_79311[7];
  assign array_update_79318[8] = add_78772 == 32'h0000_0008 ? array_update_79316 : array_update_79311[8];
  assign array_update_79318[9] = add_78772 == 32'h0000_0009 ? array_update_79316 : array_update_79311[9];
  assign array_index_79320 = array_update_72021[literal_79317 > 32'h0000_0009 ? 4'h9 : literal_79317[3:0]];
  assign array_index_79321 = array_update_79318[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_79325 = smul32b_32b_x_32b(array_index_78779[literal_79317 > 32'h0000_0009 ? 4'h9 : literal_79317[3:0]], array_index_79320[add_79315 > 32'h0000_0009 ? 4'h9 : add_79315[3:0]]);
  assign add_79327 = array_index_79321[add_79315 > 32'h0000_0009 ? 4'h9 : add_79315[3:0]] + smul_79325;
  assign array_update_79329[0] = add_79315 == 32'h0000_0000 ? add_79327 : array_index_79321[0];
  assign array_update_79329[1] = add_79315 == 32'h0000_0001 ? add_79327 : array_index_79321[1];
  assign array_update_79329[2] = add_79315 == 32'h0000_0002 ? add_79327 : array_index_79321[2];
  assign array_update_79329[3] = add_79315 == 32'h0000_0003 ? add_79327 : array_index_79321[3];
  assign array_update_79329[4] = add_79315 == 32'h0000_0004 ? add_79327 : array_index_79321[4];
  assign array_update_79329[5] = add_79315 == 32'h0000_0005 ? add_79327 : array_index_79321[5];
  assign array_update_79329[6] = add_79315 == 32'h0000_0006 ? add_79327 : array_index_79321[6];
  assign array_update_79329[7] = add_79315 == 32'h0000_0007 ? add_79327 : array_index_79321[7];
  assign array_update_79329[8] = add_79315 == 32'h0000_0008 ? add_79327 : array_index_79321[8];
  assign array_update_79329[9] = add_79315 == 32'h0000_0009 ? add_79327 : array_index_79321[9];
  assign add_79330 = literal_79317 + 32'h0000_0001;
  assign array_update_79331[0] = add_78772 == 32'h0000_0000 ? array_update_79329 : array_update_79318[0];
  assign array_update_79331[1] = add_78772 == 32'h0000_0001 ? array_update_79329 : array_update_79318[1];
  assign array_update_79331[2] = add_78772 == 32'h0000_0002 ? array_update_79329 : array_update_79318[2];
  assign array_update_79331[3] = add_78772 == 32'h0000_0003 ? array_update_79329 : array_update_79318[3];
  assign array_update_79331[4] = add_78772 == 32'h0000_0004 ? array_update_79329 : array_update_79318[4];
  assign array_update_79331[5] = add_78772 == 32'h0000_0005 ? array_update_79329 : array_update_79318[5];
  assign array_update_79331[6] = add_78772 == 32'h0000_0006 ? array_update_79329 : array_update_79318[6];
  assign array_update_79331[7] = add_78772 == 32'h0000_0007 ? array_update_79329 : array_update_79318[7];
  assign array_update_79331[8] = add_78772 == 32'h0000_0008 ? array_update_79329 : array_update_79318[8];
  assign array_update_79331[9] = add_78772 == 32'h0000_0009 ? array_update_79329 : array_update_79318[9];
  assign array_index_79333 = array_update_72021[add_79330 > 32'h0000_0009 ? 4'h9 : add_79330[3:0]];
  assign array_index_79334 = array_update_79331[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_79338 = smul32b_32b_x_32b(array_index_78779[add_79330 > 32'h0000_0009 ? 4'h9 : add_79330[3:0]], array_index_79333[add_79315 > 32'h0000_0009 ? 4'h9 : add_79315[3:0]]);
  assign add_79340 = array_index_79334[add_79315 > 32'h0000_0009 ? 4'h9 : add_79315[3:0]] + smul_79338;
  assign array_update_79342[0] = add_79315 == 32'h0000_0000 ? add_79340 : array_index_79334[0];
  assign array_update_79342[1] = add_79315 == 32'h0000_0001 ? add_79340 : array_index_79334[1];
  assign array_update_79342[2] = add_79315 == 32'h0000_0002 ? add_79340 : array_index_79334[2];
  assign array_update_79342[3] = add_79315 == 32'h0000_0003 ? add_79340 : array_index_79334[3];
  assign array_update_79342[4] = add_79315 == 32'h0000_0004 ? add_79340 : array_index_79334[4];
  assign array_update_79342[5] = add_79315 == 32'h0000_0005 ? add_79340 : array_index_79334[5];
  assign array_update_79342[6] = add_79315 == 32'h0000_0006 ? add_79340 : array_index_79334[6];
  assign array_update_79342[7] = add_79315 == 32'h0000_0007 ? add_79340 : array_index_79334[7];
  assign array_update_79342[8] = add_79315 == 32'h0000_0008 ? add_79340 : array_index_79334[8];
  assign array_update_79342[9] = add_79315 == 32'h0000_0009 ? add_79340 : array_index_79334[9];
  assign add_79343 = add_79330 + 32'h0000_0001;
  assign array_update_79344[0] = add_78772 == 32'h0000_0000 ? array_update_79342 : array_update_79331[0];
  assign array_update_79344[1] = add_78772 == 32'h0000_0001 ? array_update_79342 : array_update_79331[1];
  assign array_update_79344[2] = add_78772 == 32'h0000_0002 ? array_update_79342 : array_update_79331[2];
  assign array_update_79344[3] = add_78772 == 32'h0000_0003 ? array_update_79342 : array_update_79331[3];
  assign array_update_79344[4] = add_78772 == 32'h0000_0004 ? array_update_79342 : array_update_79331[4];
  assign array_update_79344[5] = add_78772 == 32'h0000_0005 ? array_update_79342 : array_update_79331[5];
  assign array_update_79344[6] = add_78772 == 32'h0000_0006 ? array_update_79342 : array_update_79331[6];
  assign array_update_79344[7] = add_78772 == 32'h0000_0007 ? array_update_79342 : array_update_79331[7];
  assign array_update_79344[8] = add_78772 == 32'h0000_0008 ? array_update_79342 : array_update_79331[8];
  assign array_update_79344[9] = add_78772 == 32'h0000_0009 ? array_update_79342 : array_update_79331[9];
  assign array_index_79346 = array_update_72021[add_79343 > 32'h0000_0009 ? 4'h9 : add_79343[3:0]];
  assign array_index_79347 = array_update_79344[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_79351 = smul32b_32b_x_32b(array_index_78779[add_79343 > 32'h0000_0009 ? 4'h9 : add_79343[3:0]], array_index_79346[add_79315 > 32'h0000_0009 ? 4'h9 : add_79315[3:0]]);
  assign add_79353 = array_index_79347[add_79315 > 32'h0000_0009 ? 4'h9 : add_79315[3:0]] + smul_79351;
  assign array_update_79355[0] = add_79315 == 32'h0000_0000 ? add_79353 : array_index_79347[0];
  assign array_update_79355[1] = add_79315 == 32'h0000_0001 ? add_79353 : array_index_79347[1];
  assign array_update_79355[2] = add_79315 == 32'h0000_0002 ? add_79353 : array_index_79347[2];
  assign array_update_79355[3] = add_79315 == 32'h0000_0003 ? add_79353 : array_index_79347[3];
  assign array_update_79355[4] = add_79315 == 32'h0000_0004 ? add_79353 : array_index_79347[4];
  assign array_update_79355[5] = add_79315 == 32'h0000_0005 ? add_79353 : array_index_79347[5];
  assign array_update_79355[6] = add_79315 == 32'h0000_0006 ? add_79353 : array_index_79347[6];
  assign array_update_79355[7] = add_79315 == 32'h0000_0007 ? add_79353 : array_index_79347[7];
  assign array_update_79355[8] = add_79315 == 32'h0000_0008 ? add_79353 : array_index_79347[8];
  assign array_update_79355[9] = add_79315 == 32'h0000_0009 ? add_79353 : array_index_79347[9];
  assign add_79356 = add_79343 + 32'h0000_0001;
  assign array_update_79357[0] = add_78772 == 32'h0000_0000 ? array_update_79355 : array_update_79344[0];
  assign array_update_79357[1] = add_78772 == 32'h0000_0001 ? array_update_79355 : array_update_79344[1];
  assign array_update_79357[2] = add_78772 == 32'h0000_0002 ? array_update_79355 : array_update_79344[2];
  assign array_update_79357[3] = add_78772 == 32'h0000_0003 ? array_update_79355 : array_update_79344[3];
  assign array_update_79357[4] = add_78772 == 32'h0000_0004 ? array_update_79355 : array_update_79344[4];
  assign array_update_79357[5] = add_78772 == 32'h0000_0005 ? array_update_79355 : array_update_79344[5];
  assign array_update_79357[6] = add_78772 == 32'h0000_0006 ? array_update_79355 : array_update_79344[6];
  assign array_update_79357[7] = add_78772 == 32'h0000_0007 ? array_update_79355 : array_update_79344[7];
  assign array_update_79357[8] = add_78772 == 32'h0000_0008 ? array_update_79355 : array_update_79344[8];
  assign array_update_79357[9] = add_78772 == 32'h0000_0009 ? array_update_79355 : array_update_79344[9];
  assign array_index_79359 = array_update_72021[add_79356 > 32'h0000_0009 ? 4'h9 : add_79356[3:0]];
  assign array_index_79360 = array_update_79357[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_79364 = smul32b_32b_x_32b(array_index_78779[add_79356 > 32'h0000_0009 ? 4'h9 : add_79356[3:0]], array_index_79359[add_79315 > 32'h0000_0009 ? 4'h9 : add_79315[3:0]]);
  assign add_79366 = array_index_79360[add_79315 > 32'h0000_0009 ? 4'h9 : add_79315[3:0]] + smul_79364;
  assign array_update_79368[0] = add_79315 == 32'h0000_0000 ? add_79366 : array_index_79360[0];
  assign array_update_79368[1] = add_79315 == 32'h0000_0001 ? add_79366 : array_index_79360[1];
  assign array_update_79368[2] = add_79315 == 32'h0000_0002 ? add_79366 : array_index_79360[2];
  assign array_update_79368[3] = add_79315 == 32'h0000_0003 ? add_79366 : array_index_79360[3];
  assign array_update_79368[4] = add_79315 == 32'h0000_0004 ? add_79366 : array_index_79360[4];
  assign array_update_79368[5] = add_79315 == 32'h0000_0005 ? add_79366 : array_index_79360[5];
  assign array_update_79368[6] = add_79315 == 32'h0000_0006 ? add_79366 : array_index_79360[6];
  assign array_update_79368[7] = add_79315 == 32'h0000_0007 ? add_79366 : array_index_79360[7];
  assign array_update_79368[8] = add_79315 == 32'h0000_0008 ? add_79366 : array_index_79360[8];
  assign array_update_79368[9] = add_79315 == 32'h0000_0009 ? add_79366 : array_index_79360[9];
  assign add_79369 = add_79356 + 32'h0000_0001;
  assign array_update_79370[0] = add_78772 == 32'h0000_0000 ? array_update_79368 : array_update_79357[0];
  assign array_update_79370[1] = add_78772 == 32'h0000_0001 ? array_update_79368 : array_update_79357[1];
  assign array_update_79370[2] = add_78772 == 32'h0000_0002 ? array_update_79368 : array_update_79357[2];
  assign array_update_79370[3] = add_78772 == 32'h0000_0003 ? array_update_79368 : array_update_79357[3];
  assign array_update_79370[4] = add_78772 == 32'h0000_0004 ? array_update_79368 : array_update_79357[4];
  assign array_update_79370[5] = add_78772 == 32'h0000_0005 ? array_update_79368 : array_update_79357[5];
  assign array_update_79370[6] = add_78772 == 32'h0000_0006 ? array_update_79368 : array_update_79357[6];
  assign array_update_79370[7] = add_78772 == 32'h0000_0007 ? array_update_79368 : array_update_79357[7];
  assign array_update_79370[8] = add_78772 == 32'h0000_0008 ? array_update_79368 : array_update_79357[8];
  assign array_update_79370[9] = add_78772 == 32'h0000_0009 ? array_update_79368 : array_update_79357[9];
  assign array_index_79372 = array_update_72021[add_79369 > 32'h0000_0009 ? 4'h9 : add_79369[3:0]];
  assign array_index_79373 = array_update_79370[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_79377 = smul32b_32b_x_32b(array_index_78779[add_79369 > 32'h0000_0009 ? 4'h9 : add_79369[3:0]], array_index_79372[add_79315 > 32'h0000_0009 ? 4'h9 : add_79315[3:0]]);
  assign add_79379 = array_index_79373[add_79315 > 32'h0000_0009 ? 4'h9 : add_79315[3:0]] + smul_79377;
  assign array_update_79381[0] = add_79315 == 32'h0000_0000 ? add_79379 : array_index_79373[0];
  assign array_update_79381[1] = add_79315 == 32'h0000_0001 ? add_79379 : array_index_79373[1];
  assign array_update_79381[2] = add_79315 == 32'h0000_0002 ? add_79379 : array_index_79373[2];
  assign array_update_79381[3] = add_79315 == 32'h0000_0003 ? add_79379 : array_index_79373[3];
  assign array_update_79381[4] = add_79315 == 32'h0000_0004 ? add_79379 : array_index_79373[4];
  assign array_update_79381[5] = add_79315 == 32'h0000_0005 ? add_79379 : array_index_79373[5];
  assign array_update_79381[6] = add_79315 == 32'h0000_0006 ? add_79379 : array_index_79373[6];
  assign array_update_79381[7] = add_79315 == 32'h0000_0007 ? add_79379 : array_index_79373[7];
  assign array_update_79381[8] = add_79315 == 32'h0000_0008 ? add_79379 : array_index_79373[8];
  assign array_update_79381[9] = add_79315 == 32'h0000_0009 ? add_79379 : array_index_79373[9];
  assign add_79382 = add_79369 + 32'h0000_0001;
  assign array_update_79383[0] = add_78772 == 32'h0000_0000 ? array_update_79381 : array_update_79370[0];
  assign array_update_79383[1] = add_78772 == 32'h0000_0001 ? array_update_79381 : array_update_79370[1];
  assign array_update_79383[2] = add_78772 == 32'h0000_0002 ? array_update_79381 : array_update_79370[2];
  assign array_update_79383[3] = add_78772 == 32'h0000_0003 ? array_update_79381 : array_update_79370[3];
  assign array_update_79383[4] = add_78772 == 32'h0000_0004 ? array_update_79381 : array_update_79370[4];
  assign array_update_79383[5] = add_78772 == 32'h0000_0005 ? array_update_79381 : array_update_79370[5];
  assign array_update_79383[6] = add_78772 == 32'h0000_0006 ? array_update_79381 : array_update_79370[6];
  assign array_update_79383[7] = add_78772 == 32'h0000_0007 ? array_update_79381 : array_update_79370[7];
  assign array_update_79383[8] = add_78772 == 32'h0000_0008 ? array_update_79381 : array_update_79370[8];
  assign array_update_79383[9] = add_78772 == 32'h0000_0009 ? array_update_79381 : array_update_79370[9];
  assign array_index_79385 = array_update_72021[add_79382 > 32'h0000_0009 ? 4'h9 : add_79382[3:0]];
  assign array_index_79386 = array_update_79383[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_79390 = smul32b_32b_x_32b(array_index_78779[add_79382 > 32'h0000_0009 ? 4'h9 : add_79382[3:0]], array_index_79385[add_79315 > 32'h0000_0009 ? 4'h9 : add_79315[3:0]]);
  assign add_79392 = array_index_79386[add_79315 > 32'h0000_0009 ? 4'h9 : add_79315[3:0]] + smul_79390;
  assign array_update_79394[0] = add_79315 == 32'h0000_0000 ? add_79392 : array_index_79386[0];
  assign array_update_79394[1] = add_79315 == 32'h0000_0001 ? add_79392 : array_index_79386[1];
  assign array_update_79394[2] = add_79315 == 32'h0000_0002 ? add_79392 : array_index_79386[2];
  assign array_update_79394[3] = add_79315 == 32'h0000_0003 ? add_79392 : array_index_79386[3];
  assign array_update_79394[4] = add_79315 == 32'h0000_0004 ? add_79392 : array_index_79386[4];
  assign array_update_79394[5] = add_79315 == 32'h0000_0005 ? add_79392 : array_index_79386[5];
  assign array_update_79394[6] = add_79315 == 32'h0000_0006 ? add_79392 : array_index_79386[6];
  assign array_update_79394[7] = add_79315 == 32'h0000_0007 ? add_79392 : array_index_79386[7];
  assign array_update_79394[8] = add_79315 == 32'h0000_0008 ? add_79392 : array_index_79386[8];
  assign array_update_79394[9] = add_79315 == 32'h0000_0009 ? add_79392 : array_index_79386[9];
  assign add_79395 = add_79382 + 32'h0000_0001;
  assign array_update_79396[0] = add_78772 == 32'h0000_0000 ? array_update_79394 : array_update_79383[0];
  assign array_update_79396[1] = add_78772 == 32'h0000_0001 ? array_update_79394 : array_update_79383[1];
  assign array_update_79396[2] = add_78772 == 32'h0000_0002 ? array_update_79394 : array_update_79383[2];
  assign array_update_79396[3] = add_78772 == 32'h0000_0003 ? array_update_79394 : array_update_79383[3];
  assign array_update_79396[4] = add_78772 == 32'h0000_0004 ? array_update_79394 : array_update_79383[4];
  assign array_update_79396[5] = add_78772 == 32'h0000_0005 ? array_update_79394 : array_update_79383[5];
  assign array_update_79396[6] = add_78772 == 32'h0000_0006 ? array_update_79394 : array_update_79383[6];
  assign array_update_79396[7] = add_78772 == 32'h0000_0007 ? array_update_79394 : array_update_79383[7];
  assign array_update_79396[8] = add_78772 == 32'h0000_0008 ? array_update_79394 : array_update_79383[8];
  assign array_update_79396[9] = add_78772 == 32'h0000_0009 ? array_update_79394 : array_update_79383[9];
  assign array_index_79398 = array_update_72021[add_79395 > 32'h0000_0009 ? 4'h9 : add_79395[3:0]];
  assign array_index_79399 = array_update_79396[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_79403 = smul32b_32b_x_32b(array_index_78779[add_79395 > 32'h0000_0009 ? 4'h9 : add_79395[3:0]], array_index_79398[add_79315 > 32'h0000_0009 ? 4'h9 : add_79315[3:0]]);
  assign add_79405 = array_index_79399[add_79315 > 32'h0000_0009 ? 4'h9 : add_79315[3:0]] + smul_79403;
  assign array_update_79407[0] = add_79315 == 32'h0000_0000 ? add_79405 : array_index_79399[0];
  assign array_update_79407[1] = add_79315 == 32'h0000_0001 ? add_79405 : array_index_79399[1];
  assign array_update_79407[2] = add_79315 == 32'h0000_0002 ? add_79405 : array_index_79399[2];
  assign array_update_79407[3] = add_79315 == 32'h0000_0003 ? add_79405 : array_index_79399[3];
  assign array_update_79407[4] = add_79315 == 32'h0000_0004 ? add_79405 : array_index_79399[4];
  assign array_update_79407[5] = add_79315 == 32'h0000_0005 ? add_79405 : array_index_79399[5];
  assign array_update_79407[6] = add_79315 == 32'h0000_0006 ? add_79405 : array_index_79399[6];
  assign array_update_79407[7] = add_79315 == 32'h0000_0007 ? add_79405 : array_index_79399[7];
  assign array_update_79407[8] = add_79315 == 32'h0000_0008 ? add_79405 : array_index_79399[8];
  assign array_update_79407[9] = add_79315 == 32'h0000_0009 ? add_79405 : array_index_79399[9];
  assign add_79408 = add_79395 + 32'h0000_0001;
  assign array_update_79409[0] = add_78772 == 32'h0000_0000 ? array_update_79407 : array_update_79396[0];
  assign array_update_79409[1] = add_78772 == 32'h0000_0001 ? array_update_79407 : array_update_79396[1];
  assign array_update_79409[2] = add_78772 == 32'h0000_0002 ? array_update_79407 : array_update_79396[2];
  assign array_update_79409[3] = add_78772 == 32'h0000_0003 ? array_update_79407 : array_update_79396[3];
  assign array_update_79409[4] = add_78772 == 32'h0000_0004 ? array_update_79407 : array_update_79396[4];
  assign array_update_79409[5] = add_78772 == 32'h0000_0005 ? array_update_79407 : array_update_79396[5];
  assign array_update_79409[6] = add_78772 == 32'h0000_0006 ? array_update_79407 : array_update_79396[6];
  assign array_update_79409[7] = add_78772 == 32'h0000_0007 ? array_update_79407 : array_update_79396[7];
  assign array_update_79409[8] = add_78772 == 32'h0000_0008 ? array_update_79407 : array_update_79396[8];
  assign array_update_79409[9] = add_78772 == 32'h0000_0009 ? array_update_79407 : array_update_79396[9];
  assign array_index_79411 = array_update_72021[add_79408 > 32'h0000_0009 ? 4'h9 : add_79408[3:0]];
  assign array_index_79412 = array_update_79409[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_79416 = smul32b_32b_x_32b(array_index_78779[add_79408 > 32'h0000_0009 ? 4'h9 : add_79408[3:0]], array_index_79411[add_79315 > 32'h0000_0009 ? 4'h9 : add_79315[3:0]]);
  assign add_79418 = array_index_79412[add_79315 > 32'h0000_0009 ? 4'h9 : add_79315[3:0]] + smul_79416;
  assign array_update_79420[0] = add_79315 == 32'h0000_0000 ? add_79418 : array_index_79412[0];
  assign array_update_79420[1] = add_79315 == 32'h0000_0001 ? add_79418 : array_index_79412[1];
  assign array_update_79420[2] = add_79315 == 32'h0000_0002 ? add_79418 : array_index_79412[2];
  assign array_update_79420[3] = add_79315 == 32'h0000_0003 ? add_79418 : array_index_79412[3];
  assign array_update_79420[4] = add_79315 == 32'h0000_0004 ? add_79418 : array_index_79412[4];
  assign array_update_79420[5] = add_79315 == 32'h0000_0005 ? add_79418 : array_index_79412[5];
  assign array_update_79420[6] = add_79315 == 32'h0000_0006 ? add_79418 : array_index_79412[6];
  assign array_update_79420[7] = add_79315 == 32'h0000_0007 ? add_79418 : array_index_79412[7];
  assign array_update_79420[8] = add_79315 == 32'h0000_0008 ? add_79418 : array_index_79412[8];
  assign array_update_79420[9] = add_79315 == 32'h0000_0009 ? add_79418 : array_index_79412[9];
  assign add_79421 = add_79408 + 32'h0000_0001;
  assign array_update_79422[0] = add_78772 == 32'h0000_0000 ? array_update_79420 : array_update_79409[0];
  assign array_update_79422[1] = add_78772 == 32'h0000_0001 ? array_update_79420 : array_update_79409[1];
  assign array_update_79422[2] = add_78772 == 32'h0000_0002 ? array_update_79420 : array_update_79409[2];
  assign array_update_79422[3] = add_78772 == 32'h0000_0003 ? array_update_79420 : array_update_79409[3];
  assign array_update_79422[4] = add_78772 == 32'h0000_0004 ? array_update_79420 : array_update_79409[4];
  assign array_update_79422[5] = add_78772 == 32'h0000_0005 ? array_update_79420 : array_update_79409[5];
  assign array_update_79422[6] = add_78772 == 32'h0000_0006 ? array_update_79420 : array_update_79409[6];
  assign array_update_79422[7] = add_78772 == 32'h0000_0007 ? array_update_79420 : array_update_79409[7];
  assign array_update_79422[8] = add_78772 == 32'h0000_0008 ? array_update_79420 : array_update_79409[8];
  assign array_update_79422[9] = add_78772 == 32'h0000_0009 ? array_update_79420 : array_update_79409[9];
  assign array_index_79424 = array_update_72021[add_79421 > 32'h0000_0009 ? 4'h9 : add_79421[3:0]];
  assign array_index_79425 = array_update_79422[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_79429 = smul32b_32b_x_32b(array_index_78779[add_79421 > 32'h0000_0009 ? 4'h9 : add_79421[3:0]], array_index_79424[add_79315 > 32'h0000_0009 ? 4'h9 : add_79315[3:0]]);
  assign add_79431 = array_index_79425[add_79315 > 32'h0000_0009 ? 4'h9 : add_79315[3:0]] + smul_79429;
  assign array_update_79433[0] = add_79315 == 32'h0000_0000 ? add_79431 : array_index_79425[0];
  assign array_update_79433[1] = add_79315 == 32'h0000_0001 ? add_79431 : array_index_79425[1];
  assign array_update_79433[2] = add_79315 == 32'h0000_0002 ? add_79431 : array_index_79425[2];
  assign array_update_79433[3] = add_79315 == 32'h0000_0003 ? add_79431 : array_index_79425[3];
  assign array_update_79433[4] = add_79315 == 32'h0000_0004 ? add_79431 : array_index_79425[4];
  assign array_update_79433[5] = add_79315 == 32'h0000_0005 ? add_79431 : array_index_79425[5];
  assign array_update_79433[6] = add_79315 == 32'h0000_0006 ? add_79431 : array_index_79425[6];
  assign array_update_79433[7] = add_79315 == 32'h0000_0007 ? add_79431 : array_index_79425[7];
  assign array_update_79433[8] = add_79315 == 32'h0000_0008 ? add_79431 : array_index_79425[8];
  assign array_update_79433[9] = add_79315 == 32'h0000_0009 ? add_79431 : array_index_79425[9];
  assign add_79434 = add_79421 + 32'h0000_0001;
  assign array_update_79435[0] = add_78772 == 32'h0000_0000 ? array_update_79433 : array_update_79422[0];
  assign array_update_79435[1] = add_78772 == 32'h0000_0001 ? array_update_79433 : array_update_79422[1];
  assign array_update_79435[2] = add_78772 == 32'h0000_0002 ? array_update_79433 : array_update_79422[2];
  assign array_update_79435[3] = add_78772 == 32'h0000_0003 ? array_update_79433 : array_update_79422[3];
  assign array_update_79435[4] = add_78772 == 32'h0000_0004 ? array_update_79433 : array_update_79422[4];
  assign array_update_79435[5] = add_78772 == 32'h0000_0005 ? array_update_79433 : array_update_79422[5];
  assign array_update_79435[6] = add_78772 == 32'h0000_0006 ? array_update_79433 : array_update_79422[6];
  assign array_update_79435[7] = add_78772 == 32'h0000_0007 ? array_update_79433 : array_update_79422[7];
  assign array_update_79435[8] = add_78772 == 32'h0000_0008 ? array_update_79433 : array_update_79422[8];
  assign array_update_79435[9] = add_78772 == 32'h0000_0009 ? array_update_79433 : array_update_79422[9];
  assign array_index_79437 = array_update_72021[add_79434 > 32'h0000_0009 ? 4'h9 : add_79434[3:0]];
  assign array_index_79438 = array_update_79435[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_79442 = smul32b_32b_x_32b(array_index_78779[add_79434 > 32'h0000_0009 ? 4'h9 : add_79434[3:0]], array_index_79437[add_79315 > 32'h0000_0009 ? 4'h9 : add_79315[3:0]]);
  assign add_79444 = array_index_79438[add_79315 > 32'h0000_0009 ? 4'h9 : add_79315[3:0]] + smul_79442;
  assign array_update_79445[0] = add_79315 == 32'h0000_0000 ? add_79444 : array_index_79438[0];
  assign array_update_79445[1] = add_79315 == 32'h0000_0001 ? add_79444 : array_index_79438[1];
  assign array_update_79445[2] = add_79315 == 32'h0000_0002 ? add_79444 : array_index_79438[2];
  assign array_update_79445[3] = add_79315 == 32'h0000_0003 ? add_79444 : array_index_79438[3];
  assign array_update_79445[4] = add_79315 == 32'h0000_0004 ? add_79444 : array_index_79438[4];
  assign array_update_79445[5] = add_79315 == 32'h0000_0005 ? add_79444 : array_index_79438[5];
  assign array_update_79445[6] = add_79315 == 32'h0000_0006 ? add_79444 : array_index_79438[6];
  assign array_update_79445[7] = add_79315 == 32'h0000_0007 ? add_79444 : array_index_79438[7];
  assign array_update_79445[8] = add_79315 == 32'h0000_0008 ? add_79444 : array_index_79438[8];
  assign array_update_79445[9] = add_79315 == 32'h0000_0009 ? add_79444 : array_index_79438[9];
  assign array_update_79446[0] = add_78772 == 32'h0000_0000 ? array_update_79445 : array_update_79435[0];
  assign array_update_79446[1] = add_78772 == 32'h0000_0001 ? array_update_79445 : array_update_79435[1];
  assign array_update_79446[2] = add_78772 == 32'h0000_0002 ? array_update_79445 : array_update_79435[2];
  assign array_update_79446[3] = add_78772 == 32'h0000_0003 ? array_update_79445 : array_update_79435[3];
  assign array_update_79446[4] = add_78772 == 32'h0000_0004 ? array_update_79445 : array_update_79435[4];
  assign array_update_79446[5] = add_78772 == 32'h0000_0005 ? array_update_79445 : array_update_79435[5];
  assign array_update_79446[6] = add_78772 == 32'h0000_0006 ? array_update_79445 : array_update_79435[6];
  assign array_update_79446[7] = add_78772 == 32'h0000_0007 ? array_update_79445 : array_update_79435[7];
  assign array_update_79446[8] = add_78772 == 32'h0000_0008 ? array_update_79445 : array_update_79435[8];
  assign array_update_79446[9] = add_78772 == 32'h0000_0009 ? array_update_79445 : array_update_79435[9];
  assign array_index_79448 = array_update_79446[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign add_79450 = add_79315 + 32'h0000_0001;
  assign array_update_79451[0] = add_79450 == 32'h0000_0000 ? 32'h0000_0000 : array_index_79448[0];
  assign array_update_79451[1] = add_79450 == 32'h0000_0001 ? 32'h0000_0000 : array_index_79448[1];
  assign array_update_79451[2] = add_79450 == 32'h0000_0002 ? 32'h0000_0000 : array_index_79448[2];
  assign array_update_79451[3] = add_79450 == 32'h0000_0003 ? 32'h0000_0000 : array_index_79448[3];
  assign array_update_79451[4] = add_79450 == 32'h0000_0004 ? 32'h0000_0000 : array_index_79448[4];
  assign array_update_79451[5] = add_79450 == 32'h0000_0005 ? 32'h0000_0000 : array_index_79448[5];
  assign array_update_79451[6] = add_79450 == 32'h0000_0006 ? 32'h0000_0000 : array_index_79448[6];
  assign array_update_79451[7] = add_79450 == 32'h0000_0007 ? 32'h0000_0000 : array_index_79448[7];
  assign array_update_79451[8] = add_79450 == 32'h0000_0008 ? 32'h0000_0000 : array_index_79448[8];
  assign array_update_79451[9] = add_79450 == 32'h0000_0009 ? 32'h0000_0000 : array_index_79448[9];
  assign literal_79452 = 32'h0000_0000;
  assign array_update_79453[0] = add_78772 == 32'h0000_0000 ? array_update_79451 : array_update_79446[0];
  assign array_update_79453[1] = add_78772 == 32'h0000_0001 ? array_update_79451 : array_update_79446[1];
  assign array_update_79453[2] = add_78772 == 32'h0000_0002 ? array_update_79451 : array_update_79446[2];
  assign array_update_79453[3] = add_78772 == 32'h0000_0003 ? array_update_79451 : array_update_79446[3];
  assign array_update_79453[4] = add_78772 == 32'h0000_0004 ? array_update_79451 : array_update_79446[4];
  assign array_update_79453[5] = add_78772 == 32'h0000_0005 ? array_update_79451 : array_update_79446[5];
  assign array_update_79453[6] = add_78772 == 32'h0000_0006 ? array_update_79451 : array_update_79446[6];
  assign array_update_79453[7] = add_78772 == 32'h0000_0007 ? array_update_79451 : array_update_79446[7];
  assign array_update_79453[8] = add_78772 == 32'h0000_0008 ? array_update_79451 : array_update_79446[8];
  assign array_update_79453[9] = add_78772 == 32'h0000_0009 ? array_update_79451 : array_update_79446[9];
  assign array_index_79455 = array_update_72021[literal_79452 > 32'h0000_0009 ? 4'h9 : literal_79452[3:0]];
  assign array_index_79456 = array_update_79453[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_79460 = smul32b_32b_x_32b(array_index_78779[literal_79452 > 32'h0000_0009 ? 4'h9 : literal_79452[3:0]], array_index_79455[add_79450 > 32'h0000_0009 ? 4'h9 : add_79450[3:0]]);
  assign add_79462 = array_index_79456[add_79450 > 32'h0000_0009 ? 4'h9 : add_79450[3:0]] + smul_79460;
  assign array_update_79464[0] = add_79450 == 32'h0000_0000 ? add_79462 : array_index_79456[0];
  assign array_update_79464[1] = add_79450 == 32'h0000_0001 ? add_79462 : array_index_79456[1];
  assign array_update_79464[2] = add_79450 == 32'h0000_0002 ? add_79462 : array_index_79456[2];
  assign array_update_79464[3] = add_79450 == 32'h0000_0003 ? add_79462 : array_index_79456[3];
  assign array_update_79464[4] = add_79450 == 32'h0000_0004 ? add_79462 : array_index_79456[4];
  assign array_update_79464[5] = add_79450 == 32'h0000_0005 ? add_79462 : array_index_79456[5];
  assign array_update_79464[6] = add_79450 == 32'h0000_0006 ? add_79462 : array_index_79456[6];
  assign array_update_79464[7] = add_79450 == 32'h0000_0007 ? add_79462 : array_index_79456[7];
  assign array_update_79464[8] = add_79450 == 32'h0000_0008 ? add_79462 : array_index_79456[8];
  assign array_update_79464[9] = add_79450 == 32'h0000_0009 ? add_79462 : array_index_79456[9];
  assign add_79465 = literal_79452 + 32'h0000_0001;
  assign array_update_79466[0] = add_78772 == 32'h0000_0000 ? array_update_79464 : array_update_79453[0];
  assign array_update_79466[1] = add_78772 == 32'h0000_0001 ? array_update_79464 : array_update_79453[1];
  assign array_update_79466[2] = add_78772 == 32'h0000_0002 ? array_update_79464 : array_update_79453[2];
  assign array_update_79466[3] = add_78772 == 32'h0000_0003 ? array_update_79464 : array_update_79453[3];
  assign array_update_79466[4] = add_78772 == 32'h0000_0004 ? array_update_79464 : array_update_79453[4];
  assign array_update_79466[5] = add_78772 == 32'h0000_0005 ? array_update_79464 : array_update_79453[5];
  assign array_update_79466[6] = add_78772 == 32'h0000_0006 ? array_update_79464 : array_update_79453[6];
  assign array_update_79466[7] = add_78772 == 32'h0000_0007 ? array_update_79464 : array_update_79453[7];
  assign array_update_79466[8] = add_78772 == 32'h0000_0008 ? array_update_79464 : array_update_79453[8];
  assign array_update_79466[9] = add_78772 == 32'h0000_0009 ? array_update_79464 : array_update_79453[9];
  assign array_index_79468 = array_update_72021[add_79465 > 32'h0000_0009 ? 4'h9 : add_79465[3:0]];
  assign array_index_79469 = array_update_79466[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_79473 = smul32b_32b_x_32b(array_index_78779[add_79465 > 32'h0000_0009 ? 4'h9 : add_79465[3:0]], array_index_79468[add_79450 > 32'h0000_0009 ? 4'h9 : add_79450[3:0]]);
  assign add_79475 = array_index_79469[add_79450 > 32'h0000_0009 ? 4'h9 : add_79450[3:0]] + smul_79473;
  assign array_update_79477[0] = add_79450 == 32'h0000_0000 ? add_79475 : array_index_79469[0];
  assign array_update_79477[1] = add_79450 == 32'h0000_0001 ? add_79475 : array_index_79469[1];
  assign array_update_79477[2] = add_79450 == 32'h0000_0002 ? add_79475 : array_index_79469[2];
  assign array_update_79477[3] = add_79450 == 32'h0000_0003 ? add_79475 : array_index_79469[3];
  assign array_update_79477[4] = add_79450 == 32'h0000_0004 ? add_79475 : array_index_79469[4];
  assign array_update_79477[5] = add_79450 == 32'h0000_0005 ? add_79475 : array_index_79469[5];
  assign array_update_79477[6] = add_79450 == 32'h0000_0006 ? add_79475 : array_index_79469[6];
  assign array_update_79477[7] = add_79450 == 32'h0000_0007 ? add_79475 : array_index_79469[7];
  assign array_update_79477[8] = add_79450 == 32'h0000_0008 ? add_79475 : array_index_79469[8];
  assign array_update_79477[9] = add_79450 == 32'h0000_0009 ? add_79475 : array_index_79469[9];
  assign add_79478 = add_79465 + 32'h0000_0001;
  assign array_update_79479[0] = add_78772 == 32'h0000_0000 ? array_update_79477 : array_update_79466[0];
  assign array_update_79479[1] = add_78772 == 32'h0000_0001 ? array_update_79477 : array_update_79466[1];
  assign array_update_79479[2] = add_78772 == 32'h0000_0002 ? array_update_79477 : array_update_79466[2];
  assign array_update_79479[3] = add_78772 == 32'h0000_0003 ? array_update_79477 : array_update_79466[3];
  assign array_update_79479[4] = add_78772 == 32'h0000_0004 ? array_update_79477 : array_update_79466[4];
  assign array_update_79479[5] = add_78772 == 32'h0000_0005 ? array_update_79477 : array_update_79466[5];
  assign array_update_79479[6] = add_78772 == 32'h0000_0006 ? array_update_79477 : array_update_79466[6];
  assign array_update_79479[7] = add_78772 == 32'h0000_0007 ? array_update_79477 : array_update_79466[7];
  assign array_update_79479[8] = add_78772 == 32'h0000_0008 ? array_update_79477 : array_update_79466[8];
  assign array_update_79479[9] = add_78772 == 32'h0000_0009 ? array_update_79477 : array_update_79466[9];
  assign array_index_79481 = array_update_72021[add_79478 > 32'h0000_0009 ? 4'h9 : add_79478[3:0]];
  assign array_index_79482 = array_update_79479[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_79486 = smul32b_32b_x_32b(array_index_78779[add_79478 > 32'h0000_0009 ? 4'h9 : add_79478[3:0]], array_index_79481[add_79450 > 32'h0000_0009 ? 4'h9 : add_79450[3:0]]);
  assign add_79488 = array_index_79482[add_79450 > 32'h0000_0009 ? 4'h9 : add_79450[3:0]] + smul_79486;
  assign array_update_79490[0] = add_79450 == 32'h0000_0000 ? add_79488 : array_index_79482[0];
  assign array_update_79490[1] = add_79450 == 32'h0000_0001 ? add_79488 : array_index_79482[1];
  assign array_update_79490[2] = add_79450 == 32'h0000_0002 ? add_79488 : array_index_79482[2];
  assign array_update_79490[3] = add_79450 == 32'h0000_0003 ? add_79488 : array_index_79482[3];
  assign array_update_79490[4] = add_79450 == 32'h0000_0004 ? add_79488 : array_index_79482[4];
  assign array_update_79490[5] = add_79450 == 32'h0000_0005 ? add_79488 : array_index_79482[5];
  assign array_update_79490[6] = add_79450 == 32'h0000_0006 ? add_79488 : array_index_79482[6];
  assign array_update_79490[7] = add_79450 == 32'h0000_0007 ? add_79488 : array_index_79482[7];
  assign array_update_79490[8] = add_79450 == 32'h0000_0008 ? add_79488 : array_index_79482[8];
  assign array_update_79490[9] = add_79450 == 32'h0000_0009 ? add_79488 : array_index_79482[9];
  assign add_79491 = add_79478 + 32'h0000_0001;
  assign array_update_79492[0] = add_78772 == 32'h0000_0000 ? array_update_79490 : array_update_79479[0];
  assign array_update_79492[1] = add_78772 == 32'h0000_0001 ? array_update_79490 : array_update_79479[1];
  assign array_update_79492[2] = add_78772 == 32'h0000_0002 ? array_update_79490 : array_update_79479[2];
  assign array_update_79492[3] = add_78772 == 32'h0000_0003 ? array_update_79490 : array_update_79479[3];
  assign array_update_79492[4] = add_78772 == 32'h0000_0004 ? array_update_79490 : array_update_79479[4];
  assign array_update_79492[5] = add_78772 == 32'h0000_0005 ? array_update_79490 : array_update_79479[5];
  assign array_update_79492[6] = add_78772 == 32'h0000_0006 ? array_update_79490 : array_update_79479[6];
  assign array_update_79492[7] = add_78772 == 32'h0000_0007 ? array_update_79490 : array_update_79479[7];
  assign array_update_79492[8] = add_78772 == 32'h0000_0008 ? array_update_79490 : array_update_79479[8];
  assign array_update_79492[9] = add_78772 == 32'h0000_0009 ? array_update_79490 : array_update_79479[9];
  assign array_index_79494 = array_update_72021[add_79491 > 32'h0000_0009 ? 4'h9 : add_79491[3:0]];
  assign array_index_79495 = array_update_79492[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_79499 = smul32b_32b_x_32b(array_index_78779[add_79491 > 32'h0000_0009 ? 4'h9 : add_79491[3:0]], array_index_79494[add_79450 > 32'h0000_0009 ? 4'h9 : add_79450[3:0]]);
  assign add_79501 = array_index_79495[add_79450 > 32'h0000_0009 ? 4'h9 : add_79450[3:0]] + smul_79499;
  assign array_update_79503[0] = add_79450 == 32'h0000_0000 ? add_79501 : array_index_79495[0];
  assign array_update_79503[1] = add_79450 == 32'h0000_0001 ? add_79501 : array_index_79495[1];
  assign array_update_79503[2] = add_79450 == 32'h0000_0002 ? add_79501 : array_index_79495[2];
  assign array_update_79503[3] = add_79450 == 32'h0000_0003 ? add_79501 : array_index_79495[3];
  assign array_update_79503[4] = add_79450 == 32'h0000_0004 ? add_79501 : array_index_79495[4];
  assign array_update_79503[5] = add_79450 == 32'h0000_0005 ? add_79501 : array_index_79495[5];
  assign array_update_79503[6] = add_79450 == 32'h0000_0006 ? add_79501 : array_index_79495[6];
  assign array_update_79503[7] = add_79450 == 32'h0000_0007 ? add_79501 : array_index_79495[7];
  assign array_update_79503[8] = add_79450 == 32'h0000_0008 ? add_79501 : array_index_79495[8];
  assign array_update_79503[9] = add_79450 == 32'h0000_0009 ? add_79501 : array_index_79495[9];
  assign add_79504 = add_79491 + 32'h0000_0001;
  assign array_update_79505[0] = add_78772 == 32'h0000_0000 ? array_update_79503 : array_update_79492[0];
  assign array_update_79505[1] = add_78772 == 32'h0000_0001 ? array_update_79503 : array_update_79492[1];
  assign array_update_79505[2] = add_78772 == 32'h0000_0002 ? array_update_79503 : array_update_79492[2];
  assign array_update_79505[3] = add_78772 == 32'h0000_0003 ? array_update_79503 : array_update_79492[3];
  assign array_update_79505[4] = add_78772 == 32'h0000_0004 ? array_update_79503 : array_update_79492[4];
  assign array_update_79505[5] = add_78772 == 32'h0000_0005 ? array_update_79503 : array_update_79492[5];
  assign array_update_79505[6] = add_78772 == 32'h0000_0006 ? array_update_79503 : array_update_79492[6];
  assign array_update_79505[7] = add_78772 == 32'h0000_0007 ? array_update_79503 : array_update_79492[7];
  assign array_update_79505[8] = add_78772 == 32'h0000_0008 ? array_update_79503 : array_update_79492[8];
  assign array_update_79505[9] = add_78772 == 32'h0000_0009 ? array_update_79503 : array_update_79492[9];
  assign array_index_79507 = array_update_72021[add_79504 > 32'h0000_0009 ? 4'h9 : add_79504[3:0]];
  assign array_index_79508 = array_update_79505[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_79512 = smul32b_32b_x_32b(array_index_78779[add_79504 > 32'h0000_0009 ? 4'h9 : add_79504[3:0]], array_index_79507[add_79450 > 32'h0000_0009 ? 4'h9 : add_79450[3:0]]);
  assign add_79514 = array_index_79508[add_79450 > 32'h0000_0009 ? 4'h9 : add_79450[3:0]] + smul_79512;
  assign array_update_79516[0] = add_79450 == 32'h0000_0000 ? add_79514 : array_index_79508[0];
  assign array_update_79516[1] = add_79450 == 32'h0000_0001 ? add_79514 : array_index_79508[1];
  assign array_update_79516[2] = add_79450 == 32'h0000_0002 ? add_79514 : array_index_79508[2];
  assign array_update_79516[3] = add_79450 == 32'h0000_0003 ? add_79514 : array_index_79508[3];
  assign array_update_79516[4] = add_79450 == 32'h0000_0004 ? add_79514 : array_index_79508[4];
  assign array_update_79516[5] = add_79450 == 32'h0000_0005 ? add_79514 : array_index_79508[5];
  assign array_update_79516[6] = add_79450 == 32'h0000_0006 ? add_79514 : array_index_79508[6];
  assign array_update_79516[7] = add_79450 == 32'h0000_0007 ? add_79514 : array_index_79508[7];
  assign array_update_79516[8] = add_79450 == 32'h0000_0008 ? add_79514 : array_index_79508[8];
  assign array_update_79516[9] = add_79450 == 32'h0000_0009 ? add_79514 : array_index_79508[9];
  assign add_79517 = add_79504 + 32'h0000_0001;
  assign array_update_79518[0] = add_78772 == 32'h0000_0000 ? array_update_79516 : array_update_79505[0];
  assign array_update_79518[1] = add_78772 == 32'h0000_0001 ? array_update_79516 : array_update_79505[1];
  assign array_update_79518[2] = add_78772 == 32'h0000_0002 ? array_update_79516 : array_update_79505[2];
  assign array_update_79518[3] = add_78772 == 32'h0000_0003 ? array_update_79516 : array_update_79505[3];
  assign array_update_79518[4] = add_78772 == 32'h0000_0004 ? array_update_79516 : array_update_79505[4];
  assign array_update_79518[5] = add_78772 == 32'h0000_0005 ? array_update_79516 : array_update_79505[5];
  assign array_update_79518[6] = add_78772 == 32'h0000_0006 ? array_update_79516 : array_update_79505[6];
  assign array_update_79518[7] = add_78772 == 32'h0000_0007 ? array_update_79516 : array_update_79505[7];
  assign array_update_79518[8] = add_78772 == 32'h0000_0008 ? array_update_79516 : array_update_79505[8];
  assign array_update_79518[9] = add_78772 == 32'h0000_0009 ? array_update_79516 : array_update_79505[9];
  assign array_index_79520 = array_update_72021[add_79517 > 32'h0000_0009 ? 4'h9 : add_79517[3:0]];
  assign array_index_79521 = array_update_79518[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_79525 = smul32b_32b_x_32b(array_index_78779[add_79517 > 32'h0000_0009 ? 4'h9 : add_79517[3:0]], array_index_79520[add_79450 > 32'h0000_0009 ? 4'h9 : add_79450[3:0]]);
  assign add_79527 = array_index_79521[add_79450 > 32'h0000_0009 ? 4'h9 : add_79450[3:0]] + smul_79525;
  assign array_update_79529[0] = add_79450 == 32'h0000_0000 ? add_79527 : array_index_79521[0];
  assign array_update_79529[1] = add_79450 == 32'h0000_0001 ? add_79527 : array_index_79521[1];
  assign array_update_79529[2] = add_79450 == 32'h0000_0002 ? add_79527 : array_index_79521[2];
  assign array_update_79529[3] = add_79450 == 32'h0000_0003 ? add_79527 : array_index_79521[3];
  assign array_update_79529[4] = add_79450 == 32'h0000_0004 ? add_79527 : array_index_79521[4];
  assign array_update_79529[5] = add_79450 == 32'h0000_0005 ? add_79527 : array_index_79521[5];
  assign array_update_79529[6] = add_79450 == 32'h0000_0006 ? add_79527 : array_index_79521[6];
  assign array_update_79529[7] = add_79450 == 32'h0000_0007 ? add_79527 : array_index_79521[7];
  assign array_update_79529[8] = add_79450 == 32'h0000_0008 ? add_79527 : array_index_79521[8];
  assign array_update_79529[9] = add_79450 == 32'h0000_0009 ? add_79527 : array_index_79521[9];
  assign add_79530 = add_79517 + 32'h0000_0001;
  assign array_update_79531[0] = add_78772 == 32'h0000_0000 ? array_update_79529 : array_update_79518[0];
  assign array_update_79531[1] = add_78772 == 32'h0000_0001 ? array_update_79529 : array_update_79518[1];
  assign array_update_79531[2] = add_78772 == 32'h0000_0002 ? array_update_79529 : array_update_79518[2];
  assign array_update_79531[3] = add_78772 == 32'h0000_0003 ? array_update_79529 : array_update_79518[3];
  assign array_update_79531[4] = add_78772 == 32'h0000_0004 ? array_update_79529 : array_update_79518[4];
  assign array_update_79531[5] = add_78772 == 32'h0000_0005 ? array_update_79529 : array_update_79518[5];
  assign array_update_79531[6] = add_78772 == 32'h0000_0006 ? array_update_79529 : array_update_79518[6];
  assign array_update_79531[7] = add_78772 == 32'h0000_0007 ? array_update_79529 : array_update_79518[7];
  assign array_update_79531[8] = add_78772 == 32'h0000_0008 ? array_update_79529 : array_update_79518[8];
  assign array_update_79531[9] = add_78772 == 32'h0000_0009 ? array_update_79529 : array_update_79518[9];
  assign array_index_79533 = array_update_72021[add_79530 > 32'h0000_0009 ? 4'h9 : add_79530[3:0]];
  assign array_index_79534 = array_update_79531[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_79538 = smul32b_32b_x_32b(array_index_78779[add_79530 > 32'h0000_0009 ? 4'h9 : add_79530[3:0]], array_index_79533[add_79450 > 32'h0000_0009 ? 4'h9 : add_79450[3:0]]);
  assign add_79540 = array_index_79534[add_79450 > 32'h0000_0009 ? 4'h9 : add_79450[3:0]] + smul_79538;
  assign array_update_79542[0] = add_79450 == 32'h0000_0000 ? add_79540 : array_index_79534[0];
  assign array_update_79542[1] = add_79450 == 32'h0000_0001 ? add_79540 : array_index_79534[1];
  assign array_update_79542[2] = add_79450 == 32'h0000_0002 ? add_79540 : array_index_79534[2];
  assign array_update_79542[3] = add_79450 == 32'h0000_0003 ? add_79540 : array_index_79534[3];
  assign array_update_79542[4] = add_79450 == 32'h0000_0004 ? add_79540 : array_index_79534[4];
  assign array_update_79542[5] = add_79450 == 32'h0000_0005 ? add_79540 : array_index_79534[5];
  assign array_update_79542[6] = add_79450 == 32'h0000_0006 ? add_79540 : array_index_79534[6];
  assign array_update_79542[7] = add_79450 == 32'h0000_0007 ? add_79540 : array_index_79534[7];
  assign array_update_79542[8] = add_79450 == 32'h0000_0008 ? add_79540 : array_index_79534[8];
  assign array_update_79542[9] = add_79450 == 32'h0000_0009 ? add_79540 : array_index_79534[9];
  assign add_79543 = add_79530 + 32'h0000_0001;
  assign array_update_79544[0] = add_78772 == 32'h0000_0000 ? array_update_79542 : array_update_79531[0];
  assign array_update_79544[1] = add_78772 == 32'h0000_0001 ? array_update_79542 : array_update_79531[1];
  assign array_update_79544[2] = add_78772 == 32'h0000_0002 ? array_update_79542 : array_update_79531[2];
  assign array_update_79544[3] = add_78772 == 32'h0000_0003 ? array_update_79542 : array_update_79531[3];
  assign array_update_79544[4] = add_78772 == 32'h0000_0004 ? array_update_79542 : array_update_79531[4];
  assign array_update_79544[5] = add_78772 == 32'h0000_0005 ? array_update_79542 : array_update_79531[5];
  assign array_update_79544[6] = add_78772 == 32'h0000_0006 ? array_update_79542 : array_update_79531[6];
  assign array_update_79544[7] = add_78772 == 32'h0000_0007 ? array_update_79542 : array_update_79531[7];
  assign array_update_79544[8] = add_78772 == 32'h0000_0008 ? array_update_79542 : array_update_79531[8];
  assign array_update_79544[9] = add_78772 == 32'h0000_0009 ? array_update_79542 : array_update_79531[9];
  assign array_index_79546 = array_update_72021[add_79543 > 32'h0000_0009 ? 4'h9 : add_79543[3:0]];
  assign array_index_79547 = array_update_79544[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_79551 = smul32b_32b_x_32b(array_index_78779[add_79543 > 32'h0000_0009 ? 4'h9 : add_79543[3:0]], array_index_79546[add_79450 > 32'h0000_0009 ? 4'h9 : add_79450[3:0]]);
  assign add_79553 = array_index_79547[add_79450 > 32'h0000_0009 ? 4'h9 : add_79450[3:0]] + smul_79551;
  assign array_update_79555[0] = add_79450 == 32'h0000_0000 ? add_79553 : array_index_79547[0];
  assign array_update_79555[1] = add_79450 == 32'h0000_0001 ? add_79553 : array_index_79547[1];
  assign array_update_79555[2] = add_79450 == 32'h0000_0002 ? add_79553 : array_index_79547[2];
  assign array_update_79555[3] = add_79450 == 32'h0000_0003 ? add_79553 : array_index_79547[3];
  assign array_update_79555[4] = add_79450 == 32'h0000_0004 ? add_79553 : array_index_79547[4];
  assign array_update_79555[5] = add_79450 == 32'h0000_0005 ? add_79553 : array_index_79547[5];
  assign array_update_79555[6] = add_79450 == 32'h0000_0006 ? add_79553 : array_index_79547[6];
  assign array_update_79555[7] = add_79450 == 32'h0000_0007 ? add_79553 : array_index_79547[7];
  assign array_update_79555[8] = add_79450 == 32'h0000_0008 ? add_79553 : array_index_79547[8];
  assign array_update_79555[9] = add_79450 == 32'h0000_0009 ? add_79553 : array_index_79547[9];
  assign add_79556 = add_79543 + 32'h0000_0001;
  assign array_update_79557[0] = add_78772 == 32'h0000_0000 ? array_update_79555 : array_update_79544[0];
  assign array_update_79557[1] = add_78772 == 32'h0000_0001 ? array_update_79555 : array_update_79544[1];
  assign array_update_79557[2] = add_78772 == 32'h0000_0002 ? array_update_79555 : array_update_79544[2];
  assign array_update_79557[3] = add_78772 == 32'h0000_0003 ? array_update_79555 : array_update_79544[3];
  assign array_update_79557[4] = add_78772 == 32'h0000_0004 ? array_update_79555 : array_update_79544[4];
  assign array_update_79557[5] = add_78772 == 32'h0000_0005 ? array_update_79555 : array_update_79544[5];
  assign array_update_79557[6] = add_78772 == 32'h0000_0006 ? array_update_79555 : array_update_79544[6];
  assign array_update_79557[7] = add_78772 == 32'h0000_0007 ? array_update_79555 : array_update_79544[7];
  assign array_update_79557[8] = add_78772 == 32'h0000_0008 ? array_update_79555 : array_update_79544[8];
  assign array_update_79557[9] = add_78772 == 32'h0000_0009 ? array_update_79555 : array_update_79544[9];
  assign array_index_79559 = array_update_72021[add_79556 > 32'h0000_0009 ? 4'h9 : add_79556[3:0]];
  assign array_index_79560 = array_update_79557[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_79564 = smul32b_32b_x_32b(array_index_78779[add_79556 > 32'h0000_0009 ? 4'h9 : add_79556[3:0]], array_index_79559[add_79450 > 32'h0000_0009 ? 4'h9 : add_79450[3:0]]);
  assign add_79566 = array_index_79560[add_79450 > 32'h0000_0009 ? 4'h9 : add_79450[3:0]] + smul_79564;
  assign array_update_79568[0] = add_79450 == 32'h0000_0000 ? add_79566 : array_index_79560[0];
  assign array_update_79568[1] = add_79450 == 32'h0000_0001 ? add_79566 : array_index_79560[1];
  assign array_update_79568[2] = add_79450 == 32'h0000_0002 ? add_79566 : array_index_79560[2];
  assign array_update_79568[3] = add_79450 == 32'h0000_0003 ? add_79566 : array_index_79560[3];
  assign array_update_79568[4] = add_79450 == 32'h0000_0004 ? add_79566 : array_index_79560[4];
  assign array_update_79568[5] = add_79450 == 32'h0000_0005 ? add_79566 : array_index_79560[5];
  assign array_update_79568[6] = add_79450 == 32'h0000_0006 ? add_79566 : array_index_79560[6];
  assign array_update_79568[7] = add_79450 == 32'h0000_0007 ? add_79566 : array_index_79560[7];
  assign array_update_79568[8] = add_79450 == 32'h0000_0008 ? add_79566 : array_index_79560[8];
  assign array_update_79568[9] = add_79450 == 32'h0000_0009 ? add_79566 : array_index_79560[9];
  assign add_79569 = add_79556 + 32'h0000_0001;
  assign array_update_79570[0] = add_78772 == 32'h0000_0000 ? array_update_79568 : array_update_79557[0];
  assign array_update_79570[1] = add_78772 == 32'h0000_0001 ? array_update_79568 : array_update_79557[1];
  assign array_update_79570[2] = add_78772 == 32'h0000_0002 ? array_update_79568 : array_update_79557[2];
  assign array_update_79570[3] = add_78772 == 32'h0000_0003 ? array_update_79568 : array_update_79557[3];
  assign array_update_79570[4] = add_78772 == 32'h0000_0004 ? array_update_79568 : array_update_79557[4];
  assign array_update_79570[5] = add_78772 == 32'h0000_0005 ? array_update_79568 : array_update_79557[5];
  assign array_update_79570[6] = add_78772 == 32'h0000_0006 ? array_update_79568 : array_update_79557[6];
  assign array_update_79570[7] = add_78772 == 32'h0000_0007 ? array_update_79568 : array_update_79557[7];
  assign array_update_79570[8] = add_78772 == 32'h0000_0008 ? array_update_79568 : array_update_79557[8];
  assign array_update_79570[9] = add_78772 == 32'h0000_0009 ? array_update_79568 : array_update_79557[9];
  assign array_index_79572 = array_update_72021[add_79569 > 32'h0000_0009 ? 4'h9 : add_79569[3:0]];
  assign array_index_79573 = array_update_79570[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_79577 = smul32b_32b_x_32b(array_index_78779[add_79569 > 32'h0000_0009 ? 4'h9 : add_79569[3:0]], array_index_79572[add_79450 > 32'h0000_0009 ? 4'h9 : add_79450[3:0]]);
  assign add_79579 = array_index_79573[add_79450 > 32'h0000_0009 ? 4'h9 : add_79450[3:0]] + smul_79577;
  assign array_update_79580[0] = add_79450 == 32'h0000_0000 ? add_79579 : array_index_79573[0];
  assign array_update_79580[1] = add_79450 == 32'h0000_0001 ? add_79579 : array_index_79573[1];
  assign array_update_79580[2] = add_79450 == 32'h0000_0002 ? add_79579 : array_index_79573[2];
  assign array_update_79580[3] = add_79450 == 32'h0000_0003 ? add_79579 : array_index_79573[3];
  assign array_update_79580[4] = add_79450 == 32'h0000_0004 ? add_79579 : array_index_79573[4];
  assign array_update_79580[5] = add_79450 == 32'h0000_0005 ? add_79579 : array_index_79573[5];
  assign array_update_79580[6] = add_79450 == 32'h0000_0006 ? add_79579 : array_index_79573[6];
  assign array_update_79580[7] = add_79450 == 32'h0000_0007 ? add_79579 : array_index_79573[7];
  assign array_update_79580[8] = add_79450 == 32'h0000_0008 ? add_79579 : array_index_79573[8];
  assign array_update_79580[9] = add_79450 == 32'h0000_0009 ? add_79579 : array_index_79573[9];
  assign array_update_79581[0] = add_78772 == 32'h0000_0000 ? array_update_79580 : array_update_79570[0];
  assign array_update_79581[1] = add_78772 == 32'h0000_0001 ? array_update_79580 : array_update_79570[1];
  assign array_update_79581[2] = add_78772 == 32'h0000_0002 ? array_update_79580 : array_update_79570[2];
  assign array_update_79581[3] = add_78772 == 32'h0000_0003 ? array_update_79580 : array_update_79570[3];
  assign array_update_79581[4] = add_78772 == 32'h0000_0004 ? array_update_79580 : array_update_79570[4];
  assign array_update_79581[5] = add_78772 == 32'h0000_0005 ? array_update_79580 : array_update_79570[5];
  assign array_update_79581[6] = add_78772 == 32'h0000_0006 ? array_update_79580 : array_update_79570[6];
  assign array_update_79581[7] = add_78772 == 32'h0000_0007 ? array_update_79580 : array_update_79570[7];
  assign array_update_79581[8] = add_78772 == 32'h0000_0008 ? array_update_79580 : array_update_79570[8];
  assign array_update_79581[9] = add_78772 == 32'h0000_0009 ? array_update_79580 : array_update_79570[9];
  assign array_index_79583 = array_update_79581[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign add_79585 = add_79450 + 32'h0000_0001;
  assign array_update_79586[0] = add_79585 == 32'h0000_0000 ? 32'h0000_0000 : array_index_79583[0];
  assign array_update_79586[1] = add_79585 == 32'h0000_0001 ? 32'h0000_0000 : array_index_79583[1];
  assign array_update_79586[2] = add_79585 == 32'h0000_0002 ? 32'h0000_0000 : array_index_79583[2];
  assign array_update_79586[3] = add_79585 == 32'h0000_0003 ? 32'h0000_0000 : array_index_79583[3];
  assign array_update_79586[4] = add_79585 == 32'h0000_0004 ? 32'h0000_0000 : array_index_79583[4];
  assign array_update_79586[5] = add_79585 == 32'h0000_0005 ? 32'h0000_0000 : array_index_79583[5];
  assign array_update_79586[6] = add_79585 == 32'h0000_0006 ? 32'h0000_0000 : array_index_79583[6];
  assign array_update_79586[7] = add_79585 == 32'h0000_0007 ? 32'h0000_0000 : array_index_79583[7];
  assign array_update_79586[8] = add_79585 == 32'h0000_0008 ? 32'h0000_0000 : array_index_79583[8];
  assign array_update_79586[9] = add_79585 == 32'h0000_0009 ? 32'h0000_0000 : array_index_79583[9];
  assign literal_79587 = 32'h0000_0000;
  assign array_update_79588[0] = add_78772 == 32'h0000_0000 ? array_update_79586 : array_update_79581[0];
  assign array_update_79588[1] = add_78772 == 32'h0000_0001 ? array_update_79586 : array_update_79581[1];
  assign array_update_79588[2] = add_78772 == 32'h0000_0002 ? array_update_79586 : array_update_79581[2];
  assign array_update_79588[3] = add_78772 == 32'h0000_0003 ? array_update_79586 : array_update_79581[3];
  assign array_update_79588[4] = add_78772 == 32'h0000_0004 ? array_update_79586 : array_update_79581[4];
  assign array_update_79588[5] = add_78772 == 32'h0000_0005 ? array_update_79586 : array_update_79581[5];
  assign array_update_79588[6] = add_78772 == 32'h0000_0006 ? array_update_79586 : array_update_79581[6];
  assign array_update_79588[7] = add_78772 == 32'h0000_0007 ? array_update_79586 : array_update_79581[7];
  assign array_update_79588[8] = add_78772 == 32'h0000_0008 ? array_update_79586 : array_update_79581[8];
  assign array_update_79588[9] = add_78772 == 32'h0000_0009 ? array_update_79586 : array_update_79581[9];
  assign array_index_79590 = array_update_72021[literal_79587 > 32'h0000_0009 ? 4'h9 : literal_79587[3:0]];
  assign array_index_79591 = array_update_79588[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_79595 = smul32b_32b_x_32b(array_index_78779[literal_79587 > 32'h0000_0009 ? 4'h9 : literal_79587[3:0]], array_index_79590[add_79585 > 32'h0000_0009 ? 4'h9 : add_79585[3:0]]);
  assign add_79597 = array_index_79591[add_79585 > 32'h0000_0009 ? 4'h9 : add_79585[3:0]] + smul_79595;
  assign array_update_79599[0] = add_79585 == 32'h0000_0000 ? add_79597 : array_index_79591[0];
  assign array_update_79599[1] = add_79585 == 32'h0000_0001 ? add_79597 : array_index_79591[1];
  assign array_update_79599[2] = add_79585 == 32'h0000_0002 ? add_79597 : array_index_79591[2];
  assign array_update_79599[3] = add_79585 == 32'h0000_0003 ? add_79597 : array_index_79591[3];
  assign array_update_79599[4] = add_79585 == 32'h0000_0004 ? add_79597 : array_index_79591[4];
  assign array_update_79599[5] = add_79585 == 32'h0000_0005 ? add_79597 : array_index_79591[5];
  assign array_update_79599[6] = add_79585 == 32'h0000_0006 ? add_79597 : array_index_79591[6];
  assign array_update_79599[7] = add_79585 == 32'h0000_0007 ? add_79597 : array_index_79591[7];
  assign array_update_79599[8] = add_79585 == 32'h0000_0008 ? add_79597 : array_index_79591[8];
  assign array_update_79599[9] = add_79585 == 32'h0000_0009 ? add_79597 : array_index_79591[9];
  assign add_79600 = literal_79587 + 32'h0000_0001;
  assign array_update_79601[0] = add_78772 == 32'h0000_0000 ? array_update_79599 : array_update_79588[0];
  assign array_update_79601[1] = add_78772 == 32'h0000_0001 ? array_update_79599 : array_update_79588[1];
  assign array_update_79601[2] = add_78772 == 32'h0000_0002 ? array_update_79599 : array_update_79588[2];
  assign array_update_79601[3] = add_78772 == 32'h0000_0003 ? array_update_79599 : array_update_79588[3];
  assign array_update_79601[4] = add_78772 == 32'h0000_0004 ? array_update_79599 : array_update_79588[4];
  assign array_update_79601[5] = add_78772 == 32'h0000_0005 ? array_update_79599 : array_update_79588[5];
  assign array_update_79601[6] = add_78772 == 32'h0000_0006 ? array_update_79599 : array_update_79588[6];
  assign array_update_79601[7] = add_78772 == 32'h0000_0007 ? array_update_79599 : array_update_79588[7];
  assign array_update_79601[8] = add_78772 == 32'h0000_0008 ? array_update_79599 : array_update_79588[8];
  assign array_update_79601[9] = add_78772 == 32'h0000_0009 ? array_update_79599 : array_update_79588[9];
  assign array_index_79603 = array_update_72021[add_79600 > 32'h0000_0009 ? 4'h9 : add_79600[3:0]];
  assign array_index_79604 = array_update_79601[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_79608 = smul32b_32b_x_32b(array_index_78779[add_79600 > 32'h0000_0009 ? 4'h9 : add_79600[3:0]], array_index_79603[add_79585 > 32'h0000_0009 ? 4'h9 : add_79585[3:0]]);
  assign add_79610 = array_index_79604[add_79585 > 32'h0000_0009 ? 4'h9 : add_79585[3:0]] + smul_79608;
  assign array_update_79612[0] = add_79585 == 32'h0000_0000 ? add_79610 : array_index_79604[0];
  assign array_update_79612[1] = add_79585 == 32'h0000_0001 ? add_79610 : array_index_79604[1];
  assign array_update_79612[2] = add_79585 == 32'h0000_0002 ? add_79610 : array_index_79604[2];
  assign array_update_79612[3] = add_79585 == 32'h0000_0003 ? add_79610 : array_index_79604[3];
  assign array_update_79612[4] = add_79585 == 32'h0000_0004 ? add_79610 : array_index_79604[4];
  assign array_update_79612[5] = add_79585 == 32'h0000_0005 ? add_79610 : array_index_79604[5];
  assign array_update_79612[6] = add_79585 == 32'h0000_0006 ? add_79610 : array_index_79604[6];
  assign array_update_79612[7] = add_79585 == 32'h0000_0007 ? add_79610 : array_index_79604[7];
  assign array_update_79612[8] = add_79585 == 32'h0000_0008 ? add_79610 : array_index_79604[8];
  assign array_update_79612[9] = add_79585 == 32'h0000_0009 ? add_79610 : array_index_79604[9];
  assign add_79613 = add_79600 + 32'h0000_0001;
  assign array_update_79614[0] = add_78772 == 32'h0000_0000 ? array_update_79612 : array_update_79601[0];
  assign array_update_79614[1] = add_78772 == 32'h0000_0001 ? array_update_79612 : array_update_79601[1];
  assign array_update_79614[2] = add_78772 == 32'h0000_0002 ? array_update_79612 : array_update_79601[2];
  assign array_update_79614[3] = add_78772 == 32'h0000_0003 ? array_update_79612 : array_update_79601[3];
  assign array_update_79614[4] = add_78772 == 32'h0000_0004 ? array_update_79612 : array_update_79601[4];
  assign array_update_79614[5] = add_78772 == 32'h0000_0005 ? array_update_79612 : array_update_79601[5];
  assign array_update_79614[6] = add_78772 == 32'h0000_0006 ? array_update_79612 : array_update_79601[6];
  assign array_update_79614[7] = add_78772 == 32'h0000_0007 ? array_update_79612 : array_update_79601[7];
  assign array_update_79614[8] = add_78772 == 32'h0000_0008 ? array_update_79612 : array_update_79601[8];
  assign array_update_79614[9] = add_78772 == 32'h0000_0009 ? array_update_79612 : array_update_79601[9];
  assign array_index_79616 = array_update_72021[add_79613 > 32'h0000_0009 ? 4'h9 : add_79613[3:0]];
  assign array_index_79617 = array_update_79614[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_79621 = smul32b_32b_x_32b(array_index_78779[add_79613 > 32'h0000_0009 ? 4'h9 : add_79613[3:0]], array_index_79616[add_79585 > 32'h0000_0009 ? 4'h9 : add_79585[3:0]]);
  assign add_79623 = array_index_79617[add_79585 > 32'h0000_0009 ? 4'h9 : add_79585[3:0]] + smul_79621;
  assign array_update_79625[0] = add_79585 == 32'h0000_0000 ? add_79623 : array_index_79617[0];
  assign array_update_79625[1] = add_79585 == 32'h0000_0001 ? add_79623 : array_index_79617[1];
  assign array_update_79625[2] = add_79585 == 32'h0000_0002 ? add_79623 : array_index_79617[2];
  assign array_update_79625[3] = add_79585 == 32'h0000_0003 ? add_79623 : array_index_79617[3];
  assign array_update_79625[4] = add_79585 == 32'h0000_0004 ? add_79623 : array_index_79617[4];
  assign array_update_79625[5] = add_79585 == 32'h0000_0005 ? add_79623 : array_index_79617[5];
  assign array_update_79625[6] = add_79585 == 32'h0000_0006 ? add_79623 : array_index_79617[6];
  assign array_update_79625[7] = add_79585 == 32'h0000_0007 ? add_79623 : array_index_79617[7];
  assign array_update_79625[8] = add_79585 == 32'h0000_0008 ? add_79623 : array_index_79617[8];
  assign array_update_79625[9] = add_79585 == 32'h0000_0009 ? add_79623 : array_index_79617[9];
  assign add_79626 = add_79613 + 32'h0000_0001;
  assign array_update_79627[0] = add_78772 == 32'h0000_0000 ? array_update_79625 : array_update_79614[0];
  assign array_update_79627[1] = add_78772 == 32'h0000_0001 ? array_update_79625 : array_update_79614[1];
  assign array_update_79627[2] = add_78772 == 32'h0000_0002 ? array_update_79625 : array_update_79614[2];
  assign array_update_79627[3] = add_78772 == 32'h0000_0003 ? array_update_79625 : array_update_79614[3];
  assign array_update_79627[4] = add_78772 == 32'h0000_0004 ? array_update_79625 : array_update_79614[4];
  assign array_update_79627[5] = add_78772 == 32'h0000_0005 ? array_update_79625 : array_update_79614[5];
  assign array_update_79627[6] = add_78772 == 32'h0000_0006 ? array_update_79625 : array_update_79614[6];
  assign array_update_79627[7] = add_78772 == 32'h0000_0007 ? array_update_79625 : array_update_79614[7];
  assign array_update_79627[8] = add_78772 == 32'h0000_0008 ? array_update_79625 : array_update_79614[8];
  assign array_update_79627[9] = add_78772 == 32'h0000_0009 ? array_update_79625 : array_update_79614[9];
  assign array_index_79629 = array_update_72021[add_79626 > 32'h0000_0009 ? 4'h9 : add_79626[3:0]];
  assign array_index_79630 = array_update_79627[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_79634 = smul32b_32b_x_32b(array_index_78779[add_79626 > 32'h0000_0009 ? 4'h9 : add_79626[3:0]], array_index_79629[add_79585 > 32'h0000_0009 ? 4'h9 : add_79585[3:0]]);
  assign add_79636 = array_index_79630[add_79585 > 32'h0000_0009 ? 4'h9 : add_79585[3:0]] + smul_79634;
  assign array_update_79638[0] = add_79585 == 32'h0000_0000 ? add_79636 : array_index_79630[0];
  assign array_update_79638[1] = add_79585 == 32'h0000_0001 ? add_79636 : array_index_79630[1];
  assign array_update_79638[2] = add_79585 == 32'h0000_0002 ? add_79636 : array_index_79630[2];
  assign array_update_79638[3] = add_79585 == 32'h0000_0003 ? add_79636 : array_index_79630[3];
  assign array_update_79638[4] = add_79585 == 32'h0000_0004 ? add_79636 : array_index_79630[4];
  assign array_update_79638[5] = add_79585 == 32'h0000_0005 ? add_79636 : array_index_79630[5];
  assign array_update_79638[6] = add_79585 == 32'h0000_0006 ? add_79636 : array_index_79630[6];
  assign array_update_79638[7] = add_79585 == 32'h0000_0007 ? add_79636 : array_index_79630[7];
  assign array_update_79638[8] = add_79585 == 32'h0000_0008 ? add_79636 : array_index_79630[8];
  assign array_update_79638[9] = add_79585 == 32'h0000_0009 ? add_79636 : array_index_79630[9];
  assign add_79639 = add_79626 + 32'h0000_0001;
  assign array_update_79640[0] = add_78772 == 32'h0000_0000 ? array_update_79638 : array_update_79627[0];
  assign array_update_79640[1] = add_78772 == 32'h0000_0001 ? array_update_79638 : array_update_79627[1];
  assign array_update_79640[2] = add_78772 == 32'h0000_0002 ? array_update_79638 : array_update_79627[2];
  assign array_update_79640[3] = add_78772 == 32'h0000_0003 ? array_update_79638 : array_update_79627[3];
  assign array_update_79640[4] = add_78772 == 32'h0000_0004 ? array_update_79638 : array_update_79627[4];
  assign array_update_79640[5] = add_78772 == 32'h0000_0005 ? array_update_79638 : array_update_79627[5];
  assign array_update_79640[6] = add_78772 == 32'h0000_0006 ? array_update_79638 : array_update_79627[6];
  assign array_update_79640[7] = add_78772 == 32'h0000_0007 ? array_update_79638 : array_update_79627[7];
  assign array_update_79640[8] = add_78772 == 32'h0000_0008 ? array_update_79638 : array_update_79627[8];
  assign array_update_79640[9] = add_78772 == 32'h0000_0009 ? array_update_79638 : array_update_79627[9];
  assign array_index_79642 = array_update_72021[add_79639 > 32'h0000_0009 ? 4'h9 : add_79639[3:0]];
  assign array_index_79643 = array_update_79640[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_79647 = smul32b_32b_x_32b(array_index_78779[add_79639 > 32'h0000_0009 ? 4'h9 : add_79639[3:0]], array_index_79642[add_79585 > 32'h0000_0009 ? 4'h9 : add_79585[3:0]]);
  assign add_79649 = array_index_79643[add_79585 > 32'h0000_0009 ? 4'h9 : add_79585[3:0]] + smul_79647;
  assign array_update_79651[0] = add_79585 == 32'h0000_0000 ? add_79649 : array_index_79643[0];
  assign array_update_79651[1] = add_79585 == 32'h0000_0001 ? add_79649 : array_index_79643[1];
  assign array_update_79651[2] = add_79585 == 32'h0000_0002 ? add_79649 : array_index_79643[2];
  assign array_update_79651[3] = add_79585 == 32'h0000_0003 ? add_79649 : array_index_79643[3];
  assign array_update_79651[4] = add_79585 == 32'h0000_0004 ? add_79649 : array_index_79643[4];
  assign array_update_79651[5] = add_79585 == 32'h0000_0005 ? add_79649 : array_index_79643[5];
  assign array_update_79651[6] = add_79585 == 32'h0000_0006 ? add_79649 : array_index_79643[6];
  assign array_update_79651[7] = add_79585 == 32'h0000_0007 ? add_79649 : array_index_79643[7];
  assign array_update_79651[8] = add_79585 == 32'h0000_0008 ? add_79649 : array_index_79643[8];
  assign array_update_79651[9] = add_79585 == 32'h0000_0009 ? add_79649 : array_index_79643[9];
  assign add_79652 = add_79639 + 32'h0000_0001;
  assign array_update_79653[0] = add_78772 == 32'h0000_0000 ? array_update_79651 : array_update_79640[0];
  assign array_update_79653[1] = add_78772 == 32'h0000_0001 ? array_update_79651 : array_update_79640[1];
  assign array_update_79653[2] = add_78772 == 32'h0000_0002 ? array_update_79651 : array_update_79640[2];
  assign array_update_79653[3] = add_78772 == 32'h0000_0003 ? array_update_79651 : array_update_79640[3];
  assign array_update_79653[4] = add_78772 == 32'h0000_0004 ? array_update_79651 : array_update_79640[4];
  assign array_update_79653[5] = add_78772 == 32'h0000_0005 ? array_update_79651 : array_update_79640[5];
  assign array_update_79653[6] = add_78772 == 32'h0000_0006 ? array_update_79651 : array_update_79640[6];
  assign array_update_79653[7] = add_78772 == 32'h0000_0007 ? array_update_79651 : array_update_79640[7];
  assign array_update_79653[8] = add_78772 == 32'h0000_0008 ? array_update_79651 : array_update_79640[8];
  assign array_update_79653[9] = add_78772 == 32'h0000_0009 ? array_update_79651 : array_update_79640[9];
  assign array_index_79655 = array_update_72021[add_79652 > 32'h0000_0009 ? 4'h9 : add_79652[3:0]];
  assign array_index_79656 = array_update_79653[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_79660 = smul32b_32b_x_32b(array_index_78779[add_79652 > 32'h0000_0009 ? 4'h9 : add_79652[3:0]], array_index_79655[add_79585 > 32'h0000_0009 ? 4'h9 : add_79585[3:0]]);
  assign add_79662 = array_index_79656[add_79585 > 32'h0000_0009 ? 4'h9 : add_79585[3:0]] + smul_79660;
  assign array_update_79664[0] = add_79585 == 32'h0000_0000 ? add_79662 : array_index_79656[0];
  assign array_update_79664[1] = add_79585 == 32'h0000_0001 ? add_79662 : array_index_79656[1];
  assign array_update_79664[2] = add_79585 == 32'h0000_0002 ? add_79662 : array_index_79656[2];
  assign array_update_79664[3] = add_79585 == 32'h0000_0003 ? add_79662 : array_index_79656[3];
  assign array_update_79664[4] = add_79585 == 32'h0000_0004 ? add_79662 : array_index_79656[4];
  assign array_update_79664[5] = add_79585 == 32'h0000_0005 ? add_79662 : array_index_79656[5];
  assign array_update_79664[6] = add_79585 == 32'h0000_0006 ? add_79662 : array_index_79656[6];
  assign array_update_79664[7] = add_79585 == 32'h0000_0007 ? add_79662 : array_index_79656[7];
  assign array_update_79664[8] = add_79585 == 32'h0000_0008 ? add_79662 : array_index_79656[8];
  assign array_update_79664[9] = add_79585 == 32'h0000_0009 ? add_79662 : array_index_79656[9];
  assign add_79665 = add_79652 + 32'h0000_0001;
  assign array_update_79666[0] = add_78772 == 32'h0000_0000 ? array_update_79664 : array_update_79653[0];
  assign array_update_79666[1] = add_78772 == 32'h0000_0001 ? array_update_79664 : array_update_79653[1];
  assign array_update_79666[2] = add_78772 == 32'h0000_0002 ? array_update_79664 : array_update_79653[2];
  assign array_update_79666[3] = add_78772 == 32'h0000_0003 ? array_update_79664 : array_update_79653[3];
  assign array_update_79666[4] = add_78772 == 32'h0000_0004 ? array_update_79664 : array_update_79653[4];
  assign array_update_79666[5] = add_78772 == 32'h0000_0005 ? array_update_79664 : array_update_79653[5];
  assign array_update_79666[6] = add_78772 == 32'h0000_0006 ? array_update_79664 : array_update_79653[6];
  assign array_update_79666[7] = add_78772 == 32'h0000_0007 ? array_update_79664 : array_update_79653[7];
  assign array_update_79666[8] = add_78772 == 32'h0000_0008 ? array_update_79664 : array_update_79653[8];
  assign array_update_79666[9] = add_78772 == 32'h0000_0009 ? array_update_79664 : array_update_79653[9];
  assign array_index_79668 = array_update_72021[add_79665 > 32'h0000_0009 ? 4'h9 : add_79665[3:0]];
  assign array_index_79669 = array_update_79666[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_79673 = smul32b_32b_x_32b(array_index_78779[add_79665 > 32'h0000_0009 ? 4'h9 : add_79665[3:0]], array_index_79668[add_79585 > 32'h0000_0009 ? 4'h9 : add_79585[3:0]]);
  assign add_79675 = array_index_79669[add_79585 > 32'h0000_0009 ? 4'h9 : add_79585[3:0]] + smul_79673;
  assign array_update_79677[0] = add_79585 == 32'h0000_0000 ? add_79675 : array_index_79669[0];
  assign array_update_79677[1] = add_79585 == 32'h0000_0001 ? add_79675 : array_index_79669[1];
  assign array_update_79677[2] = add_79585 == 32'h0000_0002 ? add_79675 : array_index_79669[2];
  assign array_update_79677[3] = add_79585 == 32'h0000_0003 ? add_79675 : array_index_79669[3];
  assign array_update_79677[4] = add_79585 == 32'h0000_0004 ? add_79675 : array_index_79669[4];
  assign array_update_79677[5] = add_79585 == 32'h0000_0005 ? add_79675 : array_index_79669[5];
  assign array_update_79677[6] = add_79585 == 32'h0000_0006 ? add_79675 : array_index_79669[6];
  assign array_update_79677[7] = add_79585 == 32'h0000_0007 ? add_79675 : array_index_79669[7];
  assign array_update_79677[8] = add_79585 == 32'h0000_0008 ? add_79675 : array_index_79669[8];
  assign array_update_79677[9] = add_79585 == 32'h0000_0009 ? add_79675 : array_index_79669[9];
  assign add_79678 = add_79665 + 32'h0000_0001;
  assign array_update_79679[0] = add_78772 == 32'h0000_0000 ? array_update_79677 : array_update_79666[0];
  assign array_update_79679[1] = add_78772 == 32'h0000_0001 ? array_update_79677 : array_update_79666[1];
  assign array_update_79679[2] = add_78772 == 32'h0000_0002 ? array_update_79677 : array_update_79666[2];
  assign array_update_79679[3] = add_78772 == 32'h0000_0003 ? array_update_79677 : array_update_79666[3];
  assign array_update_79679[4] = add_78772 == 32'h0000_0004 ? array_update_79677 : array_update_79666[4];
  assign array_update_79679[5] = add_78772 == 32'h0000_0005 ? array_update_79677 : array_update_79666[5];
  assign array_update_79679[6] = add_78772 == 32'h0000_0006 ? array_update_79677 : array_update_79666[6];
  assign array_update_79679[7] = add_78772 == 32'h0000_0007 ? array_update_79677 : array_update_79666[7];
  assign array_update_79679[8] = add_78772 == 32'h0000_0008 ? array_update_79677 : array_update_79666[8];
  assign array_update_79679[9] = add_78772 == 32'h0000_0009 ? array_update_79677 : array_update_79666[9];
  assign array_index_79681 = array_update_72021[add_79678 > 32'h0000_0009 ? 4'h9 : add_79678[3:0]];
  assign array_index_79682 = array_update_79679[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_79686 = smul32b_32b_x_32b(array_index_78779[add_79678 > 32'h0000_0009 ? 4'h9 : add_79678[3:0]], array_index_79681[add_79585 > 32'h0000_0009 ? 4'h9 : add_79585[3:0]]);
  assign add_79688 = array_index_79682[add_79585 > 32'h0000_0009 ? 4'h9 : add_79585[3:0]] + smul_79686;
  assign array_update_79690[0] = add_79585 == 32'h0000_0000 ? add_79688 : array_index_79682[0];
  assign array_update_79690[1] = add_79585 == 32'h0000_0001 ? add_79688 : array_index_79682[1];
  assign array_update_79690[2] = add_79585 == 32'h0000_0002 ? add_79688 : array_index_79682[2];
  assign array_update_79690[3] = add_79585 == 32'h0000_0003 ? add_79688 : array_index_79682[3];
  assign array_update_79690[4] = add_79585 == 32'h0000_0004 ? add_79688 : array_index_79682[4];
  assign array_update_79690[5] = add_79585 == 32'h0000_0005 ? add_79688 : array_index_79682[5];
  assign array_update_79690[6] = add_79585 == 32'h0000_0006 ? add_79688 : array_index_79682[6];
  assign array_update_79690[7] = add_79585 == 32'h0000_0007 ? add_79688 : array_index_79682[7];
  assign array_update_79690[8] = add_79585 == 32'h0000_0008 ? add_79688 : array_index_79682[8];
  assign array_update_79690[9] = add_79585 == 32'h0000_0009 ? add_79688 : array_index_79682[9];
  assign add_79691 = add_79678 + 32'h0000_0001;
  assign array_update_79692[0] = add_78772 == 32'h0000_0000 ? array_update_79690 : array_update_79679[0];
  assign array_update_79692[1] = add_78772 == 32'h0000_0001 ? array_update_79690 : array_update_79679[1];
  assign array_update_79692[2] = add_78772 == 32'h0000_0002 ? array_update_79690 : array_update_79679[2];
  assign array_update_79692[3] = add_78772 == 32'h0000_0003 ? array_update_79690 : array_update_79679[3];
  assign array_update_79692[4] = add_78772 == 32'h0000_0004 ? array_update_79690 : array_update_79679[4];
  assign array_update_79692[5] = add_78772 == 32'h0000_0005 ? array_update_79690 : array_update_79679[5];
  assign array_update_79692[6] = add_78772 == 32'h0000_0006 ? array_update_79690 : array_update_79679[6];
  assign array_update_79692[7] = add_78772 == 32'h0000_0007 ? array_update_79690 : array_update_79679[7];
  assign array_update_79692[8] = add_78772 == 32'h0000_0008 ? array_update_79690 : array_update_79679[8];
  assign array_update_79692[9] = add_78772 == 32'h0000_0009 ? array_update_79690 : array_update_79679[9];
  assign array_index_79694 = array_update_72021[add_79691 > 32'h0000_0009 ? 4'h9 : add_79691[3:0]];
  assign array_index_79695 = array_update_79692[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_79699 = smul32b_32b_x_32b(array_index_78779[add_79691 > 32'h0000_0009 ? 4'h9 : add_79691[3:0]], array_index_79694[add_79585 > 32'h0000_0009 ? 4'h9 : add_79585[3:0]]);
  assign add_79701 = array_index_79695[add_79585 > 32'h0000_0009 ? 4'h9 : add_79585[3:0]] + smul_79699;
  assign array_update_79703[0] = add_79585 == 32'h0000_0000 ? add_79701 : array_index_79695[0];
  assign array_update_79703[1] = add_79585 == 32'h0000_0001 ? add_79701 : array_index_79695[1];
  assign array_update_79703[2] = add_79585 == 32'h0000_0002 ? add_79701 : array_index_79695[2];
  assign array_update_79703[3] = add_79585 == 32'h0000_0003 ? add_79701 : array_index_79695[3];
  assign array_update_79703[4] = add_79585 == 32'h0000_0004 ? add_79701 : array_index_79695[4];
  assign array_update_79703[5] = add_79585 == 32'h0000_0005 ? add_79701 : array_index_79695[5];
  assign array_update_79703[6] = add_79585 == 32'h0000_0006 ? add_79701 : array_index_79695[6];
  assign array_update_79703[7] = add_79585 == 32'h0000_0007 ? add_79701 : array_index_79695[7];
  assign array_update_79703[8] = add_79585 == 32'h0000_0008 ? add_79701 : array_index_79695[8];
  assign array_update_79703[9] = add_79585 == 32'h0000_0009 ? add_79701 : array_index_79695[9];
  assign add_79704 = add_79691 + 32'h0000_0001;
  assign array_update_79705[0] = add_78772 == 32'h0000_0000 ? array_update_79703 : array_update_79692[0];
  assign array_update_79705[1] = add_78772 == 32'h0000_0001 ? array_update_79703 : array_update_79692[1];
  assign array_update_79705[2] = add_78772 == 32'h0000_0002 ? array_update_79703 : array_update_79692[2];
  assign array_update_79705[3] = add_78772 == 32'h0000_0003 ? array_update_79703 : array_update_79692[3];
  assign array_update_79705[4] = add_78772 == 32'h0000_0004 ? array_update_79703 : array_update_79692[4];
  assign array_update_79705[5] = add_78772 == 32'h0000_0005 ? array_update_79703 : array_update_79692[5];
  assign array_update_79705[6] = add_78772 == 32'h0000_0006 ? array_update_79703 : array_update_79692[6];
  assign array_update_79705[7] = add_78772 == 32'h0000_0007 ? array_update_79703 : array_update_79692[7];
  assign array_update_79705[8] = add_78772 == 32'h0000_0008 ? array_update_79703 : array_update_79692[8];
  assign array_update_79705[9] = add_78772 == 32'h0000_0009 ? array_update_79703 : array_update_79692[9];
  assign array_index_79707 = array_update_72021[add_79704 > 32'h0000_0009 ? 4'h9 : add_79704[3:0]];
  assign array_index_79708 = array_update_79705[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_79712 = smul32b_32b_x_32b(array_index_78779[add_79704 > 32'h0000_0009 ? 4'h9 : add_79704[3:0]], array_index_79707[add_79585 > 32'h0000_0009 ? 4'h9 : add_79585[3:0]]);
  assign add_79714 = array_index_79708[add_79585 > 32'h0000_0009 ? 4'h9 : add_79585[3:0]] + smul_79712;
  assign array_update_79715[0] = add_79585 == 32'h0000_0000 ? add_79714 : array_index_79708[0];
  assign array_update_79715[1] = add_79585 == 32'h0000_0001 ? add_79714 : array_index_79708[1];
  assign array_update_79715[2] = add_79585 == 32'h0000_0002 ? add_79714 : array_index_79708[2];
  assign array_update_79715[3] = add_79585 == 32'h0000_0003 ? add_79714 : array_index_79708[3];
  assign array_update_79715[4] = add_79585 == 32'h0000_0004 ? add_79714 : array_index_79708[4];
  assign array_update_79715[5] = add_79585 == 32'h0000_0005 ? add_79714 : array_index_79708[5];
  assign array_update_79715[6] = add_79585 == 32'h0000_0006 ? add_79714 : array_index_79708[6];
  assign array_update_79715[7] = add_79585 == 32'h0000_0007 ? add_79714 : array_index_79708[7];
  assign array_update_79715[8] = add_79585 == 32'h0000_0008 ? add_79714 : array_index_79708[8];
  assign array_update_79715[9] = add_79585 == 32'h0000_0009 ? add_79714 : array_index_79708[9];
  assign array_update_79716[0] = add_78772 == 32'h0000_0000 ? array_update_79715 : array_update_79705[0];
  assign array_update_79716[1] = add_78772 == 32'h0000_0001 ? array_update_79715 : array_update_79705[1];
  assign array_update_79716[2] = add_78772 == 32'h0000_0002 ? array_update_79715 : array_update_79705[2];
  assign array_update_79716[3] = add_78772 == 32'h0000_0003 ? array_update_79715 : array_update_79705[3];
  assign array_update_79716[4] = add_78772 == 32'h0000_0004 ? array_update_79715 : array_update_79705[4];
  assign array_update_79716[5] = add_78772 == 32'h0000_0005 ? array_update_79715 : array_update_79705[5];
  assign array_update_79716[6] = add_78772 == 32'h0000_0006 ? array_update_79715 : array_update_79705[6];
  assign array_update_79716[7] = add_78772 == 32'h0000_0007 ? array_update_79715 : array_update_79705[7];
  assign array_update_79716[8] = add_78772 == 32'h0000_0008 ? array_update_79715 : array_update_79705[8];
  assign array_update_79716[9] = add_78772 == 32'h0000_0009 ? array_update_79715 : array_update_79705[9];
  assign array_index_79718 = array_update_79716[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign add_79720 = add_79585 + 32'h0000_0001;
  assign array_update_79721[0] = add_79720 == 32'h0000_0000 ? 32'h0000_0000 : array_index_79718[0];
  assign array_update_79721[1] = add_79720 == 32'h0000_0001 ? 32'h0000_0000 : array_index_79718[1];
  assign array_update_79721[2] = add_79720 == 32'h0000_0002 ? 32'h0000_0000 : array_index_79718[2];
  assign array_update_79721[3] = add_79720 == 32'h0000_0003 ? 32'h0000_0000 : array_index_79718[3];
  assign array_update_79721[4] = add_79720 == 32'h0000_0004 ? 32'h0000_0000 : array_index_79718[4];
  assign array_update_79721[5] = add_79720 == 32'h0000_0005 ? 32'h0000_0000 : array_index_79718[5];
  assign array_update_79721[6] = add_79720 == 32'h0000_0006 ? 32'h0000_0000 : array_index_79718[6];
  assign array_update_79721[7] = add_79720 == 32'h0000_0007 ? 32'h0000_0000 : array_index_79718[7];
  assign array_update_79721[8] = add_79720 == 32'h0000_0008 ? 32'h0000_0000 : array_index_79718[8];
  assign array_update_79721[9] = add_79720 == 32'h0000_0009 ? 32'h0000_0000 : array_index_79718[9];
  assign literal_79722 = 32'h0000_0000;
  assign array_update_79723[0] = add_78772 == 32'h0000_0000 ? array_update_79721 : array_update_79716[0];
  assign array_update_79723[1] = add_78772 == 32'h0000_0001 ? array_update_79721 : array_update_79716[1];
  assign array_update_79723[2] = add_78772 == 32'h0000_0002 ? array_update_79721 : array_update_79716[2];
  assign array_update_79723[3] = add_78772 == 32'h0000_0003 ? array_update_79721 : array_update_79716[3];
  assign array_update_79723[4] = add_78772 == 32'h0000_0004 ? array_update_79721 : array_update_79716[4];
  assign array_update_79723[5] = add_78772 == 32'h0000_0005 ? array_update_79721 : array_update_79716[5];
  assign array_update_79723[6] = add_78772 == 32'h0000_0006 ? array_update_79721 : array_update_79716[6];
  assign array_update_79723[7] = add_78772 == 32'h0000_0007 ? array_update_79721 : array_update_79716[7];
  assign array_update_79723[8] = add_78772 == 32'h0000_0008 ? array_update_79721 : array_update_79716[8];
  assign array_update_79723[9] = add_78772 == 32'h0000_0009 ? array_update_79721 : array_update_79716[9];
  assign array_index_79725 = array_update_72021[literal_79722 > 32'h0000_0009 ? 4'h9 : literal_79722[3:0]];
  assign array_index_79726 = array_update_79723[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_79730 = smul32b_32b_x_32b(array_index_78779[literal_79722 > 32'h0000_0009 ? 4'h9 : literal_79722[3:0]], array_index_79725[add_79720 > 32'h0000_0009 ? 4'h9 : add_79720[3:0]]);
  assign add_79732 = array_index_79726[add_79720 > 32'h0000_0009 ? 4'h9 : add_79720[3:0]] + smul_79730;
  assign array_update_79734[0] = add_79720 == 32'h0000_0000 ? add_79732 : array_index_79726[0];
  assign array_update_79734[1] = add_79720 == 32'h0000_0001 ? add_79732 : array_index_79726[1];
  assign array_update_79734[2] = add_79720 == 32'h0000_0002 ? add_79732 : array_index_79726[2];
  assign array_update_79734[3] = add_79720 == 32'h0000_0003 ? add_79732 : array_index_79726[3];
  assign array_update_79734[4] = add_79720 == 32'h0000_0004 ? add_79732 : array_index_79726[4];
  assign array_update_79734[5] = add_79720 == 32'h0000_0005 ? add_79732 : array_index_79726[5];
  assign array_update_79734[6] = add_79720 == 32'h0000_0006 ? add_79732 : array_index_79726[6];
  assign array_update_79734[7] = add_79720 == 32'h0000_0007 ? add_79732 : array_index_79726[7];
  assign array_update_79734[8] = add_79720 == 32'h0000_0008 ? add_79732 : array_index_79726[8];
  assign array_update_79734[9] = add_79720 == 32'h0000_0009 ? add_79732 : array_index_79726[9];
  assign add_79735 = literal_79722 + 32'h0000_0001;
  assign array_update_79736[0] = add_78772 == 32'h0000_0000 ? array_update_79734 : array_update_79723[0];
  assign array_update_79736[1] = add_78772 == 32'h0000_0001 ? array_update_79734 : array_update_79723[1];
  assign array_update_79736[2] = add_78772 == 32'h0000_0002 ? array_update_79734 : array_update_79723[2];
  assign array_update_79736[3] = add_78772 == 32'h0000_0003 ? array_update_79734 : array_update_79723[3];
  assign array_update_79736[4] = add_78772 == 32'h0000_0004 ? array_update_79734 : array_update_79723[4];
  assign array_update_79736[5] = add_78772 == 32'h0000_0005 ? array_update_79734 : array_update_79723[5];
  assign array_update_79736[6] = add_78772 == 32'h0000_0006 ? array_update_79734 : array_update_79723[6];
  assign array_update_79736[7] = add_78772 == 32'h0000_0007 ? array_update_79734 : array_update_79723[7];
  assign array_update_79736[8] = add_78772 == 32'h0000_0008 ? array_update_79734 : array_update_79723[8];
  assign array_update_79736[9] = add_78772 == 32'h0000_0009 ? array_update_79734 : array_update_79723[9];
  assign array_index_79738 = array_update_72021[add_79735 > 32'h0000_0009 ? 4'h9 : add_79735[3:0]];
  assign array_index_79739 = array_update_79736[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_79743 = smul32b_32b_x_32b(array_index_78779[add_79735 > 32'h0000_0009 ? 4'h9 : add_79735[3:0]], array_index_79738[add_79720 > 32'h0000_0009 ? 4'h9 : add_79720[3:0]]);
  assign add_79745 = array_index_79739[add_79720 > 32'h0000_0009 ? 4'h9 : add_79720[3:0]] + smul_79743;
  assign array_update_79747[0] = add_79720 == 32'h0000_0000 ? add_79745 : array_index_79739[0];
  assign array_update_79747[1] = add_79720 == 32'h0000_0001 ? add_79745 : array_index_79739[1];
  assign array_update_79747[2] = add_79720 == 32'h0000_0002 ? add_79745 : array_index_79739[2];
  assign array_update_79747[3] = add_79720 == 32'h0000_0003 ? add_79745 : array_index_79739[3];
  assign array_update_79747[4] = add_79720 == 32'h0000_0004 ? add_79745 : array_index_79739[4];
  assign array_update_79747[5] = add_79720 == 32'h0000_0005 ? add_79745 : array_index_79739[5];
  assign array_update_79747[6] = add_79720 == 32'h0000_0006 ? add_79745 : array_index_79739[6];
  assign array_update_79747[7] = add_79720 == 32'h0000_0007 ? add_79745 : array_index_79739[7];
  assign array_update_79747[8] = add_79720 == 32'h0000_0008 ? add_79745 : array_index_79739[8];
  assign array_update_79747[9] = add_79720 == 32'h0000_0009 ? add_79745 : array_index_79739[9];
  assign add_79748 = add_79735 + 32'h0000_0001;
  assign array_update_79749[0] = add_78772 == 32'h0000_0000 ? array_update_79747 : array_update_79736[0];
  assign array_update_79749[1] = add_78772 == 32'h0000_0001 ? array_update_79747 : array_update_79736[1];
  assign array_update_79749[2] = add_78772 == 32'h0000_0002 ? array_update_79747 : array_update_79736[2];
  assign array_update_79749[3] = add_78772 == 32'h0000_0003 ? array_update_79747 : array_update_79736[3];
  assign array_update_79749[4] = add_78772 == 32'h0000_0004 ? array_update_79747 : array_update_79736[4];
  assign array_update_79749[5] = add_78772 == 32'h0000_0005 ? array_update_79747 : array_update_79736[5];
  assign array_update_79749[6] = add_78772 == 32'h0000_0006 ? array_update_79747 : array_update_79736[6];
  assign array_update_79749[7] = add_78772 == 32'h0000_0007 ? array_update_79747 : array_update_79736[7];
  assign array_update_79749[8] = add_78772 == 32'h0000_0008 ? array_update_79747 : array_update_79736[8];
  assign array_update_79749[9] = add_78772 == 32'h0000_0009 ? array_update_79747 : array_update_79736[9];
  assign array_index_79751 = array_update_72021[add_79748 > 32'h0000_0009 ? 4'h9 : add_79748[3:0]];
  assign array_index_79752 = array_update_79749[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_79756 = smul32b_32b_x_32b(array_index_78779[add_79748 > 32'h0000_0009 ? 4'h9 : add_79748[3:0]], array_index_79751[add_79720 > 32'h0000_0009 ? 4'h9 : add_79720[3:0]]);
  assign add_79758 = array_index_79752[add_79720 > 32'h0000_0009 ? 4'h9 : add_79720[3:0]] + smul_79756;
  assign array_update_79760[0] = add_79720 == 32'h0000_0000 ? add_79758 : array_index_79752[0];
  assign array_update_79760[1] = add_79720 == 32'h0000_0001 ? add_79758 : array_index_79752[1];
  assign array_update_79760[2] = add_79720 == 32'h0000_0002 ? add_79758 : array_index_79752[2];
  assign array_update_79760[3] = add_79720 == 32'h0000_0003 ? add_79758 : array_index_79752[3];
  assign array_update_79760[4] = add_79720 == 32'h0000_0004 ? add_79758 : array_index_79752[4];
  assign array_update_79760[5] = add_79720 == 32'h0000_0005 ? add_79758 : array_index_79752[5];
  assign array_update_79760[6] = add_79720 == 32'h0000_0006 ? add_79758 : array_index_79752[6];
  assign array_update_79760[7] = add_79720 == 32'h0000_0007 ? add_79758 : array_index_79752[7];
  assign array_update_79760[8] = add_79720 == 32'h0000_0008 ? add_79758 : array_index_79752[8];
  assign array_update_79760[9] = add_79720 == 32'h0000_0009 ? add_79758 : array_index_79752[9];
  assign add_79761 = add_79748 + 32'h0000_0001;
  assign array_update_79762[0] = add_78772 == 32'h0000_0000 ? array_update_79760 : array_update_79749[0];
  assign array_update_79762[1] = add_78772 == 32'h0000_0001 ? array_update_79760 : array_update_79749[1];
  assign array_update_79762[2] = add_78772 == 32'h0000_0002 ? array_update_79760 : array_update_79749[2];
  assign array_update_79762[3] = add_78772 == 32'h0000_0003 ? array_update_79760 : array_update_79749[3];
  assign array_update_79762[4] = add_78772 == 32'h0000_0004 ? array_update_79760 : array_update_79749[4];
  assign array_update_79762[5] = add_78772 == 32'h0000_0005 ? array_update_79760 : array_update_79749[5];
  assign array_update_79762[6] = add_78772 == 32'h0000_0006 ? array_update_79760 : array_update_79749[6];
  assign array_update_79762[7] = add_78772 == 32'h0000_0007 ? array_update_79760 : array_update_79749[7];
  assign array_update_79762[8] = add_78772 == 32'h0000_0008 ? array_update_79760 : array_update_79749[8];
  assign array_update_79762[9] = add_78772 == 32'h0000_0009 ? array_update_79760 : array_update_79749[9];
  assign array_index_79764 = array_update_72021[add_79761 > 32'h0000_0009 ? 4'h9 : add_79761[3:0]];
  assign array_index_79765 = array_update_79762[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_79769 = smul32b_32b_x_32b(array_index_78779[add_79761 > 32'h0000_0009 ? 4'h9 : add_79761[3:0]], array_index_79764[add_79720 > 32'h0000_0009 ? 4'h9 : add_79720[3:0]]);
  assign add_79771 = array_index_79765[add_79720 > 32'h0000_0009 ? 4'h9 : add_79720[3:0]] + smul_79769;
  assign array_update_79773[0] = add_79720 == 32'h0000_0000 ? add_79771 : array_index_79765[0];
  assign array_update_79773[1] = add_79720 == 32'h0000_0001 ? add_79771 : array_index_79765[1];
  assign array_update_79773[2] = add_79720 == 32'h0000_0002 ? add_79771 : array_index_79765[2];
  assign array_update_79773[3] = add_79720 == 32'h0000_0003 ? add_79771 : array_index_79765[3];
  assign array_update_79773[4] = add_79720 == 32'h0000_0004 ? add_79771 : array_index_79765[4];
  assign array_update_79773[5] = add_79720 == 32'h0000_0005 ? add_79771 : array_index_79765[5];
  assign array_update_79773[6] = add_79720 == 32'h0000_0006 ? add_79771 : array_index_79765[6];
  assign array_update_79773[7] = add_79720 == 32'h0000_0007 ? add_79771 : array_index_79765[7];
  assign array_update_79773[8] = add_79720 == 32'h0000_0008 ? add_79771 : array_index_79765[8];
  assign array_update_79773[9] = add_79720 == 32'h0000_0009 ? add_79771 : array_index_79765[9];
  assign add_79774 = add_79761 + 32'h0000_0001;
  assign array_update_79775[0] = add_78772 == 32'h0000_0000 ? array_update_79773 : array_update_79762[0];
  assign array_update_79775[1] = add_78772 == 32'h0000_0001 ? array_update_79773 : array_update_79762[1];
  assign array_update_79775[2] = add_78772 == 32'h0000_0002 ? array_update_79773 : array_update_79762[2];
  assign array_update_79775[3] = add_78772 == 32'h0000_0003 ? array_update_79773 : array_update_79762[3];
  assign array_update_79775[4] = add_78772 == 32'h0000_0004 ? array_update_79773 : array_update_79762[4];
  assign array_update_79775[5] = add_78772 == 32'h0000_0005 ? array_update_79773 : array_update_79762[5];
  assign array_update_79775[6] = add_78772 == 32'h0000_0006 ? array_update_79773 : array_update_79762[6];
  assign array_update_79775[7] = add_78772 == 32'h0000_0007 ? array_update_79773 : array_update_79762[7];
  assign array_update_79775[8] = add_78772 == 32'h0000_0008 ? array_update_79773 : array_update_79762[8];
  assign array_update_79775[9] = add_78772 == 32'h0000_0009 ? array_update_79773 : array_update_79762[9];
  assign array_index_79777 = array_update_72021[add_79774 > 32'h0000_0009 ? 4'h9 : add_79774[3:0]];
  assign array_index_79778 = array_update_79775[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_79782 = smul32b_32b_x_32b(array_index_78779[add_79774 > 32'h0000_0009 ? 4'h9 : add_79774[3:0]], array_index_79777[add_79720 > 32'h0000_0009 ? 4'h9 : add_79720[3:0]]);
  assign add_79784 = array_index_79778[add_79720 > 32'h0000_0009 ? 4'h9 : add_79720[3:0]] + smul_79782;
  assign array_update_79786[0] = add_79720 == 32'h0000_0000 ? add_79784 : array_index_79778[0];
  assign array_update_79786[1] = add_79720 == 32'h0000_0001 ? add_79784 : array_index_79778[1];
  assign array_update_79786[2] = add_79720 == 32'h0000_0002 ? add_79784 : array_index_79778[2];
  assign array_update_79786[3] = add_79720 == 32'h0000_0003 ? add_79784 : array_index_79778[3];
  assign array_update_79786[4] = add_79720 == 32'h0000_0004 ? add_79784 : array_index_79778[4];
  assign array_update_79786[5] = add_79720 == 32'h0000_0005 ? add_79784 : array_index_79778[5];
  assign array_update_79786[6] = add_79720 == 32'h0000_0006 ? add_79784 : array_index_79778[6];
  assign array_update_79786[7] = add_79720 == 32'h0000_0007 ? add_79784 : array_index_79778[7];
  assign array_update_79786[8] = add_79720 == 32'h0000_0008 ? add_79784 : array_index_79778[8];
  assign array_update_79786[9] = add_79720 == 32'h0000_0009 ? add_79784 : array_index_79778[9];
  assign add_79787 = add_79774 + 32'h0000_0001;
  assign array_update_79788[0] = add_78772 == 32'h0000_0000 ? array_update_79786 : array_update_79775[0];
  assign array_update_79788[1] = add_78772 == 32'h0000_0001 ? array_update_79786 : array_update_79775[1];
  assign array_update_79788[2] = add_78772 == 32'h0000_0002 ? array_update_79786 : array_update_79775[2];
  assign array_update_79788[3] = add_78772 == 32'h0000_0003 ? array_update_79786 : array_update_79775[3];
  assign array_update_79788[4] = add_78772 == 32'h0000_0004 ? array_update_79786 : array_update_79775[4];
  assign array_update_79788[5] = add_78772 == 32'h0000_0005 ? array_update_79786 : array_update_79775[5];
  assign array_update_79788[6] = add_78772 == 32'h0000_0006 ? array_update_79786 : array_update_79775[6];
  assign array_update_79788[7] = add_78772 == 32'h0000_0007 ? array_update_79786 : array_update_79775[7];
  assign array_update_79788[8] = add_78772 == 32'h0000_0008 ? array_update_79786 : array_update_79775[8];
  assign array_update_79788[9] = add_78772 == 32'h0000_0009 ? array_update_79786 : array_update_79775[9];
  assign array_index_79790 = array_update_72021[add_79787 > 32'h0000_0009 ? 4'h9 : add_79787[3:0]];
  assign array_index_79791 = array_update_79788[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_79795 = smul32b_32b_x_32b(array_index_78779[add_79787 > 32'h0000_0009 ? 4'h9 : add_79787[3:0]], array_index_79790[add_79720 > 32'h0000_0009 ? 4'h9 : add_79720[3:0]]);
  assign add_79797 = array_index_79791[add_79720 > 32'h0000_0009 ? 4'h9 : add_79720[3:0]] + smul_79795;
  assign array_update_79799[0] = add_79720 == 32'h0000_0000 ? add_79797 : array_index_79791[0];
  assign array_update_79799[1] = add_79720 == 32'h0000_0001 ? add_79797 : array_index_79791[1];
  assign array_update_79799[2] = add_79720 == 32'h0000_0002 ? add_79797 : array_index_79791[2];
  assign array_update_79799[3] = add_79720 == 32'h0000_0003 ? add_79797 : array_index_79791[3];
  assign array_update_79799[4] = add_79720 == 32'h0000_0004 ? add_79797 : array_index_79791[4];
  assign array_update_79799[5] = add_79720 == 32'h0000_0005 ? add_79797 : array_index_79791[5];
  assign array_update_79799[6] = add_79720 == 32'h0000_0006 ? add_79797 : array_index_79791[6];
  assign array_update_79799[7] = add_79720 == 32'h0000_0007 ? add_79797 : array_index_79791[7];
  assign array_update_79799[8] = add_79720 == 32'h0000_0008 ? add_79797 : array_index_79791[8];
  assign array_update_79799[9] = add_79720 == 32'h0000_0009 ? add_79797 : array_index_79791[9];
  assign add_79800 = add_79787 + 32'h0000_0001;
  assign array_update_79801[0] = add_78772 == 32'h0000_0000 ? array_update_79799 : array_update_79788[0];
  assign array_update_79801[1] = add_78772 == 32'h0000_0001 ? array_update_79799 : array_update_79788[1];
  assign array_update_79801[2] = add_78772 == 32'h0000_0002 ? array_update_79799 : array_update_79788[2];
  assign array_update_79801[3] = add_78772 == 32'h0000_0003 ? array_update_79799 : array_update_79788[3];
  assign array_update_79801[4] = add_78772 == 32'h0000_0004 ? array_update_79799 : array_update_79788[4];
  assign array_update_79801[5] = add_78772 == 32'h0000_0005 ? array_update_79799 : array_update_79788[5];
  assign array_update_79801[6] = add_78772 == 32'h0000_0006 ? array_update_79799 : array_update_79788[6];
  assign array_update_79801[7] = add_78772 == 32'h0000_0007 ? array_update_79799 : array_update_79788[7];
  assign array_update_79801[8] = add_78772 == 32'h0000_0008 ? array_update_79799 : array_update_79788[8];
  assign array_update_79801[9] = add_78772 == 32'h0000_0009 ? array_update_79799 : array_update_79788[9];
  assign array_index_79803 = array_update_72021[add_79800 > 32'h0000_0009 ? 4'h9 : add_79800[3:0]];
  assign array_index_79804 = array_update_79801[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_79808 = smul32b_32b_x_32b(array_index_78779[add_79800 > 32'h0000_0009 ? 4'h9 : add_79800[3:0]], array_index_79803[add_79720 > 32'h0000_0009 ? 4'h9 : add_79720[3:0]]);
  assign add_79810 = array_index_79804[add_79720 > 32'h0000_0009 ? 4'h9 : add_79720[3:0]] + smul_79808;
  assign array_update_79812[0] = add_79720 == 32'h0000_0000 ? add_79810 : array_index_79804[0];
  assign array_update_79812[1] = add_79720 == 32'h0000_0001 ? add_79810 : array_index_79804[1];
  assign array_update_79812[2] = add_79720 == 32'h0000_0002 ? add_79810 : array_index_79804[2];
  assign array_update_79812[3] = add_79720 == 32'h0000_0003 ? add_79810 : array_index_79804[3];
  assign array_update_79812[4] = add_79720 == 32'h0000_0004 ? add_79810 : array_index_79804[4];
  assign array_update_79812[5] = add_79720 == 32'h0000_0005 ? add_79810 : array_index_79804[5];
  assign array_update_79812[6] = add_79720 == 32'h0000_0006 ? add_79810 : array_index_79804[6];
  assign array_update_79812[7] = add_79720 == 32'h0000_0007 ? add_79810 : array_index_79804[7];
  assign array_update_79812[8] = add_79720 == 32'h0000_0008 ? add_79810 : array_index_79804[8];
  assign array_update_79812[9] = add_79720 == 32'h0000_0009 ? add_79810 : array_index_79804[9];
  assign add_79813 = add_79800 + 32'h0000_0001;
  assign array_update_79814[0] = add_78772 == 32'h0000_0000 ? array_update_79812 : array_update_79801[0];
  assign array_update_79814[1] = add_78772 == 32'h0000_0001 ? array_update_79812 : array_update_79801[1];
  assign array_update_79814[2] = add_78772 == 32'h0000_0002 ? array_update_79812 : array_update_79801[2];
  assign array_update_79814[3] = add_78772 == 32'h0000_0003 ? array_update_79812 : array_update_79801[3];
  assign array_update_79814[4] = add_78772 == 32'h0000_0004 ? array_update_79812 : array_update_79801[4];
  assign array_update_79814[5] = add_78772 == 32'h0000_0005 ? array_update_79812 : array_update_79801[5];
  assign array_update_79814[6] = add_78772 == 32'h0000_0006 ? array_update_79812 : array_update_79801[6];
  assign array_update_79814[7] = add_78772 == 32'h0000_0007 ? array_update_79812 : array_update_79801[7];
  assign array_update_79814[8] = add_78772 == 32'h0000_0008 ? array_update_79812 : array_update_79801[8];
  assign array_update_79814[9] = add_78772 == 32'h0000_0009 ? array_update_79812 : array_update_79801[9];
  assign array_index_79816 = array_update_72021[add_79813 > 32'h0000_0009 ? 4'h9 : add_79813[3:0]];
  assign array_index_79817 = array_update_79814[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_79821 = smul32b_32b_x_32b(array_index_78779[add_79813 > 32'h0000_0009 ? 4'h9 : add_79813[3:0]], array_index_79816[add_79720 > 32'h0000_0009 ? 4'h9 : add_79720[3:0]]);
  assign add_79823 = array_index_79817[add_79720 > 32'h0000_0009 ? 4'h9 : add_79720[3:0]] + smul_79821;
  assign array_update_79825[0] = add_79720 == 32'h0000_0000 ? add_79823 : array_index_79817[0];
  assign array_update_79825[1] = add_79720 == 32'h0000_0001 ? add_79823 : array_index_79817[1];
  assign array_update_79825[2] = add_79720 == 32'h0000_0002 ? add_79823 : array_index_79817[2];
  assign array_update_79825[3] = add_79720 == 32'h0000_0003 ? add_79823 : array_index_79817[3];
  assign array_update_79825[4] = add_79720 == 32'h0000_0004 ? add_79823 : array_index_79817[4];
  assign array_update_79825[5] = add_79720 == 32'h0000_0005 ? add_79823 : array_index_79817[5];
  assign array_update_79825[6] = add_79720 == 32'h0000_0006 ? add_79823 : array_index_79817[6];
  assign array_update_79825[7] = add_79720 == 32'h0000_0007 ? add_79823 : array_index_79817[7];
  assign array_update_79825[8] = add_79720 == 32'h0000_0008 ? add_79823 : array_index_79817[8];
  assign array_update_79825[9] = add_79720 == 32'h0000_0009 ? add_79823 : array_index_79817[9];
  assign add_79826 = add_79813 + 32'h0000_0001;
  assign array_update_79827[0] = add_78772 == 32'h0000_0000 ? array_update_79825 : array_update_79814[0];
  assign array_update_79827[1] = add_78772 == 32'h0000_0001 ? array_update_79825 : array_update_79814[1];
  assign array_update_79827[2] = add_78772 == 32'h0000_0002 ? array_update_79825 : array_update_79814[2];
  assign array_update_79827[3] = add_78772 == 32'h0000_0003 ? array_update_79825 : array_update_79814[3];
  assign array_update_79827[4] = add_78772 == 32'h0000_0004 ? array_update_79825 : array_update_79814[4];
  assign array_update_79827[5] = add_78772 == 32'h0000_0005 ? array_update_79825 : array_update_79814[5];
  assign array_update_79827[6] = add_78772 == 32'h0000_0006 ? array_update_79825 : array_update_79814[6];
  assign array_update_79827[7] = add_78772 == 32'h0000_0007 ? array_update_79825 : array_update_79814[7];
  assign array_update_79827[8] = add_78772 == 32'h0000_0008 ? array_update_79825 : array_update_79814[8];
  assign array_update_79827[9] = add_78772 == 32'h0000_0009 ? array_update_79825 : array_update_79814[9];
  assign array_index_79829 = array_update_72021[add_79826 > 32'h0000_0009 ? 4'h9 : add_79826[3:0]];
  assign array_index_79830 = array_update_79827[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_79834 = smul32b_32b_x_32b(array_index_78779[add_79826 > 32'h0000_0009 ? 4'h9 : add_79826[3:0]], array_index_79829[add_79720 > 32'h0000_0009 ? 4'h9 : add_79720[3:0]]);
  assign add_79836 = array_index_79830[add_79720 > 32'h0000_0009 ? 4'h9 : add_79720[3:0]] + smul_79834;
  assign array_update_79838[0] = add_79720 == 32'h0000_0000 ? add_79836 : array_index_79830[0];
  assign array_update_79838[1] = add_79720 == 32'h0000_0001 ? add_79836 : array_index_79830[1];
  assign array_update_79838[2] = add_79720 == 32'h0000_0002 ? add_79836 : array_index_79830[2];
  assign array_update_79838[3] = add_79720 == 32'h0000_0003 ? add_79836 : array_index_79830[3];
  assign array_update_79838[4] = add_79720 == 32'h0000_0004 ? add_79836 : array_index_79830[4];
  assign array_update_79838[5] = add_79720 == 32'h0000_0005 ? add_79836 : array_index_79830[5];
  assign array_update_79838[6] = add_79720 == 32'h0000_0006 ? add_79836 : array_index_79830[6];
  assign array_update_79838[7] = add_79720 == 32'h0000_0007 ? add_79836 : array_index_79830[7];
  assign array_update_79838[8] = add_79720 == 32'h0000_0008 ? add_79836 : array_index_79830[8];
  assign array_update_79838[9] = add_79720 == 32'h0000_0009 ? add_79836 : array_index_79830[9];
  assign add_79839 = add_79826 + 32'h0000_0001;
  assign array_update_79840[0] = add_78772 == 32'h0000_0000 ? array_update_79838 : array_update_79827[0];
  assign array_update_79840[1] = add_78772 == 32'h0000_0001 ? array_update_79838 : array_update_79827[1];
  assign array_update_79840[2] = add_78772 == 32'h0000_0002 ? array_update_79838 : array_update_79827[2];
  assign array_update_79840[3] = add_78772 == 32'h0000_0003 ? array_update_79838 : array_update_79827[3];
  assign array_update_79840[4] = add_78772 == 32'h0000_0004 ? array_update_79838 : array_update_79827[4];
  assign array_update_79840[5] = add_78772 == 32'h0000_0005 ? array_update_79838 : array_update_79827[5];
  assign array_update_79840[6] = add_78772 == 32'h0000_0006 ? array_update_79838 : array_update_79827[6];
  assign array_update_79840[7] = add_78772 == 32'h0000_0007 ? array_update_79838 : array_update_79827[7];
  assign array_update_79840[8] = add_78772 == 32'h0000_0008 ? array_update_79838 : array_update_79827[8];
  assign array_update_79840[9] = add_78772 == 32'h0000_0009 ? array_update_79838 : array_update_79827[9];
  assign array_index_79842 = array_update_72021[add_79839 > 32'h0000_0009 ? 4'h9 : add_79839[3:0]];
  assign array_index_79843 = array_update_79840[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_79847 = smul32b_32b_x_32b(array_index_78779[add_79839 > 32'h0000_0009 ? 4'h9 : add_79839[3:0]], array_index_79842[add_79720 > 32'h0000_0009 ? 4'h9 : add_79720[3:0]]);
  assign add_79849 = array_index_79843[add_79720 > 32'h0000_0009 ? 4'h9 : add_79720[3:0]] + smul_79847;
  assign array_update_79850[0] = add_79720 == 32'h0000_0000 ? add_79849 : array_index_79843[0];
  assign array_update_79850[1] = add_79720 == 32'h0000_0001 ? add_79849 : array_index_79843[1];
  assign array_update_79850[2] = add_79720 == 32'h0000_0002 ? add_79849 : array_index_79843[2];
  assign array_update_79850[3] = add_79720 == 32'h0000_0003 ? add_79849 : array_index_79843[3];
  assign array_update_79850[4] = add_79720 == 32'h0000_0004 ? add_79849 : array_index_79843[4];
  assign array_update_79850[5] = add_79720 == 32'h0000_0005 ? add_79849 : array_index_79843[5];
  assign array_update_79850[6] = add_79720 == 32'h0000_0006 ? add_79849 : array_index_79843[6];
  assign array_update_79850[7] = add_79720 == 32'h0000_0007 ? add_79849 : array_index_79843[7];
  assign array_update_79850[8] = add_79720 == 32'h0000_0008 ? add_79849 : array_index_79843[8];
  assign array_update_79850[9] = add_79720 == 32'h0000_0009 ? add_79849 : array_index_79843[9];
  assign array_update_79851[0] = add_78772 == 32'h0000_0000 ? array_update_79850 : array_update_79840[0];
  assign array_update_79851[1] = add_78772 == 32'h0000_0001 ? array_update_79850 : array_update_79840[1];
  assign array_update_79851[2] = add_78772 == 32'h0000_0002 ? array_update_79850 : array_update_79840[2];
  assign array_update_79851[3] = add_78772 == 32'h0000_0003 ? array_update_79850 : array_update_79840[3];
  assign array_update_79851[4] = add_78772 == 32'h0000_0004 ? array_update_79850 : array_update_79840[4];
  assign array_update_79851[5] = add_78772 == 32'h0000_0005 ? array_update_79850 : array_update_79840[5];
  assign array_update_79851[6] = add_78772 == 32'h0000_0006 ? array_update_79850 : array_update_79840[6];
  assign array_update_79851[7] = add_78772 == 32'h0000_0007 ? array_update_79850 : array_update_79840[7];
  assign array_update_79851[8] = add_78772 == 32'h0000_0008 ? array_update_79850 : array_update_79840[8];
  assign array_update_79851[9] = add_78772 == 32'h0000_0009 ? array_update_79850 : array_update_79840[9];
  assign array_index_79853 = array_update_79851[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign add_79855 = add_79720 + 32'h0000_0001;
  assign array_update_79856[0] = add_79855 == 32'h0000_0000 ? 32'h0000_0000 : array_index_79853[0];
  assign array_update_79856[1] = add_79855 == 32'h0000_0001 ? 32'h0000_0000 : array_index_79853[1];
  assign array_update_79856[2] = add_79855 == 32'h0000_0002 ? 32'h0000_0000 : array_index_79853[2];
  assign array_update_79856[3] = add_79855 == 32'h0000_0003 ? 32'h0000_0000 : array_index_79853[3];
  assign array_update_79856[4] = add_79855 == 32'h0000_0004 ? 32'h0000_0000 : array_index_79853[4];
  assign array_update_79856[5] = add_79855 == 32'h0000_0005 ? 32'h0000_0000 : array_index_79853[5];
  assign array_update_79856[6] = add_79855 == 32'h0000_0006 ? 32'h0000_0000 : array_index_79853[6];
  assign array_update_79856[7] = add_79855 == 32'h0000_0007 ? 32'h0000_0000 : array_index_79853[7];
  assign array_update_79856[8] = add_79855 == 32'h0000_0008 ? 32'h0000_0000 : array_index_79853[8];
  assign array_update_79856[9] = add_79855 == 32'h0000_0009 ? 32'h0000_0000 : array_index_79853[9];
  assign literal_79857 = 32'h0000_0000;
  assign array_update_79858[0] = add_78772 == 32'h0000_0000 ? array_update_79856 : array_update_79851[0];
  assign array_update_79858[1] = add_78772 == 32'h0000_0001 ? array_update_79856 : array_update_79851[1];
  assign array_update_79858[2] = add_78772 == 32'h0000_0002 ? array_update_79856 : array_update_79851[2];
  assign array_update_79858[3] = add_78772 == 32'h0000_0003 ? array_update_79856 : array_update_79851[3];
  assign array_update_79858[4] = add_78772 == 32'h0000_0004 ? array_update_79856 : array_update_79851[4];
  assign array_update_79858[5] = add_78772 == 32'h0000_0005 ? array_update_79856 : array_update_79851[5];
  assign array_update_79858[6] = add_78772 == 32'h0000_0006 ? array_update_79856 : array_update_79851[6];
  assign array_update_79858[7] = add_78772 == 32'h0000_0007 ? array_update_79856 : array_update_79851[7];
  assign array_update_79858[8] = add_78772 == 32'h0000_0008 ? array_update_79856 : array_update_79851[8];
  assign array_update_79858[9] = add_78772 == 32'h0000_0009 ? array_update_79856 : array_update_79851[9];
  assign array_index_79860 = array_update_72021[literal_79857 > 32'h0000_0009 ? 4'h9 : literal_79857[3:0]];
  assign array_index_79861 = array_update_79858[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_79865 = smul32b_32b_x_32b(array_index_78779[literal_79857 > 32'h0000_0009 ? 4'h9 : literal_79857[3:0]], array_index_79860[add_79855 > 32'h0000_0009 ? 4'h9 : add_79855[3:0]]);
  assign add_79867 = array_index_79861[add_79855 > 32'h0000_0009 ? 4'h9 : add_79855[3:0]] + smul_79865;
  assign array_update_79869[0] = add_79855 == 32'h0000_0000 ? add_79867 : array_index_79861[0];
  assign array_update_79869[1] = add_79855 == 32'h0000_0001 ? add_79867 : array_index_79861[1];
  assign array_update_79869[2] = add_79855 == 32'h0000_0002 ? add_79867 : array_index_79861[2];
  assign array_update_79869[3] = add_79855 == 32'h0000_0003 ? add_79867 : array_index_79861[3];
  assign array_update_79869[4] = add_79855 == 32'h0000_0004 ? add_79867 : array_index_79861[4];
  assign array_update_79869[5] = add_79855 == 32'h0000_0005 ? add_79867 : array_index_79861[5];
  assign array_update_79869[6] = add_79855 == 32'h0000_0006 ? add_79867 : array_index_79861[6];
  assign array_update_79869[7] = add_79855 == 32'h0000_0007 ? add_79867 : array_index_79861[7];
  assign array_update_79869[8] = add_79855 == 32'h0000_0008 ? add_79867 : array_index_79861[8];
  assign array_update_79869[9] = add_79855 == 32'h0000_0009 ? add_79867 : array_index_79861[9];
  assign add_79870 = literal_79857 + 32'h0000_0001;
  assign array_update_79871[0] = add_78772 == 32'h0000_0000 ? array_update_79869 : array_update_79858[0];
  assign array_update_79871[1] = add_78772 == 32'h0000_0001 ? array_update_79869 : array_update_79858[1];
  assign array_update_79871[2] = add_78772 == 32'h0000_0002 ? array_update_79869 : array_update_79858[2];
  assign array_update_79871[3] = add_78772 == 32'h0000_0003 ? array_update_79869 : array_update_79858[3];
  assign array_update_79871[4] = add_78772 == 32'h0000_0004 ? array_update_79869 : array_update_79858[4];
  assign array_update_79871[5] = add_78772 == 32'h0000_0005 ? array_update_79869 : array_update_79858[5];
  assign array_update_79871[6] = add_78772 == 32'h0000_0006 ? array_update_79869 : array_update_79858[6];
  assign array_update_79871[7] = add_78772 == 32'h0000_0007 ? array_update_79869 : array_update_79858[7];
  assign array_update_79871[8] = add_78772 == 32'h0000_0008 ? array_update_79869 : array_update_79858[8];
  assign array_update_79871[9] = add_78772 == 32'h0000_0009 ? array_update_79869 : array_update_79858[9];
  assign array_index_79873 = array_update_72021[add_79870 > 32'h0000_0009 ? 4'h9 : add_79870[3:0]];
  assign array_index_79874 = array_update_79871[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_79878 = smul32b_32b_x_32b(array_index_78779[add_79870 > 32'h0000_0009 ? 4'h9 : add_79870[3:0]], array_index_79873[add_79855 > 32'h0000_0009 ? 4'h9 : add_79855[3:0]]);
  assign add_79880 = array_index_79874[add_79855 > 32'h0000_0009 ? 4'h9 : add_79855[3:0]] + smul_79878;
  assign array_update_79882[0] = add_79855 == 32'h0000_0000 ? add_79880 : array_index_79874[0];
  assign array_update_79882[1] = add_79855 == 32'h0000_0001 ? add_79880 : array_index_79874[1];
  assign array_update_79882[2] = add_79855 == 32'h0000_0002 ? add_79880 : array_index_79874[2];
  assign array_update_79882[3] = add_79855 == 32'h0000_0003 ? add_79880 : array_index_79874[3];
  assign array_update_79882[4] = add_79855 == 32'h0000_0004 ? add_79880 : array_index_79874[4];
  assign array_update_79882[5] = add_79855 == 32'h0000_0005 ? add_79880 : array_index_79874[5];
  assign array_update_79882[6] = add_79855 == 32'h0000_0006 ? add_79880 : array_index_79874[6];
  assign array_update_79882[7] = add_79855 == 32'h0000_0007 ? add_79880 : array_index_79874[7];
  assign array_update_79882[8] = add_79855 == 32'h0000_0008 ? add_79880 : array_index_79874[8];
  assign array_update_79882[9] = add_79855 == 32'h0000_0009 ? add_79880 : array_index_79874[9];
  assign add_79883 = add_79870 + 32'h0000_0001;
  assign array_update_79884[0] = add_78772 == 32'h0000_0000 ? array_update_79882 : array_update_79871[0];
  assign array_update_79884[1] = add_78772 == 32'h0000_0001 ? array_update_79882 : array_update_79871[1];
  assign array_update_79884[2] = add_78772 == 32'h0000_0002 ? array_update_79882 : array_update_79871[2];
  assign array_update_79884[3] = add_78772 == 32'h0000_0003 ? array_update_79882 : array_update_79871[3];
  assign array_update_79884[4] = add_78772 == 32'h0000_0004 ? array_update_79882 : array_update_79871[4];
  assign array_update_79884[5] = add_78772 == 32'h0000_0005 ? array_update_79882 : array_update_79871[5];
  assign array_update_79884[6] = add_78772 == 32'h0000_0006 ? array_update_79882 : array_update_79871[6];
  assign array_update_79884[7] = add_78772 == 32'h0000_0007 ? array_update_79882 : array_update_79871[7];
  assign array_update_79884[8] = add_78772 == 32'h0000_0008 ? array_update_79882 : array_update_79871[8];
  assign array_update_79884[9] = add_78772 == 32'h0000_0009 ? array_update_79882 : array_update_79871[9];
  assign array_index_79886 = array_update_72021[add_79883 > 32'h0000_0009 ? 4'h9 : add_79883[3:0]];
  assign array_index_79887 = array_update_79884[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_79891 = smul32b_32b_x_32b(array_index_78779[add_79883 > 32'h0000_0009 ? 4'h9 : add_79883[3:0]], array_index_79886[add_79855 > 32'h0000_0009 ? 4'h9 : add_79855[3:0]]);
  assign add_79893 = array_index_79887[add_79855 > 32'h0000_0009 ? 4'h9 : add_79855[3:0]] + smul_79891;
  assign array_update_79895[0] = add_79855 == 32'h0000_0000 ? add_79893 : array_index_79887[0];
  assign array_update_79895[1] = add_79855 == 32'h0000_0001 ? add_79893 : array_index_79887[1];
  assign array_update_79895[2] = add_79855 == 32'h0000_0002 ? add_79893 : array_index_79887[2];
  assign array_update_79895[3] = add_79855 == 32'h0000_0003 ? add_79893 : array_index_79887[3];
  assign array_update_79895[4] = add_79855 == 32'h0000_0004 ? add_79893 : array_index_79887[4];
  assign array_update_79895[5] = add_79855 == 32'h0000_0005 ? add_79893 : array_index_79887[5];
  assign array_update_79895[6] = add_79855 == 32'h0000_0006 ? add_79893 : array_index_79887[6];
  assign array_update_79895[7] = add_79855 == 32'h0000_0007 ? add_79893 : array_index_79887[7];
  assign array_update_79895[8] = add_79855 == 32'h0000_0008 ? add_79893 : array_index_79887[8];
  assign array_update_79895[9] = add_79855 == 32'h0000_0009 ? add_79893 : array_index_79887[9];
  assign add_79896 = add_79883 + 32'h0000_0001;
  assign array_update_79897[0] = add_78772 == 32'h0000_0000 ? array_update_79895 : array_update_79884[0];
  assign array_update_79897[1] = add_78772 == 32'h0000_0001 ? array_update_79895 : array_update_79884[1];
  assign array_update_79897[2] = add_78772 == 32'h0000_0002 ? array_update_79895 : array_update_79884[2];
  assign array_update_79897[3] = add_78772 == 32'h0000_0003 ? array_update_79895 : array_update_79884[3];
  assign array_update_79897[4] = add_78772 == 32'h0000_0004 ? array_update_79895 : array_update_79884[4];
  assign array_update_79897[5] = add_78772 == 32'h0000_0005 ? array_update_79895 : array_update_79884[5];
  assign array_update_79897[6] = add_78772 == 32'h0000_0006 ? array_update_79895 : array_update_79884[6];
  assign array_update_79897[7] = add_78772 == 32'h0000_0007 ? array_update_79895 : array_update_79884[7];
  assign array_update_79897[8] = add_78772 == 32'h0000_0008 ? array_update_79895 : array_update_79884[8];
  assign array_update_79897[9] = add_78772 == 32'h0000_0009 ? array_update_79895 : array_update_79884[9];
  assign array_index_79899 = array_update_72021[add_79896 > 32'h0000_0009 ? 4'h9 : add_79896[3:0]];
  assign array_index_79900 = array_update_79897[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_79904 = smul32b_32b_x_32b(array_index_78779[add_79896 > 32'h0000_0009 ? 4'h9 : add_79896[3:0]], array_index_79899[add_79855 > 32'h0000_0009 ? 4'h9 : add_79855[3:0]]);
  assign add_79906 = array_index_79900[add_79855 > 32'h0000_0009 ? 4'h9 : add_79855[3:0]] + smul_79904;
  assign array_update_79908[0] = add_79855 == 32'h0000_0000 ? add_79906 : array_index_79900[0];
  assign array_update_79908[1] = add_79855 == 32'h0000_0001 ? add_79906 : array_index_79900[1];
  assign array_update_79908[2] = add_79855 == 32'h0000_0002 ? add_79906 : array_index_79900[2];
  assign array_update_79908[3] = add_79855 == 32'h0000_0003 ? add_79906 : array_index_79900[3];
  assign array_update_79908[4] = add_79855 == 32'h0000_0004 ? add_79906 : array_index_79900[4];
  assign array_update_79908[5] = add_79855 == 32'h0000_0005 ? add_79906 : array_index_79900[5];
  assign array_update_79908[6] = add_79855 == 32'h0000_0006 ? add_79906 : array_index_79900[6];
  assign array_update_79908[7] = add_79855 == 32'h0000_0007 ? add_79906 : array_index_79900[7];
  assign array_update_79908[8] = add_79855 == 32'h0000_0008 ? add_79906 : array_index_79900[8];
  assign array_update_79908[9] = add_79855 == 32'h0000_0009 ? add_79906 : array_index_79900[9];
  assign add_79909 = add_79896 + 32'h0000_0001;
  assign array_update_79910[0] = add_78772 == 32'h0000_0000 ? array_update_79908 : array_update_79897[0];
  assign array_update_79910[1] = add_78772 == 32'h0000_0001 ? array_update_79908 : array_update_79897[1];
  assign array_update_79910[2] = add_78772 == 32'h0000_0002 ? array_update_79908 : array_update_79897[2];
  assign array_update_79910[3] = add_78772 == 32'h0000_0003 ? array_update_79908 : array_update_79897[3];
  assign array_update_79910[4] = add_78772 == 32'h0000_0004 ? array_update_79908 : array_update_79897[4];
  assign array_update_79910[5] = add_78772 == 32'h0000_0005 ? array_update_79908 : array_update_79897[5];
  assign array_update_79910[6] = add_78772 == 32'h0000_0006 ? array_update_79908 : array_update_79897[6];
  assign array_update_79910[7] = add_78772 == 32'h0000_0007 ? array_update_79908 : array_update_79897[7];
  assign array_update_79910[8] = add_78772 == 32'h0000_0008 ? array_update_79908 : array_update_79897[8];
  assign array_update_79910[9] = add_78772 == 32'h0000_0009 ? array_update_79908 : array_update_79897[9];
  assign array_index_79912 = array_update_72021[add_79909 > 32'h0000_0009 ? 4'h9 : add_79909[3:0]];
  assign array_index_79913 = array_update_79910[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_79917 = smul32b_32b_x_32b(array_index_78779[add_79909 > 32'h0000_0009 ? 4'h9 : add_79909[3:0]], array_index_79912[add_79855 > 32'h0000_0009 ? 4'h9 : add_79855[3:0]]);
  assign add_79919 = array_index_79913[add_79855 > 32'h0000_0009 ? 4'h9 : add_79855[3:0]] + smul_79917;
  assign array_update_79921[0] = add_79855 == 32'h0000_0000 ? add_79919 : array_index_79913[0];
  assign array_update_79921[1] = add_79855 == 32'h0000_0001 ? add_79919 : array_index_79913[1];
  assign array_update_79921[2] = add_79855 == 32'h0000_0002 ? add_79919 : array_index_79913[2];
  assign array_update_79921[3] = add_79855 == 32'h0000_0003 ? add_79919 : array_index_79913[3];
  assign array_update_79921[4] = add_79855 == 32'h0000_0004 ? add_79919 : array_index_79913[4];
  assign array_update_79921[5] = add_79855 == 32'h0000_0005 ? add_79919 : array_index_79913[5];
  assign array_update_79921[6] = add_79855 == 32'h0000_0006 ? add_79919 : array_index_79913[6];
  assign array_update_79921[7] = add_79855 == 32'h0000_0007 ? add_79919 : array_index_79913[7];
  assign array_update_79921[8] = add_79855 == 32'h0000_0008 ? add_79919 : array_index_79913[8];
  assign array_update_79921[9] = add_79855 == 32'h0000_0009 ? add_79919 : array_index_79913[9];
  assign add_79922 = add_79909 + 32'h0000_0001;
  assign array_update_79923[0] = add_78772 == 32'h0000_0000 ? array_update_79921 : array_update_79910[0];
  assign array_update_79923[1] = add_78772 == 32'h0000_0001 ? array_update_79921 : array_update_79910[1];
  assign array_update_79923[2] = add_78772 == 32'h0000_0002 ? array_update_79921 : array_update_79910[2];
  assign array_update_79923[3] = add_78772 == 32'h0000_0003 ? array_update_79921 : array_update_79910[3];
  assign array_update_79923[4] = add_78772 == 32'h0000_0004 ? array_update_79921 : array_update_79910[4];
  assign array_update_79923[5] = add_78772 == 32'h0000_0005 ? array_update_79921 : array_update_79910[5];
  assign array_update_79923[6] = add_78772 == 32'h0000_0006 ? array_update_79921 : array_update_79910[6];
  assign array_update_79923[7] = add_78772 == 32'h0000_0007 ? array_update_79921 : array_update_79910[7];
  assign array_update_79923[8] = add_78772 == 32'h0000_0008 ? array_update_79921 : array_update_79910[8];
  assign array_update_79923[9] = add_78772 == 32'h0000_0009 ? array_update_79921 : array_update_79910[9];
  assign array_index_79925 = array_update_72021[add_79922 > 32'h0000_0009 ? 4'h9 : add_79922[3:0]];
  assign array_index_79926 = array_update_79923[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_79930 = smul32b_32b_x_32b(array_index_78779[add_79922 > 32'h0000_0009 ? 4'h9 : add_79922[3:0]], array_index_79925[add_79855 > 32'h0000_0009 ? 4'h9 : add_79855[3:0]]);
  assign add_79932 = array_index_79926[add_79855 > 32'h0000_0009 ? 4'h9 : add_79855[3:0]] + smul_79930;
  assign array_update_79934[0] = add_79855 == 32'h0000_0000 ? add_79932 : array_index_79926[0];
  assign array_update_79934[1] = add_79855 == 32'h0000_0001 ? add_79932 : array_index_79926[1];
  assign array_update_79934[2] = add_79855 == 32'h0000_0002 ? add_79932 : array_index_79926[2];
  assign array_update_79934[3] = add_79855 == 32'h0000_0003 ? add_79932 : array_index_79926[3];
  assign array_update_79934[4] = add_79855 == 32'h0000_0004 ? add_79932 : array_index_79926[4];
  assign array_update_79934[5] = add_79855 == 32'h0000_0005 ? add_79932 : array_index_79926[5];
  assign array_update_79934[6] = add_79855 == 32'h0000_0006 ? add_79932 : array_index_79926[6];
  assign array_update_79934[7] = add_79855 == 32'h0000_0007 ? add_79932 : array_index_79926[7];
  assign array_update_79934[8] = add_79855 == 32'h0000_0008 ? add_79932 : array_index_79926[8];
  assign array_update_79934[9] = add_79855 == 32'h0000_0009 ? add_79932 : array_index_79926[9];
  assign add_79935 = add_79922 + 32'h0000_0001;
  assign array_update_79936[0] = add_78772 == 32'h0000_0000 ? array_update_79934 : array_update_79923[0];
  assign array_update_79936[1] = add_78772 == 32'h0000_0001 ? array_update_79934 : array_update_79923[1];
  assign array_update_79936[2] = add_78772 == 32'h0000_0002 ? array_update_79934 : array_update_79923[2];
  assign array_update_79936[3] = add_78772 == 32'h0000_0003 ? array_update_79934 : array_update_79923[3];
  assign array_update_79936[4] = add_78772 == 32'h0000_0004 ? array_update_79934 : array_update_79923[4];
  assign array_update_79936[5] = add_78772 == 32'h0000_0005 ? array_update_79934 : array_update_79923[5];
  assign array_update_79936[6] = add_78772 == 32'h0000_0006 ? array_update_79934 : array_update_79923[6];
  assign array_update_79936[7] = add_78772 == 32'h0000_0007 ? array_update_79934 : array_update_79923[7];
  assign array_update_79936[8] = add_78772 == 32'h0000_0008 ? array_update_79934 : array_update_79923[8];
  assign array_update_79936[9] = add_78772 == 32'h0000_0009 ? array_update_79934 : array_update_79923[9];
  assign array_index_79938 = array_update_72021[add_79935 > 32'h0000_0009 ? 4'h9 : add_79935[3:0]];
  assign array_index_79939 = array_update_79936[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_79943 = smul32b_32b_x_32b(array_index_78779[add_79935 > 32'h0000_0009 ? 4'h9 : add_79935[3:0]], array_index_79938[add_79855 > 32'h0000_0009 ? 4'h9 : add_79855[3:0]]);
  assign add_79945 = array_index_79939[add_79855 > 32'h0000_0009 ? 4'h9 : add_79855[3:0]] + smul_79943;
  assign array_update_79947[0] = add_79855 == 32'h0000_0000 ? add_79945 : array_index_79939[0];
  assign array_update_79947[1] = add_79855 == 32'h0000_0001 ? add_79945 : array_index_79939[1];
  assign array_update_79947[2] = add_79855 == 32'h0000_0002 ? add_79945 : array_index_79939[2];
  assign array_update_79947[3] = add_79855 == 32'h0000_0003 ? add_79945 : array_index_79939[3];
  assign array_update_79947[4] = add_79855 == 32'h0000_0004 ? add_79945 : array_index_79939[4];
  assign array_update_79947[5] = add_79855 == 32'h0000_0005 ? add_79945 : array_index_79939[5];
  assign array_update_79947[6] = add_79855 == 32'h0000_0006 ? add_79945 : array_index_79939[6];
  assign array_update_79947[7] = add_79855 == 32'h0000_0007 ? add_79945 : array_index_79939[7];
  assign array_update_79947[8] = add_79855 == 32'h0000_0008 ? add_79945 : array_index_79939[8];
  assign array_update_79947[9] = add_79855 == 32'h0000_0009 ? add_79945 : array_index_79939[9];
  assign add_79948 = add_79935 + 32'h0000_0001;
  assign array_update_79949[0] = add_78772 == 32'h0000_0000 ? array_update_79947 : array_update_79936[0];
  assign array_update_79949[1] = add_78772 == 32'h0000_0001 ? array_update_79947 : array_update_79936[1];
  assign array_update_79949[2] = add_78772 == 32'h0000_0002 ? array_update_79947 : array_update_79936[2];
  assign array_update_79949[3] = add_78772 == 32'h0000_0003 ? array_update_79947 : array_update_79936[3];
  assign array_update_79949[4] = add_78772 == 32'h0000_0004 ? array_update_79947 : array_update_79936[4];
  assign array_update_79949[5] = add_78772 == 32'h0000_0005 ? array_update_79947 : array_update_79936[5];
  assign array_update_79949[6] = add_78772 == 32'h0000_0006 ? array_update_79947 : array_update_79936[6];
  assign array_update_79949[7] = add_78772 == 32'h0000_0007 ? array_update_79947 : array_update_79936[7];
  assign array_update_79949[8] = add_78772 == 32'h0000_0008 ? array_update_79947 : array_update_79936[8];
  assign array_update_79949[9] = add_78772 == 32'h0000_0009 ? array_update_79947 : array_update_79936[9];
  assign array_index_79951 = array_update_72021[add_79948 > 32'h0000_0009 ? 4'h9 : add_79948[3:0]];
  assign array_index_79952 = array_update_79949[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_79956 = smul32b_32b_x_32b(array_index_78779[add_79948 > 32'h0000_0009 ? 4'h9 : add_79948[3:0]], array_index_79951[add_79855 > 32'h0000_0009 ? 4'h9 : add_79855[3:0]]);
  assign add_79958 = array_index_79952[add_79855 > 32'h0000_0009 ? 4'h9 : add_79855[3:0]] + smul_79956;
  assign array_update_79960[0] = add_79855 == 32'h0000_0000 ? add_79958 : array_index_79952[0];
  assign array_update_79960[1] = add_79855 == 32'h0000_0001 ? add_79958 : array_index_79952[1];
  assign array_update_79960[2] = add_79855 == 32'h0000_0002 ? add_79958 : array_index_79952[2];
  assign array_update_79960[3] = add_79855 == 32'h0000_0003 ? add_79958 : array_index_79952[3];
  assign array_update_79960[4] = add_79855 == 32'h0000_0004 ? add_79958 : array_index_79952[4];
  assign array_update_79960[5] = add_79855 == 32'h0000_0005 ? add_79958 : array_index_79952[5];
  assign array_update_79960[6] = add_79855 == 32'h0000_0006 ? add_79958 : array_index_79952[6];
  assign array_update_79960[7] = add_79855 == 32'h0000_0007 ? add_79958 : array_index_79952[7];
  assign array_update_79960[8] = add_79855 == 32'h0000_0008 ? add_79958 : array_index_79952[8];
  assign array_update_79960[9] = add_79855 == 32'h0000_0009 ? add_79958 : array_index_79952[9];
  assign add_79961 = add_79948 + 32'h0000_0001;
  assign array_update_79962[0] = add_78772 == 32'h0000_0000 ? array_update_79960 : array_update_79949[0];
  assign array_update_79962[1] = add_78772 == 32'h0000_0001 ? array_update_79960 : array_update_79949[1];
  assign array_update_79962[2] = add_78772 == 32'h0000_0002 ? array_update_79960 : array_update_79949[2];
  assign array_update_79962[3] = add_78772 == 32'h0000_0003 ? array_update_79960 : array_update_79949[3];
  assign array_update_79962[4] = add_78772 == 32'h0000_0004 ? array_update_79960 : array_update_79949[4];
  assign array_update_79962[5] = add_78772 == 32'h0000_0005 ? array_update_79960 : array_update_79949[5];
  assign array_update_79962[6] = add_78772 == 32'h0000_0006 ? array_update_79960 : array_update_79949[6];
  assign array_update_79962[7] = add_78772 == 32'h0000_0007 ? array_update_79960 : array_update_79949[7];
  assign array_update_79962[8] = add_78772 == 32'h0000_0008 ? array_update_79960 : array_update_79949[8];
  assign array_update_79962[9] = add_78772 == 32'h0000_0009 ? array_update_79960 : array_update_79949[9];
  assign array_index_79964 = array_update_72021[add_79961 > 32'h0000_0009 ? 4'h9 : add_79961[3:0]];
  assign array_index_79965 = array_update_79962[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_79969 = smul32b_32b_x_32b(array_index_78779[add_79961 > 32'h0000_0009 ? 4'h9 : add_79961[3:0]], array_index_79964[add_79855 > 32'h0000_0009 ? 4'h9 : add_79855[3:0]]);
  assign add_79971 = array_index_79965[add_79855 > 32'h0000_0009 ? 4'h9 : add_79855[3:0]] + smul_79969;
  assign array_update_79973[0] = add_79855 == 32'h0000_0000 ? add_79971 : array_index_79965[0];
  assign array_update_79973[1] = add_79855 == 32'h0000_0001 ? add_79971 : array_index_79965[1];
  assign array_update_79973[2] = add_79855 == 32'h0000_0002 ? add_79971 : array_index_79965[2];
  assign array_update_79973[3] = add_79855 == 32'h0000_0003 ? add_79971 : array_index_79965[3];
  assign array_update_79973[4] = add_79855 == 32'h0000_0004 ? add_79971 : array_index_79965[4];
  assign array_update_79973[5] = add_79855 == 32'h0000_0005 ? add_79971 : array_index_79965[5];
  assign array_update_79973[6] = add_79855 == 32'h0000_0006 ? add_79971 : array_index_79965[6];
  assign array_update_79973[7] = add_79855 == 32'h0000_0007 ? add_79971 : array_index_79965[7];
  assign array_update_79973[8] = add_79855 == 32'h0000_0008 ? add_79971 : array_index_79965[8];
  assign array_update_79973[9] = add_79855 == 32'h0000_0009 ? add_79971 : array_index_79965[9];
  assign add_79974 = add_79961 + 32'h0000_0001;
  assign array_update_79975[0] = add_78772 == 32'h0000_0000 ? array_update_79973 : array_update_79962[0];
  assign array_update_79975[1] = add_78772 == 32'h0000_0001 ? array_update_79973 : array_update_79962[1];
  assign array_update_79975[2] = add_78772 == 32'h0000_0002 ? array_update_79973 : array_update_79962[2];
  assign array_update_79975[3] = add_78772 == 32'h0000_0003 ? array_update_79973 : array_update_79962[3];
  assign array_update_79975[4] = add_78772 == 32'h0000_0004 ? array_update_79973 : array_update_79962[4];
  assign array_update_79975[5] = add_78772 == 32'h0000_0005 ? array_update_79973 : array_update_79962[5];
  assign array_update_79975[6] = add_78772 == 32'h0000_0006 ? array_update_79973 : array_update_79962[6];
  assign array_update_79975[7] = add_78772 == 32'h0000_0007 ? array_update_79973 : array_update_79962[7];
  assign array_update_79975[8] = add_78772 == 32'h0000_0008 ? array_update_79973 : array_update_79962[8];
  assign array_update_79975[9] = add_78772 == 32'h0000_0009 ? array_update_79973 : array_update_79962[9];
  assign array_index_79977 = array_update_72021[add_79974 > 32'h0000_0009 ? 4'h9 : add_79974[3:0]];
  assign array_index_79978 = array_update_79975[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_79982 = smul32b_32b_x_32b(array_index_78779[add_79974 > 32'h0000_0009 ? 4'h9 : add_79974[3:0]], array_index_79977[add_79855 > 32'h0000_0009 ? 4'h9 : add_79855[3:0]]);
  assign add_79984 = array_index_79978[add_79855 > 32'h0000_0009 ? 4'h9 : add_79855[3:0]] + smul_79982;
  assign array_update_79985[0] = add_79855 == 32'h0000_0000 ? add_79984 : array_index_79978[0];
  assign array_update_79985[1] = add_79855 == 32'h0000_0001 ? add_79984 : array_index_79978[1];
  assign array_update_79985[2] = add_79855 == 32'h0000_0002 ? add_79984 : array_index_79978[2];
  assign array_update_79985[3] = add_79855 == 32'h0000_0003 ? add_79984 : array_index_79978[3];
  assign array_update_79985[4] = add_79855 == 32'h0000_0004 ? add_79984 : array_index_79978[4];
  assign array_update_79985[5] = add_79855 == 32'h0000_0005 ? add_79984 : array_index_79978[5];
  assign array_update_79985[6] = add_79855 == 32'h0000_0006 ? add_79984 : array_index_79978[6];
  assign array_update_79985[7] = add_79855 == 32'h0000_0007 ? add_79984 : array_index_79978[7];
  assign array_update_79985[8] = add_79855 == 32'h0000_0008 ? add_79984 : array_index_79978[8];
  assign array_update_79985[9] = add_79855 == 32'h0000_0009 ? add_79984 : array_index_79978[9];
  assign array_update_79986[0] = add_78772 == 32'h0000_0000 ? array_update_79985 : array_update_79975[0];
  assign array_update_79986[1] = add_78772 == 32'h0000_0001 ? array_update_79985 : array_update_79975[1];
  assign array_update_79986[2] = add_78772 == 32'h0000_0002 ? array_update_79985 : array_update_79975[2];
  assign array_update_79986[3] = add_78772 == 32'h0000_0003 ? array_update_79985 : array_update_79975[3];
  assign array_update_79986[4] = add_78772 == 32'h0000_0004 ? array_update_79985 : array_update_79975[4];
  assign array_update_79986[5] = add_78772 == 32'h0000_0005 ? array_update_79985 : array_update_79975[5];
  assign array_update_79986[6] = add_78772 == 32'h0000_0006 ? array_update_79985 : array_update_79975[6];
  assign array_update_79986[7] = add_78772 == 32'h0000_0007 ? array_update_79985 : array_update_79975[7];
  assign array_update_79986[8] = add_78772 == 32'h0000_0008 ? array_update_79985 : array_update_79975[8];
  assign array_update_79986[9] = add_78772 == 32'h0000_0009 ? array_update_79985 : array_update_79975[9];
  assign array_index_79988 = array_update_79986[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign add_79990 = add_79855 + 32'h0000_0001;
  assign array_update_79991[0] = add_79990 == 32'h0000_0000 ? 32'h0000_0000 : array_index_79988[0];
  assign array_update_79991[1] = add_79990 == 32'h0000_0001 ? 32'h0000_0000 : array_index_79988[1];
  assign array_update_79991[2] = add_79990 == 32'h0000_0002 ? 32'h0000_0000 : array_index_79988[2];
  assign array_update_79991[3] = add_79990 == 32'h0000_0003 ? 32'h0000_0000 : array_index_79988[3];
  assign array_update_79991[4] = add_79990 == 32'h0000_0004 ? 32'h0000_0000 : array_index_79988[4];
  assign array_update_79991[5] = add_79990 == 32'h0000_0005 ? 32'h0000_0000 : array_index_79988[5];
  assign array_update_79991[6] = add_79990 == 32'h0000_0006 ? 32'h0000_0000 : array_index_79988[6];
  assign array_update_79991[7] = add_79990 == 32'h0000_0007 ? 32'h0000_0000 : array_index_79988[7];
  assign array_update_79991[8] = add_79990 == 32'h0000_0008 ? 32'h0000_0000 : array_index_79988[8];
  assign array_update_79991[9] = add_79990 == 32'h0000_0009 ? 32'h0000_0000 : array_index_79988[9];
  assign literal_79992 = 32'h0000_0000;
  assign array_update_79993[0] = add_78772 == 32'h0000_0000 ? array_update_79991 : array_update_79986[0];
  assign array_update_79993[1] = add_78772 == 32'h0000_0001 ? array_update_79991 : array_update_79986[1];
  assign array_update_79993[2] = add_78772 == 32'h0000_0002 ? array_update_79991 : array_update_79986[2];
  assign array_update_79993[3] = add_78772 == 32'h0000_0003 ? array_update_79991 : array_update_79986[3];
  assign array_update_79993[4] = add_78772 == 32'h0000_0004 ? array_update_79991 : array_update_79986[4];
  assign array_update_79993[5] = add_78772 == 32'h0000_0005 ? array_update_79991 : array_update_79986[5];
  assign array_update_79993[6] = add_78772 == 32'h0000_0006 ? array_update_79991 : array_update_79986[6];
  assign array_update_79993[7] = add_78772 == 32'h0000_0007 ? array_update_79991 : array_update_79986[7];
  assign array_update_79993[8] = add_78772 == 32'h0000_0008 ? array_update_79991 : array_update_79986[8];
  assign array_update_79993[9] = add_78772 == 32'h0000_0009 ? array_update_79991 : array_update_79986[9];
  assign array_index_79995 = array_update_72021[literal_79992 > 32'h0000_0009 ? 4'h9 : literal_79992[3:0]];
  assign array_index_79996 = array_update_79993[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_80000 = smul32b_32b_x_32b(array_index_78779[literal_79992 > 32'h0000_0009 ? 4'h9 : literal_79992[3:0]], array_index_79995[add_79990 > 32'h0000_0009 ? 4'h9 : add_79990[3:0]]);
  assign add_80002 = array_index_79996[add_79990 > 32'h0000_0009 ? 4'h9 : add_79990[3:0]] + smul_80000;
  assign array_update_80004[0] = add_79990 == 32'h0000_0000 ? add_80002 : array_index_79996[0];
  assign array_update_80004[1] = add_79990 == 32'h0000_0001 ? add_80002 : array_index_79996[1];
  assign array_update_80004[2] = add_79990 == 32'h0000_0002 ? add_80002 : array_index_79996[2];
  assign array_update_80004[3] = add_79990 == 32'h0000_0003 ? add_80002 : array_index_79996[3];
  assign array_update_80004[4] = add_79990 == 32'h0000_0004 ? add_80002 : array_index_79996[4];
  assign array_update_80004[5] = add_79990 == 32'h0000_0005 ? add_80002 : array_index_79996[5];
  assign array_update_80004[6] = add_79990 == 32'h0000_0006 ? add_80002 : array_index_79996[6];
  assign array_update_80004[7] = add_79990 == 32'h0000_0007 ? add_80002 : array_index_79996[7];
  assign array_update_80004[8] = add_79990 == 32'h0000_0008 ? add_80002 : array_index_79996[8];
  assign array_update_80004[9] = add_79990 == 32'h0000_0009 ? add_80002 : array_index_79996[9];
  assign add_80005 = literal_79992 + 32'h0000_0001;
  assign array_update_80006[0] = add_78772 == 32'h0000_0000 ? array_update_80004 : array_update_79993[0];
  assign array_update_80006[1] = add_78772 == 32'h0000_0001 ? array_update_80004 : array_update_79993[1];
  assign array_update_80006[2] = add_78772 == 32'h0000_0002 ? array_update_80004 : array_update_79993[2];
  assign array_update_80006[3] = add_78772 == 32'h0000_0003 ? array_update_80004 : array_update_79993[3];
  assign array_update_80006[4] = add_78772 == 32'h0000_0004 ? array_update_80004 : array_update_79993[4];
  assign array_update_80006[5] = add_78772 == 32'h0000_0005 ? array_update_80004 : array_update_79993[5];
  assign array_update_80006[6] = add_78772 == 32'h0000_0006 ? array_update_80004 : array_update_79993[6];
  assign array_update_80006[7] = add_78772 == 32'h0000_0007 ? array_update_80004 : array_update_79993[7];
  assign array_update_80006[8] = add_78772 == 32'h0000_0008 ? array_update_80004 : array_update_79993[8];
  assign array_update_80006[9] = add_78772 == 32'h0000_0009 ? array_update_80004 : array_update_79993[9];
  assign array_index_80008 = array_update_72021[add_80005 > 32'h0000_0009 ? 4'h9 : add_80005[3:0]];
  assign array_index_80009 = array_update_80006[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_80013 = smul32b_32b_x_32b(array_index_78779[add_80005 > 32'h0000_0009 ? 4'h9 : add_80005[3:0]], array_index_80008[add_79990 > 32'h0000_0009 ? 4'h9 : add_79990[3:0]]);
  assign add_80015 = array_index_80009[add_79990 > 32'h0000_0009 ? 4'h9 : add_79990[3:0]] + smul_80013;
  assign array_update_80017[0] = add_79990 == 32'h0000_0000 ? add_80015 : array_index_80009[0];
  assign array_update_80017[1] = add_79990 == 32'h0000_0001 ? add_80015 : array_index_80009[1];
  assign array_update_80017[2] = add_79990 == 32'h0000_0002 ? add_80015 : array_index_80009[2];
  assign array_update_80017[3] = add_79990 == 32'h0000_0003 ? add_80015 : array_index_80009[3];
  assign array_update_80017[4] = add_79990 == 32'h0000_0004 ? add_80015 : array_index_80009[4];
  assign array_update_80017[5] = add_79990 == 32'h0000_0005 ? add_80015 : array_index_80009[5];
  assign array_update_80017[6] = add_79990 == 32'h0000_0006 ? add_80015 : array_index_80009[6];
  assign array_update_80017[7] = add_79990 == 32'h0000_0007 ? add_80015 : array_index_80009[7];
  assign array_update_80017[8] = add_79990 == 32'h0000_0008 ? add_80015 : array_index_80009[8];
  assign array_update_80017[9] = add_79990 == 32'h0000_0009 ? add_80015 : array_index_80009[9];
  assign add_80018 = add_80005 + 32'h0000_0001;
  assign array_update_80019[0] = add_78772 == 32'h0000_0000 ? array_update_80017 : array_update_80006[0];
  assign array_update_80019[1] = add_78772 == 32'h0000_0001 ? array_update_80017 : array_update_80006[1];
  assign array_update_80019[2] = add_78772 == 32'h0000_0002 ? array_update_80017 : array_update_80006[2];
  assign array_update_80019[3] = add_78772 == 32'h0000_0003 ? array_update_80017 : array_update_80006[3];
  assign array_update_80019[4] = add_78772 == 32'h0000_0004 ? array_update_80017 : array_update_80006[4];
  assign array_update_80019[5] = add_78772 == 32'h0000_0005 ? array_update_80017 : array_update_80006[5];
  assign array_update_80019[6] = add_78772 == 32'h0000_0006 ? array_update_80017 : array_update_80006[6];
  assign array_update_80019[7] = add_78772 == 32'h0000_0007 ? array_update_80017 : array_update_80006[7];
  assign array_update_80019[8] = add_78772 == 32'h0000_0008 ? array_update_80017 : array_update_80006[8];
  assign array_update_80019[9] = add_78772 == 32'h0000_0009 ? array_update_80017 : array_update_80006[9];
  assign array_index_80021 = array_update_72021[add_80018 > 32'h0000_0009 ? 4'h9 : add_80018[3:0]];
  assign array_index_80022 = array_update_80019[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_80026 = smul32b_32b_x_32b(array_index_78779[add_80018 > 32'h0000_0009 ? 4'h9 : add_80018[3:0]], array_index_80021[add_79990 > 32'h0000_0009 ? 4'h9 : add_79990[3:0]]);
  assign add_80028 = array_index_80022[add_79990 > 32'h0000_0009 ? 4'h9 : add_79990[3:0]] + smul_80026;
  assign array_update_80030[0] = add_79990 == 32'h0000_0000 ? add_80028 : array_index_80022[0];
  assign array_update_80030[1] = add_79990 == 32'h0000_0001 ? add_80028 : array_index_80022[1];
  assign array_update_80030[2] = add_79990 == 32'h0000_0002 ? add_80028 : array_index_80022[2];
  assign array_update_80030[3] = add_79990 == 32'h0000_0003 ? add_80028 : array_index_80022[3];
  assign array_update_80030[4] = add_79990 == 32'h0000_0004 ? add_80028 : array_index_80022[4];
  assign array_update_80030[5] = add_79990 == 32'h0000_0005 ? add_80028 : array_index_80022[5];
  assign array_update_80030[6] = add_79990 == 32'h0000_0006 ? add_80028 : array_index_80022[6];
  assign array_update_80030[7] = add_79990 == 32'h0000_0007 ? add_80028 : array_index_80022[7];
  assign array_update_80030[8] = add_79990 == 32'h0000_0008 ? add_80028 : array_index_80022[8];
  assign array_update_80030[9] = add_79990 == 32'h0000_0009 ? add_80028 : array_index_80022[9];
  assign add_80031 = add_80018 + 32'h0000_0001;
  assign array_update_80032[0] = add_78772 == 32'h0000_0000 ? array_update_80030 : array_update_80019[0];
  assign array_update_80032[1] = add_78772 == 32'h0000_0001 ? array_update_80030 : array_update_80019[1];
  assign array_update_80032[2] = add_78772 == 32'h0000_0002 ? array_update_80030 : array_update_80019[2];
  assign array_update_80032[3] = add_78772 == 32'h0000_0003 ? array_update_80030 : array_update_80019[3];
  assign array_update_80032[4] = add_78772 == 32'h0000_0004 ? array_update_80030 : array_update_80019[4];
  assign array_update_80032[5] = add_78772 == 32'h0000_0005 ? array_update_80030 : array_update_80019[5];
  assign array_update_80032[6] = add_78772 == 32'h0000_0006 ? array_update_80030 : array_update_80019[6];
  assign array_update_80032[7] = add_78772 == 32'h0000_0007 ? array_update_80030 : array_update_80019[7];
  assign array_update_80032[8] = add_78772 == 32'h0000_0008 ? array_update_80030 : array_update_80019[8];
  assign array_update_80032[9] = add_78772 == 32'h0000_0009 ? array_update_80030 : array_update_80019[9];
  assign array_index_80034 = array_update_72021[add_80031 > 32'h0000_0009 ? 4'h9 : add_80031[3:0]];
  assign array_index_80035 = array_update_80032[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_80039 = smul32b_32b_x_32b(array_index_78779[add_80031 > 32'h0000_0009 ? 4'h9 : add_80031[3:0]], array_index_80034[add_79990 > 32'h0000_0009 ? 4'h9 : add_79990[3:0]]);
  assign add_80041 = array_index_80035[add_79990 > 32'h0000_0009 ? 4'h9 : add_79990[3:0]] + smul_80039;
  assign array_update_80043[0] = add_79990 == 32'h0000_0000 ? add_80041 : array_index_80035[0];
  assign array_update_80043[1] = add_79990 == 32'h0000_0001 ? add_80041 : array_index_80035[1];
  assign array_update_80043[2] = add_79990 == 32'h0000_0002 ? add_80041 : array_index_80035[2];
  assign array_update_80043[3] = add_79990 == 32'h0000_0003 ? add_80041 : array_index_80035[3];
  assign array_update_80043[4] = add_79990 == 32'h0000_0004 ? add_80041 : array_index_80035[4];
  assign array_update_80043[5] = add_79990 == 32'h0000_0005 ? add_80041 : array_index_80035[5];
  assign array_update_80043[6] = add_79990 == 32'h0000_0006 ? add_80041 : array_index_80035[6];
  assign array_update_80043[7] = add_79990 == 32'h0000_0007 ? add_80041 : array_index_80035[7];
  assign array_update_80043[8] = add_79990 == 32'h0000_0008 ? add_80041 : array_index_80035[8];
  assign array_update_80043[9] = add_79990 == 32'h0000_0009 ? add_80041 : array_index_80035[9];
  assign add_80044 = add_80031 + 32'h0000_0001;
  assign array_update_80045[0] = add_78772 == 32'h0000_0000 ? array_update_80043 : array_update_80032[0];
  assign array_update_80045[1] = add_78772 == 32'h0000_0001 ? array_update_80043 : array_update_80032[1];
  assign array_update_80045[2] = add_78772 == 32'h0000_0002 ? array_update_80043 : array_update_80032[2];
  assign array_update_80045[3] = add_78772 == 32'h0000_0003 ? array_update_80043 : array_update_80032[3];
  assign array_update_80045[4] = add_78772 == 32'h0000_0004 ? array_update_80043 : array_update_80032[4];
  assign array_update_80045[5] = add_78772 == 32'h0000_0005 ? array_update_80043 : array_update_80032[5];
  assign array_update_80045[6] = add_78772 == 32'h0000_0006 ? array_update_80043 : array_update_80032[6];
  assign array_update_80045[7] = add_78772 == 32'h0000_0007 ? array_update_80043 : array_update_80032[7];
  assign array_update_80045[8] = add_78772 == 32'h0000_0008 ? array_update_80043 : array_update_80032[8];
  assign array_update_80045[9] = add_78772 == 32'h0000_0009 ? array_update_80043 : array_update_80032[9];
  assign array_index_80047 = array_update_72021[add_80044 > 32'h0000_0009 ? 4'h9 : add_80044[3:0]];
  assign array_index_80048 = array_update_80045[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_80052 = smul32b_32b_x_32b(array_index_78779[add_80044 > 32'h0000_0009 ? 4'h9 : add_80044[3:0]], array_index_80047[add_79990 > 32'h0000_0009 ? 4'h9 : add_79990[3:0]]);
  assign add_80054 = array_index_80048[add_79990 > 32'h0000_0009 ? 4'h9 : add_79990[3:0]] + smul_80052;
  assign array_update_80056[0] = add_79990 == 32'h0000_0000 ? add_80054 : array_index_80048[0];
  assign array_update_80056[1] = add_79990 == 32'h0000_0001 ? add_80054 : array_index_80048[1];
  assign array_update_80056[2] = add_79990 == 32'h0000_0002 ? add_80054 : array_index_80048[2];
  assign array_update_80056[3] = add_79990 == 32'h0000_0003 ? add_80054 : array_index_80048[3];
  assign array_update_80056[4] = add_79990 == 32'h0000_0004 ? add_80054 : array_index_80048[4];
  assign array_update_80056[5] = add_79990 == 32'h0000_0005 ? add_80054 : array_index_80048[5];
  assign array_update_80056[6] = add_79990 == 32'h0000_0006 ? add_80054 : array_index_80048[6];
  assign array_update_80056[7] = add_79990 == 32'h0000_0007 ? add_80054 : array_index_80048[7];
  assign array_update_80056[8] = add_79990 == 32'h0000_0008 ? add_80054 : array_index_80048[8];
  assign array_update_80056[9] = add_79990 == 32'h0000_0009 ? add_80054 : array_index_80048[9];
  assign add_80057 = add_80044 + 32'h0000_0001;
  assign array_update_80058[0] = add_78772 == 32'h0000_0000 ? array_update_80056 : array_update_80045[0];
  assign array_update_80058[1] = add_78772 == 32'h0000_0001 ? array_update_80056 : array_update_80045[1];
  assign array_update_80058[2] = add_78772 == 32'h0000_0002 ? array_update_80056 : array_update_80045[2];
  assign array_update_80058[3] = add_78772 == 32'h0000_0003 ? array_update_80056 : array_update_80045[3];
  assign array_update_80058[4] = add_78772 == 32'h0000_0004 ? array_update_80056 : array_update_80045[4];
  assign array_update_80058[5] = add_78772 == 32'h0000_0005 ? array_update_80056 : array_update_80045[5];
  assign array_update_80058[6] = add_78772 == 32'h0000_0006 ? array_update_80056 : array_update_80045[6];
  assign array_update_80058[7] = add_78772 == 32'h0000_0007 ? array_update_80056 : array_update_80045[7];
  assign array_update_80058[8] = add_78772 == 32'h0000_0008 ? array_update_80056 : array_update_80045[8];
  assign array_update_80058[9] = add_78772 == 32'h0000_0009 ? array_update_80056 : array_update_80045[9];
  assign array_index_80060 = array_update_72021[add_80057 > 32'h0000_0009 ? 4'h9 : add_80057[3:0]];
  assign array_index_80061 = array_update_80058[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_80065 = smul32b_32b_x_32b(array_index_78779[add_80057 > 32'h0000_0009 ? 4'h9 : add_80057[3:0]], array_index_80060[add_79990 > 32'h0000_0009 ? 4'h9 : add_79990[3:0]]);
  assign add_80067 = array_index_80061[add_79990 > 32'h0000_0009 ? 4'h9 : add_79990[3:0]] + smul_80065;
  assign array_update_80069[0] = add_79990 == 32'h0000_0000 ? add_80067 : array_index_80061[0];
  assign array_update_80069[1] = add_79990 == 32'h0000_0001 ? add_80067 : array_index_80061[1];
  assign array_update_80069[2] = add_79990 == 32'h0000_0002 ? add_80067 : array_index_80061[2];
  assign array_update_80069[3] = add_79990 == 32'h0000_0003 ? add_80067 : array_index_80061[3];
  assign array_update_80069[4] = add_79990 == 32'h0000_0004 ? add_80067 : array_index_80061[4];
  assign array_update_80069[5] = add_79990 == 32'h0000_0005 ? add_80067 : array_index_80061[5];
  assign array_update_80069[6] = add_79990 == 32'h0000_0006 ? add_80067 : array_index_80061[6];
  assign array_update_80069[7] = add_79990 == 32'h0000_0007 ? add_80067 : array_index_80061[7];
  assign array_update_80069[8] = add_79990 == 32'h0000_0008 ? add_80067 : array_index_80061[8];
  assign array_update_80069[9] = add_79990 == 32'h0000_0009 ? add_80067 : array_index_80061[9];
  assign add_80070 = add_80057 + 32'h0000_0001;
  assign array_update_80071[0] = add_78772 == 32'h0000_0000 ? array_update_80069 : array_update_80058[0];
  assign array_update_80071[1] = add_78772 == 32'h0000_0001 ? array_update_80069 : array_update_80058[1];
  assign array_update_80071[2] = add_78772 == 32'h0000_0002 ? array_update_80069 : array_update_80058[2];
  assign array_update_80071[3] = add_78772 == 32'h0000_0003 ? array_update_80069 : array_update_80058[3];
  assign array_update_80071[4] = add_78772 == 32'h0000_0004 ? array_update_80069 : array_update_80058[4];
  assign array_update_80071[5] = add_78772 == 32'h0000_0005 ? array_update_80069 : array_update_80058[5];
  assign array_update_80071[6] = add_78772 == 32'h0000_0006 ? array_update_80069 : array_update_80058[6];
  assign array_update_80071[7] = add_78772 == 32'h0000_0007 ? array_update_80069 : array_update_80058[7];
  assign array_update_80071[8] = add_78772 == 32'h0000_0008 ? array_update_80069 : array_update_80058[8];
  assign array_update_80071[9] = add_78772 == 32'h0000_0009 ? array_update_80069 : array_update_80058[9];
  assign array_index_80073 = array_update_72021[add_80070 > 32'h0000_0009 ? 4'h9 : add_80070[3:0]];
  assign array_index_80074 = array_update_80071[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_80078 = smul32b_32b_x_32b(array_index_78779[add_80070 > 32'h0000_0009 ? 4'h9 : add_80070[3:0]], array_index_80073[add_79990 > 32'h0000_0009 ? 4'h9 : add_79990[3:0]]);
  assign add_80080 = array_index_80074[add_79990 > 32'h0000_0009 ? 4'h9 : add_79990[3:0]] + smul_80078;
  assign array_update_80082[0] = add_79990 == 32'h0000_0000 ? add_80080 : array_index_80074[0];
  assign array_update_80082[1] = add_79990 == 32'h0000_0001 ? add_80080 : array_index_80074[1];
  assign array_update_80082[2] = add_79990 == 32'h0000_0002 ? add_80080 : array_index_80074[2];
  assign array_update_80082[3] = add_79990 == 32'h0000_0003 ? add_80080 : array_index_80074[3];
  assign array_update_80082[4] = add_79990 == 32'h0000_0004 ? add_80080 : array_index_80074[4];
  assign array_update_80082[5] = add_79990 == 32'h0000_0005 ? add_80080 : array_index_80074[5];
  assign array_update_80082[6] = add_79990 == 32'h0000_0006 ? add_80080 : array_index_80074[6];
  assign array_update_80082[7] = add_79990 == 32'h0000_0007 ? add_80080 : array_index_80074[7];
  assign array_update_80082[8] = add_79990 == 32'h0000_0008 ? add_80080 : array_index_80074[8];
  assign array_update_80082[9] = add_79990 == 32'h0000_0009 ? add_80080 : array_index_80074[9];
  assign add_80083 = add_80070 + 32'h0000_0001;
  assign array_update_80084[0] = add_78772 == 32'h0000_0000 ? array_update_80082 : array_update_80071[0];
  assign array_update_80084[1] = add_78772 == 32'h0000_0001 ? array_update_80082 : array_update_80071[1];
  assign array_update_80084[2] = add_78772 == 32'h0000_0002 ? array_update_80082 : array_update_80071[2];
  assign array_update_80084[3] = add_78772 == 32'h0000_0003 ? array_update_80082 : array_update_80071[3];
  assign array_update_80084[4] = add_78772 == 32'h0000_0004 ? array_update_80082 : array_update_80071[4];
  assign array_update_80084[5] = add_78772 == 32'h0000_0005 ? array_update_80082 : array_update_80071[5];
  assign array_update_80084[6] = add_78772 == 32'h0000_0006 ? array_update_80082 : array_update_80071[6];
  assign array_update_80084[7] = add_78772 == 32'h0000_0007 ? array_update_80082 : array_update_80071[7];
  assign array_update_80084[8] = add_78772 == 32'h0000_0008 ? array_update_80082 : array_update_80071[8];
  assign array_update_80084[9] = add_78772 == 32'h0000_0009 ? array_update_80082 : array_update_80071[9];
  assign array_index_80086 = array_update_72021[add_80083 > 32'h0000_0009 ? 4'h9 : add_80083[3:0]];
  assign array_index_80087 = array_update_80084[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_80091 = smul32b_32b_x_32b(array_index_78779[add_80083 > 32'h0000_0009 ? 4'h9 : add_80083[3:0]], array_index_80086[add_79990 > 32'h0000_0009 ? 4'h9 : add_79990[3:0]]);
  assign add_80093 = array_index_80087[add_79990 > 32'h0000_0009 ? 4'h9 : add_79990[3:0]] + smul_80091;
  assign array_update_80095[0] = add_79990 == 32'h0000_0000 ? add_80093 : array_index_80087[0];
  assign array_update_80095[1] = add_79990 == 32'h0000_0001 ? add_80093 : array_index_80087[1];
  assign array_update_80095[2] = add_79990 == 32'h0000_0002 ? add_80093 : array_index_80087[2];
  assign array_update_80095[3] = add_79990 == 32'h0000_0003 ? add_80093 : array_index_80087[3];
  assign array_update_80095[4] = add_79990 == 32'h0000_0004 ? add_80093 : array_index_80087[4];
  assign array_update_80095[5] = add_79990 == 32'h0000_0005 ? add_80093 : array_index_80087[5];
  assign array_update_80095[6] = add_79990 == 32'h0000_0006 ? add_80093 : array_index_80087[6];
  assign array_update_80095[7] = add_79990 == 32'h0000_0007 ? add_80093 : array_index_80087[7];
  assign array_update_80095[8] = add_79990 == 32'h0000_0008 ? add_80093 : array_index_80087[8];
  assign array_update_80095[9] = add_79990 == 32'h0000_0009 ? add_80093 : array_index_80087[9];
  assign add_80096 = add_80083 + 32'h0000_0001;
  assign array_update_80097[0] = add_78772 == 32'h0000_0000 ? array_update_80095 : array_update_80084[0];
  assign array_update_80097[1] = add_78772 == 32'h0000_0001 ? array_update_80095 : array_update_80084[1];
  assign array_update_80097[2] = add_78772 == 32'h0000_0002 ? array_update_80095 : array_update_80084[2];
  assign array_update_80097[3] = add_78772 == 32'h0000_0003 ? array_update_80095 : array_update_80084[3];
  assign array_update_80097[4] = add_78772 == 32'h0000_0004 ? array_update_80095 : array_update_80084[4];
  assign array_update_80097[5] = add_78772 == 32'h0000_0005 ? array_update_80095 : array_update_80084[5];
  assign array_update_80097[6] = add_78772 == 32'h0000_0006 ? array_update_80095 : array_update_80084[6];
  assign array_update_80097[7] = add_78772 == 32'h0000_0007 ? array_update_80095 : array_update_80084[7];
  assign array_update_80097[8] = add_78772 == 32'h0000_0008 ? array_update_80095 : array_update_80084[8];
  assign array_update_80097[9] = add_78772 == 32'h0000_0009 ? array_update_80095 : array_update_80084[9];
  assign array_index_80099 = array_update_72021[add_80096 > 32'h0000_0009 ? 4'h9 : add_80096[3:0]];
  assign array_index_80100 = array_update_80097[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_80104 = smul32b_32b_x_32b(array_index_78779[add_80096 > 32'h0000_0009 ? 4'h9 : add_80096[3:0]], array_index_80099[add_79990 > 32'h0000_0009 ? 4'h9 : add_79990[3:0]]);
  assign add_80106 = array_index_80100[add_79990 > 32'h0000_0009 ? 4'h9 : add_79990[3:0]] + smul_80104;
  assign array_update_80108[0] = add_79990 == 32'h0000_0000 ? add_80106 : array_index_80100[0];
  assign array_update_80108[1] = add_79990 == 32'h0000_0001 ? add_80106 : array_index_80100[1];
  assign array_update_80108[2] = add_79990 == 32'h0000_0002 ? add_80106 : array_index_80100[2];
  assign array_update_80108[3] = add_79990 == 32'h0000_0003 ? add_80106 : array_index_80100[3];
  assign array_update_80108[4] = add_79990 == 32'h0000_0004 ? add_80106 : array_index_80100[4];
  assign array_update_80108[5] = add_79990 == 32'h0000_0005 ? add_80106 : array_index_80100[5];
  assign array_update_80108[6] = add_79990 == 32'h0000_0006 ? add_80106 : array_index_80100[6];
  assign array_update_80108[7] = add_79990 == 32'h0000_0007 ? add_80106 : array_index_80100[7];
  assign array_update_80108[8] = add_79990 == 32'h0000_0008 ? add_80106 : array_index_80100[8];
  assign array_update_80108[9] = add_79990 == 32'h0000_0009 ? add_80106 : array_index_80100[9];
  assign add_80109 = add_80096 + 32'h0000_0001;
  assign array_update_80110[0] = add_78772 == 32'h0000_0000 ? array_update_80108 : array_update_80097[0];
  assign array_update_80110[1] = add_78772 == 32'h0000_0001 ? array_update_80108 : array_update_80097[1];
  assign array_update_80110[2] = add_78772 == 32'h0000_0002 ? array_update_80108 : array_update_80097[2];
  assign array_update_80110[3] = add_78772 == 32'h0000_0003 ? array_update_80108 : array_update_80097[3];
  assign array_update_80110[4] = add_78772 == 32'h0000_0004 ? array_update_80108 : array_update_80097[4];
  assign array_update_80110[5] = add_78772 == 32'h0000_0005 ? array_update_80108 : array_update_80097[5];
  assign array_update_80110[6] = add_78772 == 32'h0000_0006 ? array_update_80108 : array_update_80097[6];
  assign array_update_80110[7] = add_78772 == 32'h0000_0007 ? array_update_80108 : array_update_80097[7];
  assign array_update_80110[8] = add_78772 == 32'h0000_0008 ? array_update_80108 : array_update_80097[8];
  assign array_update_80110[9] = add_78772 == 32'h0000_0009 ? array_update_80108 : array_update_80097[9];
  assign array_index_80112 = array_update_72021[add_80109 > 32'h0000_0009 ? 4'h9 : add_80109[3:0]];
  assign array_index_80113 = array_update_80110[add_78772 > 32'h0000_0009 ? 4'h9 : add_78772[3:0]];
  assign smul_80117 = smul32b_32b_x_32b(array_index_78779[add_80109 > 32'h0000_0009 ? 4'h9 : add_80109[3:0]], array_index_80112[add_79990 > 32'h0000_0009 ? 4'h9 : add_79990[3:0]]);
  assign add_80119 = array_index_80113[add_79990 > 32'h0000_0009 ? 4'h9 : add_79990[3:0]] + smul_80117;
  assign array_update_80120[0] = add_79990 == 32'h0000_0000 ? add_80119 : array_index_80113[0];
  assign array_update_80120[1] = add_79990 == 32'h0000_0001 ? add_80119 : array_index_80113[1];
  assign array_update_80120[2] = add_79990 == 32'h0000_0002 ? add_80119 : array_index_80113[2];
  assign array_update_80120[3] = add_79990 == 32'h0000_0003 ? add_80119 : array_index_80113[3];
  assign array_update_80120[4] = add_79990 == 32'h0000_0004 ? add_80119 : array_index_80113[4];
  assign array_update_80120[5] = add_79990 == 32'h0000_0005 ? add_80119 : array_index_80113[5];
  assign array_update_80120[6] = add_79990 == 32'h0000_0006 ? add_80119 : array_index_80113[6];
  assign array_update_80120[7] = add_79990 == 32'h0000_0007 ? add_80119 : array_index_80113[7];
  assign array_update_80120[8] = add_79990 == 32'h0000_0008 ? add_80119 : array_index_80113[8];
  assign array_update_80120[9] = add_79990 == 32'h0000_0009 ? add_80119 : array_index_80113[9];
  assign array_update_80122[0] = add_78772 == 32'h0000_0000 ? array_update_80120 : array_update_80110[0];
  assign array_update_80122[1] = add_78772 == 32'h0000_0001 ? array_update_80120 : array_update_80110[1];
  assign array_update_80122[2] = add_78772 == 32'h0000_0002 ? array_update_80120 : array_update_80110[2];
  assign array_update_80122[3] = add_78772 == 32'h0000_0003 ? array_update_80120 : array_update_80110[3];
  assign array_update_80122[4] = add_78772 == 32'h0000_0004 ? array_update_80120 : array_update_80110[4];
  assign array_update_80122[5] = add_78772 == 32'h0000_0005 ? array_update_80120 : array_update_80110[5];
  assign array_update_80122[6] = add_78772 == 32'h0000_0006 ? array_update_80120 : array_update_80110[6];
  assign array_update_80122[7] = add_78772 == 32'h0000_0007 ? array_update_80120 : array_update_80110[7];
  assign array_update_80122[8] = add_78772 == 32'h0000_0008 ? array_update_80120 : array_update_80110[8];
  assign array_update_80122[9] = add_78772 == 32'h0000_0009 ? array_update_80120 : array_update_80110[9];
  assign add_80123 = add_78772 + 32'h0000_0001;
  assign array_index_80124 = array_update_80122[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign literal_80126 = 32'h0000_0000;
  assign array_update_80127[0] = literal_80126 == 32'h0000_0000 ? 32'h0000_0000 : array_index_80124[0];
  assign array_update_80127[1] = literal_80126 == 32'h0000_0001 ? 32'h0000_0000 : array_index_80124[1];
  assign array_update_80127[2] = literal_80126 == 32'h0000_0002 ? 32'h0000_0000 : array_index_80124[2];
  assign array_update_80127[3] = literal_80126 == 32'h0000_0003 ? 32'h0000_0000 : array_index_80124[3];
  assign array_update_80127[4] = literal_80126 == 32'h0000_0004 ? 32'h0000_0000 : array_index_80124[4];
  assign array_update_80127[5] = literal_80126 == 32'h0000_0005 ? 32'h0000_0000 : array_index_80124[5];
  assign array_update_80127[6] = literal_80126 == 32'h0000_0006 ? 32'h0000_0000 : array_index_80124[6];
  assign array_update_80127[7] = literal_80126 == 32'h0000_0007 ? 32'h0000_0000 : array_index_80124[7];
  assign array_update_80127[8] = literal_80126 == 32'h0000_0008 ? 32'h0000_0000 : array_index_80124[8];
  assign array_update_80127[9] = literal_80126 == 32'h0000_0009 ? 32'h0000_0000 : array_index_80124[9];
  assign literal_80128 = 32'h0000_0000;
  assign array_update_80129[0] = add_80123 == 32'h0000_0000 ? array_update_80127 : array_update_80122[0];
  assign array_update_80129[1] = add_80123 == 32'h0000_0001 ? array_update_80127 : array_update_80122[1];
  assign array_update_80129[2] = add_80123 == 32'h0000_0002 ? array_update_80127 : array_update_80122[2];
  assign array_update_80129[3] = add_80123 == 32'h0000_0003 ? array_update_80127 : array_update_80122[3];
  assign array_update_80129[4] = add_80123 == 32'h0000_0004 ? array_update_80127 : array_update_80122[4];
  assign array_update_80129[5] = add_80123 == 32'h0000_0005 ? array_update_80127 : array_update_80122[5];
  assign array_update_80129[6] = add_80123 == 32'h0000_0006 ? array_update_80127 : array_update_80122[6];
  assign array_update_80129[7] = add_80123 == 32'h0000_0007 ? array_update_80127 : array_update_80122[7];
  assign array_update_80129[8] = add_80123 == 32'h0000_0008 ? array_update_80127 : array_update_80122[8];
  assign array_update_80129[9] = add_80123 == 32'h0000_0009 ? array_update_80127 : array_update_80122[9];
  assign array_index_80130 = array_update_72020[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign array_index_80131 = array_update_72021[literal_80128 > 32'h0000_0009 ? 4'h9 : literal_80128[3:0]];
  assign array_index_80132 = array_update_80129[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_80136 = smul32b_32b_x_32b(array_index_80130[literal_80128 > 32'h0000_0009 ? 4'h9 : literal_80128[3:0]], array_index_80131[literal_80126 > 32'h0000_0009 ? 4'h9 : literal_80126[3:0]]);
  assign add_80138 = array_index_80132[literal_80126 > 32'h0000_0009 ? 4'h9 : literal_80126[3:0]] + smul_80136;
  assign array_update_80140[0] = literal_80126 == 32'h0000_0000 ? add_80138 : array_index_80132[0];
  assign array_update_80140[1] = literal_80126 == 32'h0000_0001 ? add_80138 : array_index_80132[1];
  assign array_update_80140[2] = literal_80126 == 32'h0000_0002 ? add_80138 : array_index_80132[2];
  assign array_update_80140[3] = literal_80126 == 32'h0000_0003 ? add_80138 : array_index_80132[3];
  assign array_update_80140[4] = literal_80126 == 32'h0000_0004 ? add_80138 : array_index_80132[4];
  assign array_update_80140[5] = literal_80126 == 32'h0000_0005 ? add_80138 : array_index_80132[5];
  assign array_update_80140[6] = literal_80126 == 32'h0000_0006 ? add_80138 : array_index_80132[6];
  assign array_update_80140[7] = literal_80126 == 32'h0000_0007 ? add_80138 : array_index_80132[7];
  assign array_update_80140[8] = literal_80126 == 32'h0000_0008 ? add_80138 : array_index_80132[8];
  assign array_update_80140[9] = literal_80126 == 32'h0000_0009 ? add_80138 : array_index_80132[9];
  assign add_80141 = literal_80128 + 32'h0000_0001;
  assign array_update_80142[0] = add_80123 == 32'h0000_0000 ? array_update_80140 : array_update_80129[0];
  assign array_update_80142[1] = add_80123 == 32'h0000_0001 ? array_update_80140 : array_update_80129[1];
  assign array_update_80142[2] = add_80123 == 32'h0000_0002 ? array_update_80140 : array_update_80129[2];
  assign array_update_80142[3] = add_80123 == 32'h0000_0003 ? array_update_80140 : array_update_80129[3];
  assign array_update_80142[4] = add_80123 == 32'h0000_0004 ? array_update_80140 : array_update_80129[4];
  assign array_update_80142[5] = add_80123 == 32'h0000_0005 ? array_update_80140 : array_update_80129[5];
  assign array_update_80142[6] = add_80123 == 32'h0000_0006 ? array_update_80140 : array_update_80129[6];
  assign array_update_80142[7] = add_80123 == 32'h0000_0007 ? array_update_80140 : array_update_80129[7];
  assign array_update_80142[8] = add_80123 == 32'h0000_0008 ? array_update_80140 : array_update_80129[8];
  assign array_update_80142[9] = add_80123 == 32'h0000_0009 ? array_update_80140 : array_update_80129[9];
  assign array_index_80144 = array_update_72021[add_80141 > 32'h0000_0009 ? 4'h9 : add_80141[3:0]];
  assign array_index_80145 = array_update_80142[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_80149 = smul32b_32b_x_32b(array_index_80130[add_80141 > 32'h0000_0009 ? 4'h9 : add_80141[3:0]], array_index_80144[literal_80126 > 32'h0000_0009 ? 4'h9 : literal_80126[3:0]]);
  assign add_80151 = array_index_80145[literal_80126 > 32'h0000_0009 ? 4'h9 : literal_80126[3:0]] + smul_80149;
  assign array_update_80153[0] = literal_80126 == 32'h0000_0000 ? add_80151 : array_index_80145[0];
  assign array_update_80153[1] = literal_80126 == 32'h0000_0001 ? add_80151 : array_index_80145[1];
  assign array_update_80153[2] = literal_80126 == 32'h0000_0002 ? add_80151 : array_index_80145[2];
  assign array_update_80153[3] = literal_80126 == 32'h0000_0003 ? add_80151 : array_index_80145[3];
  assign array_update_80153[4] = literal_80126 == 32'h0000_0004 ? add_80151 : array_index_80145[4];
  assign array_update_80153[5] = literal_80126 == 32'h0000_0005 ? add_80151 : array_index_80145[5];
  assign array_update_80153[6] = literal_80126 == 32'h0000_0006 ? add_80151 : array_index_80145[6];
  assign array_update_80153[7] = literal_80126 == 32'h0000_0007 ? add_80151 : array_index_80145[7];
  assign array_update_80153[8] = literal_80126 == 32'h0000_0008 ? add_80151 : array_index_80145[8];
  assign array_update_80153[9] = literal_80126 == 32'h0000_0009 ? add_80151 : array_index_80145[9];
  assign add_80154 = add_80141 + 32'h0000_0001;
  assign array_update_80155[0] = add_80123 == 32'h0000_0000 ? array_update_80153 : array_update_80142[0];
  assign array_update_80155[1] = add_80123 == 32'h0000_0001 ? array_update_80153 : array_update_80142[1];
  assign array_update_80155[2] = add_80123 == 32'h0000_0002 ? array_update_80153 : array_update_80142[2];
  assign array_update_80155[3] = add_80123 == 32'h0000_0003 ? array_update_80153 : array_update_80142[3];
  assign array_update_80155[4] = add_80123 == 32'h0000_0004 ? array_update_80153 : array_update_80142[4];
  assign array_update_80155[5] = add_80123 == 32'h0000_0005 ? array_update_80153 : array_update_80142[5];
  assign array_update_80155[6] = add_80123 == 32'h0000_0006 ? array_update_80153 : array_update_80142[6];
  assign array_update_80155[7] = add_80123 == 32'h0000_0007 ? array_update_80153 : array_update_80142[7];
  assign array_update_80155[8] = add_80123 == 32'h0000_0008 ? array_update_80153 : array_update_80142[8];
  assign array_update_80155[9] = add_80123 == 32'h0000_0009 ? array_update_80153 : array_update_80142[9];
  assign array_index_80157 = array_update_72021[add_80154 > 32'h0000_0009 ? 4'h9 : add_80154[3:0]];
  assign array_index_80158 = array_update_80155[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_80162 = smul32b_32b_x_32b(array_index_80130[add_80154 > 32'h0000_0009 ? 4'h9 : add_80154[3:0]], array_index_80157[literal_80126 > 32'h0000_0009 ? 4'h9 : literal_80126[3:0]]);
  assign add_80164 = array_index_80158[literal_80126 > 32'h0000_0009 ? 4'h9 : literal_80126[3:0]] + smul_80162;
  assign array_update_80166[0] = literal_80126 == 32'h0000_0000 ? add_80164 : array_index_80158[0];
  assign array_update_80166[1] = literal_80126 == 32'h0000_0001 ? add_80164 : array_index_80158[1];
  assign array_update_80166[2] = literal_80126 == 32'h0000_0002 ? add_80164 : array_index_80158[2];
  assign array_update_80166[3] = literal_80126 == 32'h0000_0003 ? add_80164 : array_index_80158[3];
  assign array_update_80166[4] = literal_80126 == 32'h0000_0004 ? add_80164 : array_index_80158[4];
  assign array_update_80166[5] = literal_80126 == 32'h0000_0005 ? add_80164 : array_index_80158[5];
  assign array_update_80166[6] = literal_80126 == 32'h0000_0006 ? add_80164 : array_index_80158[6];
  assign array_update_80166[7] = literal_80126 == 32'h0000_0007 ? add_80164 : array_index_80158[7];
  assign array_update_80166[8] = literal_80126 == 32'h0000_0008 ? add_80164 : array_index_80158[8];
  assign array_update_80166[9] = literal_80126 == 32'h0000_0009 ? add_80164 : array_index_80158[9];
  assign add_80167 = add_80154 + 32'h0000_0001;
  assign array_update_80168[0] = add_80123 == 32'h0000_0000 ? array_update_80166 : array_update_80155[0];
  assign array_update_80168[1] = add_80123 == 32'h0000_0001 ? array_update_80166 : array_update_80155[1];
  assign array_update_80168[2] = add_80123 == 32'h0000_0002 ? array_update_80166 : array_update_80155[2];
  assign array_update_80168[3] = add_80123 == 32'h0000_0003 ? array_update_80166 : array_update_80155[3];
  assign array_update_80168[4] = add_80123 == 32'h0000_0004 ? array_update_80166 : array_update_80155[4];
  assign array_update_80168[5] = add_80123 == 32'h0000_0005 ? array_update_80166 : array_update_80155[5];
  assign array_update_80168[6] = add_80123 == 32'h0000_0006 ? array_update_80166 : array_update_80155[6];
  assign array_update_80168[7] = add_80123 == 32'h0000_0007 ? array_update_80166 : array_update_80155[7];
  assign array_update_80168[8] = add_80123 == 32'h0000_0008 ? array_update_80166 : array_update_80155[8];
  assign array_update_80168[9] = add_80123 == 32'h0000_0009 ? array_update_80166 : array_update_80155[9];
  assign array_index_80170 = array_update_72021[add_80167 > 32'h0000_0009 ? 4'h9 : add_80167[3:0]];
  assign array_index_80171 = array_update_80168[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_80175 = smul32b_32b_x_32b(array_index_80130[add_80167 > 32'h0000_0009 ? 4'h9 : add_80167[3:0]], array_index_80170[literal_80126 > 32'h0000_0009 ? 4'h9 : literal_80126[3:0]]);
  assign add_80177 = array_index_80171[literal_80126 > 32'h0000_0009 ? 4'h9 : literal_80126[3:0]] + smul_80175;
  assign array_update_80179[0] = literal_80126 == 32'h0000_0000 ? add_80177 : array_index_80171[0];
  assign array_update_80179[1] = literal_80126 == 32'h0000_0001 ? add_80177 : array_index_80171[1];
  assign array_update_80179[2] = literal_80126 == 32'h0000_0002 ? add_80177 : array_index_80171[2];
  assign array_update_80179[3] = literal_80126 == 32'h0000_0003 ? add_80177 : array_index_80171[3];
  assign array_update_80179[4] = literal_80126 == 32'h0000_0004 ? add_80177 : array_index_80171[4];
  assign array_update_80179[5] = literal_80126 == 32'h0000_0005 ? add_80177 : array_index_80171[5];
  assign array_update_80179[6] = literal_80126 == 32'h0000_0006 ? add_80177 : array_index_80171[6];
  assign array_update_80179[7] = literal_80126 == 32'h0000_0007 ? add_80177 : array_index_80171[7];
  assign array_update_80179[8] = literal_80126 == 32'h0000_0008 ? add_80177 : array_index_80171[8];
  assign array_update_80179[9] = literal_80126 == 32'h0000_0009 ? add_80177 : array_index_80171[9];
  assign add_80180 = add_80167 + 32'h0000_0001;
  assign array_update_80181[0] = add_80123 == 32'h0000_0000 ? array_update_80179 : array_update_80168[0];
  assign array_update_80181[1] = add_80123 == 32'h0000_0001 ? array_update_80179 : array_update_80168[1];
  assign array_update_80181[2] = add_80123 == 32'h0000_0002 ? array_update_80179 : array_update_80168[2];
  assign array_update_80181[3] = add_80123 == 32'h0000_0003 ? array_update_80179 : array_update_80168[3];
  assign array_update_80181[4] = add_80123 == 32'h0000_0004 ? array_update_80179 : array_update_80168[4];
  assign array_update_80181[5] = add_80123 == 32'h0000_0005 ? array_update_80179 : array_update_80168[5];
  assign array_update_80181[6] = add_80123 == 32'h0000_0006 ? array_update_80179 : array_update_80168[6];
  assign array_update_80181[7] = add_80123 == 32'h0000_0007 ? array_update_80179 : array_update_80168[7];
  assign array_update_80181[8] = add_80123 == 32'h0000_0008 ? array_update_80179 : array_update_80168[8];
  assign array_update_80181[9] = add_80123 == 32'h0000_0009 ? array_update_80179 : array_update_80168[9];
  assign array_index_80183 = array_update_72021[add_80180 > 32'h0000_0009 ? 4'h9 : add_80180[3:0]];
  assign array_index_80184 = array_update_80181[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_80188 = smul32b_32b_x_32b(array_index_80130[add_80180 > 32'h0000_0009 ? 4'h9 : add_80180[3:0]], array_index_80183[literal_80126 > 32'h0000_0009 ? 4'h9 : literal_80126[3:0]]);
  assign add_80190 = array_index_80184[literal_80126 > 32'h0000_0009 ? 4'h9 : literal_80126[3:0]] + smul_80188;
  assign array_update_80192[0] = literal_80126 == 32'h0000_0000 ? add_80190 : array_index_80184[0];
  assign array_update_80192[1] = literal_80126 == 32'h0000_0001 ? add_80190 : array_index_80184[1];
  assign array_update_80192[2] = literal_80126 == 32'h0000_0002 ? add_80190 : array_index_80184[2];
  assign array_update_80192[3] = literal_80126 == 32'h0000_0003 ? add_80190 : array_index_80184[3];
  assign array_update_80192[4] = literal_80126 == 32'h0000_0004 ? add_80190 : array_index_80184[4];
  assign array_update_80192[5] = literal_80126 == 32'h0000_0005 ? add_80190 : array_index_80184[5];
  assign array_update_80192[6] = literal_80126 == 32'h0000_0006 ? add_80190 : array_index_80184[6];
  assign array_update_80192[7] = literal_80126 == 32'h0000_0007 ? add_80190 : array_index_80184[7];
  assign array_update_80192[8] = literal_80126 == 32'h0000_0008 ? add_80190 : array_index_80184[8];
  assign array_update_80192[9] = literal_80126 == 32'h0000_0009 ? add_80190 : array_index_80184[9];
  assign add_80193 = add_80180 + 32'h0000_0001;
  assign array_update_80194[0] = add_80123 == 32'h0000_0000 ? array_update_80192 : array_update_80181[0];
  assign array_update_80194[1] = add_80123 == 32'h0000_0001 ? array_update_80192 : array_update_80181[1];
  assign array_update_80194[2] = add_80123 == 32'h0000_0002 ? array_update_80192 : array_update_80181[2];
  assign array_update_80194[3] = add_80123 == 32'h0000_0003 ? array_update_80192 : array_update_80181[3];
  assign array_update_80194[4] = add_80123 == 32'h0000_0004 ? array_update_80192 : array_update_80181[4];
  assign array_update_80194[5] = add_80123 == 32'h0000_0005 ? array_update_80192 : array_update_80181[5];
  assign array_update_80194[6] = add_80123 == 32'h0000_0006 ? array_update_80192 : array_update_80181[6];
  assign array_update_80194[7] = add_80123 == 32'h0000_0007 ? array_update_80192 : array_update_80181[7];
  assign array_update_80194[8] = add_80123 == 32'h0000_0008 ? array_update_80192 : array_update_80181[8];
  assign array_update_80194[9] = add_80123 == 32'h0000_0009 ? array_update_80192 : array_update_80181[9];
  assign array_index_80196 = array_update_72021[add_80193 > 32'h0000_0009 ? 4'h9 : add_80193[3:0]];
  assign array_index_80197 = array_update_80194[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_80201 = smul32b_32b_x_32b(array_index_80130[add_80193 > 32'h0000_0009 ? 4'h9 : add_80193[3:0]], array_index_80196[literal_80126 > 32'h0000_0009 ? 4'h9 : literal_80126[3:0]]);
  assign add_80203 = array_index_80197[literal_80126 > 32'h0000_0009 ? 4'h9 : literal_80126[3:0]] + smul_80201;
  assign array_update_80205[0] = literal_80126 == 32'h0000_0000 ? add_80203 : array_index_80197[0];
  assign array_update_80205[1] = literal_80126 == 32'h0000_0001 ? add_80203 : array_index_80197[1];
  assign array_update_80205[2] = literal_80126 == 32'h0000_0002 ? add_80203 : array_index_80197[2];
  assign array_update_80205[3] = literal_80126 == 32'h0000_0003 ? add_80203 : array_index_80197[3];
  assign array_update_80205[4] = literal_80126 == 32'h0000_0004 ? add_80203 : array_index_80197[4];
  assign array_update_80205[5] = literal_80126 == 32'h0000_0005 ? add_80203 : array_index_80197[5];
  assign array_update_80205[6] = literal_80126 == 32'h0000_0006 ? add_80203 : array_index_80197[6];
  assign array_update_80205[7] = literal_80126 == 32'h0000_0007 ? add_80203 : array_index_80197[7];
  assign array_update_80205[8] = literal_80126 == 32'h0000_0008 ? add_80203 : array_index_80197[8];
  assign array_update_80205[9] = literal_80126 == 32'h0000_0009 ? add_80203 : array_index_80197[9];
  assign add_80206 = add_80193 + 32'h0000_0001;
  assign array_update_80207[0] = add_80123 == 32'h0000_0000 ? array_update_80205 : array_update_80194[0];
  assign array_update_80207[1] = add_80123 == 32'h0000_0001 ? array_update_80205 : array_update_80194[1];
  assign array_update_80207[2] = add_80123 == 32'h0000_0002 ? array_update_80205 : array_update_80194[2];
  assign array_update_80207[3] = add_80123 == 32'h0000_0003 ? array_update_80205 : array_update_80194[3];
  assign array_update_80207[4] = add_80123 == 32'h0000_0004 ? array_update_80205 : array_update_80194[4];
  assign array_update_80207[5] = add_80123 == 32'h0000_0005 ? array_update_80205 : array_update_80194[5];
  assign array_update_80207[6] = add_80123 == 32'h0000_0006 ? array_update_80205 : array_update_80194[6];
  assign array_update_80207[7] = add_80123 == 32'h0000_0007 ? array_update_80205 : array_update_80194[7];
  assign array_update_80207[8] = add_80123 == 32'h0000_0008 ? array_update_80205 : array_update_80194[8];
  assign array_update_80207[9] = add_80123 == 32'h0000_0009 ? array_update_80205 : array_update_80194[9];
  assign array_index_80209 = array_update_72021[add_80206 > 32'h0000_0009 ? 4'h9 : add_80206[3:0]];
  assign array_index_80210 = array_update_80207[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_80214 = smul32b_32b_x_32b(array_index_80130[add_80206 > 32'h0000_0009 ? 4'h9 : add_80206[3:0]], array_index_80209[literal_80126 > 32'h0000_0009 ? 4'h9 : literal_80126[3:0]]);
  assign add_80216 = array_index_80210[literal_80126 > 32'h0000_0009 ? 4'h9 : literal_80126[3:0]] + smul_80214;
  assign array_update_80218[0] = literal_80126 == 32'h0000_0000 ? add_80216 : array_index_80210[0];
  assign array_update_80218[1] = literal_80126 == 32'h0000_0001 ? add_80216 : array_index_80210[1];
  assign array_update_80218[2] = literal_80126 == 32'h0000_0002 ? add_80216 : array_index_80210[2];
  assign array_update_80218[3] = literal_80126 == 32'h0000_0003 ? add_80216 : array_index_80210[3];
  assign array_update_80218[4] = literal_80126 == 32'h0000_0004 ? add_80216 : array_index_80210[4];
  assign array_update_80218[5] = literal_80126 == 32'h0000_0005 ? add_80216 : array_index_80210[5];
  assign array_update_80218[6] = literal_80126 == 32'h0000_0006 ? add_80216 : array_index_80210[6];
  assign array_update_80218[7] = literal_80126 == 32'h0000_0007 ? add_80216 : array_index_80210[7];
  assign array_update_80218[8] = literal_80126 == 32'h0000_0008 ? add_80216 : array_index_80210[8];
  assign array_update_80218[9] = literal_80126 == 32'h0000_0009 ? add_80216 : array_index_80210[9];
  assign add_80219 = add_80206 + 32'h0000_0001;
  assign array_update_80220[0] = add_80123 == 32'h0000_0000 ? array_update_80218 : array_update_80207[0];
  assign array_update_80220[1] = add_80123 == 32'h0000_0001 ? array_update_80218 : array_update_80207[1];
  assign array_update_80220[2] = add_80123 == 32'h0000_0002 ? array_update_80218 : array_update_80207[2];
  assign array_update_80220[3] = add_80123 == 32'h0000_0003 ? array_update_80218 : array_update_80207[3];
  assign array_update_80220[4] = add_80123 == 32'h0000_0004 ? array_update_80218 : array_update_80207[4];
  assign array_update_80220[5] = add_80123 == 32'h0000_0005 ? array_update_80218 : array_update_80207[5];
  assign array_update_80220[6] = add_80123 == 32'h0000_0006 ? array_update_80218 : array_update_80207[6];
  assign array_update_80220[7] = add_80123 == 32'h0000_0007 ? array_update_80218 : array_update_80207[7];
  assign array_update_80220[8] = add_80123 == 32'h0000_0008 ? array_update_80218 : array_update_80207[8];
  assign array_update_80220[9] = add_80123 == 32'h0000_0009 ? array_update_80218 : array_update_80207[9];
  assign array_index_80222 = array_update_72021[add_80219 > 32'h0000_0009 ? 4'h9 : add_80219[3:0]];
  assign array_index_80223 = array_update_80220[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_80227 = smul32b_32b_x_32b(array_index_80130[add_80219 > 32'h0000_0009 ? 4'h9 : add_80219[3:0]], array_index_80222[literal_80126 > 32'h0000_0009 ? 4'h9 : literal_80126[3:0]]);
  assign add_80229 = array_index_80223[literal_80126 > 32'h0000_0009 ? 4'h9 : literal_80126[3:0]] + smul_80227;
  assign array_update_80231[0] = literal_80126 == 32'h0000_0000 ? add_80229 : array_index_80223[0];
  assign array_update_80231[1] = literal_80126 == 32'h0000_0001 ? add_80229 : array_index_80223[1];
  assign array_update_80231[2] = literal_80126 == 32'h0000_0002 ? add_80229 : array_index_80223[2];
  assign array_update_80231[3] = literal_80126 == 32'h0000_0003 ? add_80229 : array_index_80223[3];
  assign array_update_80231[4] = literal_80126 == 32'h0000_0004 ? add_80229 : array_index_80223[4];
  assign array_update_80231[5] = literal_80126 == 32'h0000_0005 ? add_80229 : array_index_80223[5];
  assign array_update_80231[6] = literal_80126 == 32'h0000_0006 ? add_80229 : array_index_80223[6];
  assign array_update_80231[7] = literal_80126 == 32'h0000_0007 ? add_80229 : array_index_80223[7];
  assign array_update_80231[8] = literal_80126 == 32'h0000_0008 ? add_80229 : array_index_80223[8];
  assign array_update_80231[9] = literal_80126 == 32'h0000_0009 ? add_80229 : array_index_80223[9];
  assign add_80232 = add_80219 + 32'h0000_0001;
  assign array_update_80233[0] = add_80123 == 32'h0000_0000 ? array_update_80231 : array_update_80220[0];
  assign array_update_80233[1] = add_80123 == 32'h0000_0001 ? array_update_80231 : array_update_80220[1];
  assign array_update_80233[2] = add_80123 == 32'h0000_0002 ? array_update_80231 : array_update_80220[2];
  assign array_update_80233[3] = add_80123 == 32'h0000_0003 ? array_update_80231 : array_update_80220[3];
  assign array_update_80233[4] = add_80123 == 32'h0000_0004 ? array_update_80231 : array_update_80220[4];
  assign array_update_80233[5] = add_80123 == 32'h0000_0005 ? array_update_80231 : array_update_80220[5];
  assign array_update_80233[6] = add_80123 == 32'h0000_0006 ? array_update_80231 : array_update_80220[6];
  assign array_update_80233[7] = add_80123 == 32'h0000_0007 ? array_update_80231 : array_update_80220[7];
  assign array_update_80233[8] = add_80123 == 32'h0000_0008 ? array_update_80231 : array_update_80220[8];
  assign array_update_80233[9] = add_80123 == 32'h0000_0009 ? array_update_80231 : array_update_80220[9];
  assign array_index_80235 = array_update_72021[add_80232 > 32'h0000_0009 ? 4'h9 : add_80232[3:0]];
  assign array_index_80236 = array_update_80233[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_80240 = smul32b_32b_x_32b(array_index_80130[add_80232 > 32'h0000_0009 ? 4'h9 : add_80232[3:0]], array_index_80235[literal_80126 > 32'h0000_0009 ? 4'h9 : literal_80126[3:0]]);
  assign add_80242 = array_index_80236[literal_80126 > 32'h0000_0009 ? 4'h9 : literal_80126[3:0]] + smul_80240;
  assign array_update_80244[0] = literal_80126 == 32'h0000_0000 ? add_80242 : array_index_80236[0];
  assign array_update_80244[1] = literal_80126 == 32'h0000_0001 ? add_80242 : array_index_80236[1];
  assign array_update_80244[2] = literal_80126 == 32'h0000_0002 ? add_80242 : array_index_80236[2];
  assign array_update_80244[3] = literal_80126 == 32'h0000_0003 ? add_80242 : array_index_80236[3];
  assign array_update_80244[4] = literal_80126 == 32'h0000_0004 ? add_80242 : array_index_80236[4];
  assign array_update_80244[5] = literal_80126 == 32'h0000_0005 ? add_80242 : array_index_80236[5];
  assign array_update_80244[6] = literal_80126 == 32'h0000_0006 ? add_80242 : array_index_80236[6];
  assign array_update_80244[7] = literal_80126 == 32'h0000_0007 ? add_80242 : array_index_80236[7];
  assign array_update_80244[8] = literal_80126 == 32'h0000_0008 ? add_80242 : array_index_80236[8];
  assign array_update_80244[9] = literal_80126 == 32'h0000_0009 ? add_80242 : array_index_80236[9];
  assign add_80245 = add_80232 + 32'h0000_0001;
  assign array_update_80246[0] = add_80123 == 32'h0000_0000 ? array_update_80244 : array_update_80233[0];
  assign array_update_80246[1] = add_80123 == 32'h0000_0001 ? array_update_80244 : array_update_80233[1];
  assign array_update_80246[2] = add_80123 == 32'h0000_0002 ? array_update_80244 : array_update_80233[2];
  assign array_update_80246[3] = add_80123 == 32'h0000_0003 ? array_update_80244 : array_update_80233[3];
  assign array_update_80246[4] = add_80123 == 32'h0000_0004 ? array_update_80244 : array_update_80233[4];
  assign array_update_80246[5] = add_80123 == 32'h0000_0005 ? array_update_80244 : array_update_80233[5];
  assign array_update_80246[6] = add_80123 == 32'h0000_0006 ? array_update_80244 : array_update_80233[6];
  assign array_update_80246[7] = add_80123 == 32'h0000_0007 ? array_update_80244 : array_update_80233[7];
  assign array_update_80246[8] = add_80123 == 32'h0000_0008 ? array_update_80244 : array_update_80233[8];
  assign array_update_80246[9] = add_80123 == 32'h0000_0009 ? array_update_80244 : array_update_80233[9];
  assign array_index_80248 = array_update_72021[add_80245 > 32'h0000_0009 ? 4'h9 : add_80245[3:0]];
  assign array_index_80249 = array_update_80246[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_80253 = smul32b_32b_x_32b(array_index_80130[add_80245 > 32'h0000_0009 ? 4'h9 : add_80245[3:0]], array_index_80248[literal_80126 > 32'h0000_0009 ? 4'h9 : literal_80126[3:0]]);
  assign add_80255 = array_index_80249[literal_80126 > 32'h0000_0009 ? 4'h9 : literal_80126[3:0]] + smul_80253;
  assign array_update_80256[0] = literal_80126 == 32'h0000_0000 ? add_80255 : array_index_80249[0];
  assign array_update_80256[1] = literal_80126 == 32'h0000_0001 ? add_80255 : array_index_80249[1];
  assign array_update_80256[2] = literal_80126 == 32'h0000_0002 ? add_80255 : array_index_80249[2];
  assign array_update_80256[3] = literal_80126 == 32'h0000_0003 ? add_80255 : array_index_80249[3];
  assign array_update_80256[4] = literal_80126 == 32'h0000_0004 ? add_80255 : array_index_80249[4];
  assign array_update_80256[5] = literal_80126 == 32'h0000_0005 ? add_80255 : array_index_80249[5];
  assign array_update_80256[6] = literal_80126 == 32'h0000_0006 ? add_80255 : array_index_80249[6];
  assign array_update_80256[7] = literal_80126 == 32'h0000_0007 ? add_80255 : array_index_80249[7];
  assign array_update_80256[8] = literal_80126 == 32'h0000_0008 ? add_80255 : array_index_80249[8];
  assign array_update_80256[9] = literal_80126 == 32'h0000_0009 ? add_80255 : array_index_80249[9];
  assign array_update_80257[0] = add_80123 == 32'h0000_0000 ? array_update_80256 : array_update_80246[0];
  assign array_update_80257[1] = add_80123 == 32'h0000_0001 ? array_update_80256 : array_update_80246[1];
  assign array_update_80257[2] = add_80123 == 32'h0000_0002 ? array_update_80256 : array_update_80246[2];
  assign array_update_80257[3] = add_80123 == 32'h0000_0003 ? array_update_80256 : array_update_80246[3];
  assign array_update_80257[4] = add_80123 == 32'h0000_0004 ? array_update_80256 : array_update_80246[4];
  assign array_update_80257[5] = add_80123 == 32'h0000_0005 ? array_update_80256 : array_update_80246[5];
  assign array_update_80257[6] = add_80123 == 32'h0000_0006 ? array_update_80256 : array_update_80246[6];
  assign array_update_80257[7] = add_80123 == 32'h0000_0007 ? array_update_80256 : array_update_80246[7];
  assign array_update_80257[8] = add_80123 == 32'h0000_0008 ? array_update_80256 : array_update_80246[8];
  assign array_update_80257[9] = add_80123 == 32'h0000_0009 ? array_update_80256 : array_update_80246[9];
  assign array_index_80259 = array_update_80257[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign add_80261 = literal_80126 + 32'h0000_0001;
  assign array_update_80262[0] = add_80261 == 32'h0000_0000 ? 32'h0000_0000 : array_index_80259[0];
  assign array_update_80262[1] = add_80261 == 32'h0000_0001 ? 32'h0000_0000 : array_index_80259[1];
  assign array_update_80262[2] = add_80261 == 32'h0000_0002 ? 32'h0000_0000 : array_index_80259[2];
  assign array_update_80262[3] = add_80261 == 32'h0000_0003 ? 32'h0000_0000 : array_index_80259[3];
  assign array_update_80262[4] = add_80261 == 32'h0000_0004 ? 32'h0000_0000 : array_index_80259[4];
  assign array_update_80262[5] = add_80261 == 32'h0000_0005 ? 32'h0000_0000 : array_index_80259[5];
  assign array_update_80262[6] = add_80261 == 32'h0000_0006 ? 32'h0000_0000 : array_index_80259[6];
  assign array_update_80262[7] = add_80261 == 32'h0000_0007 ? 32'h0000_0000 : array_index_80259[7];
  assign array_update_80262[8] = add_80261 == 32'h0000_0008 ? 32'h0000_0000 : array_index_80259[8];
  assign array_update_80262[9] = add_80261 == 32'h0000_0009 ? 32'h0000_0000 : array_index_80259[9];
  assign literal_80263 = 32'h0000_0000;
  assign array_update_80264[0] = add_80123 == 32'h0000_0000 ? array_update_80262 : array_update_80257[0];
  assign array_update_80264[1] = add_80123 == 32'h0000_0001 ? array_update_80262 : array_update_80257[1];
  assign array_update_80264[2] = add_80123 == 32'h0000_0002 ? array_update_80262 : array_update_80257[2];
  assign array_update_80264[3] = add_80123 == 32'h0000_0003 ? array_update_80262 : array_update_80257[3];
  assign array_update_80264[4] = add_80123 == 32'h0000_0004 ? array_update_80262 : array_update_80257[4];
  assign array_update_80264[5] = add_80123 == 32'h0000_0005 ? array_update_80262 : array_update_80257[5];
  assign array_update_80264[6] = add_80123 == 32'h0000_0006 ? array_update_80262 : array_update_80257[6];
  assign array_update_80264[7] = add_80123 == 32'h0000_0007 ? array_update_80262 : array_update_80257[7];
  assign array_update_80264[8] = add_80123 == 32'h0000_0008 ? array_update_80262 : array_update_80257[8];
  assign array_update_80264[9] = add_80123 == 32'h0000_0009 ? array_update_80262 : array_update_80257[9];
  assign array_index_80266 = array_update_72021[literal_80263 > 32'h0000_0009 ? 4'h9 : literal_80263[3:0]];
  assign array_index_80267 = array_update_80264[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_80271 = smul32b_32b_x_32b(array_index_80130[literal_80263 > 32'h0000_0009 ? 4'h9 : literal_80263[3:0]], array_index_80266[add_80261 > 32'h0000_0009 ? 4'h9 : add_80261[3:0]]);
  assign add_80273 = array_index_80267[add_80261 > 32'h0000_0009 ? 4'h9 : add_80261[3:0]] + smul_80271;
  assign array_update_80275[0] = add_80261 == 32'h0000_0000 ? add_80273 : array_index_80267[0];
  assign array_update_80275[1] = add_80261 == 32'h0000_0001 ? add_80273 : array_index_80267[1];
  assign array_update_80275[2] = add_80261 == 32'h0000_0002 ? add_80273 : array_index_80267[2];
  assign array_update_80275[3] = add_80261 == 32'h0000_0003 ? add_80273 : array_index_80267[3];
  assign array_update_80275[4] = add_80261 == 32'h0000_0004 ? add_80273 : array_index_80267[4];
  assign array_update_80275[5] = add_80261 == 32'h0000_0005 ? add_80273 : array_index_80267[5];
  assign array_update_80275[6] = add_80261 == 32'h0000_0006 ? add_80273 : array_index_80267[6];
  assign array_update_80275[7] = add_80261 == 32'h0000_0007 ? add_80273 : array_index_80267[7];
  assign array_update_80275[8] = add_80261 == 32'h0000_0008 ? add_80273 : array_index_80267[8];
  assign array_update_80275[9] = add_80261 == 32'h0000_0009 ? add_80273 : array_index_80267[9];
  assign add_80276 = literal_80263 + 32'h0000_0001;
  assign array_update_80277[0] = add_80123 == 32'h0000_0000 ? array_update_80275 : array_update_80264[0];
  assign array_update_80277[1] = add_80123 == 32'h0000_0001 ? array_update_80275 : array_update_80264[1];
  assign array_update_80277[2] = add_80123 == 32'h0000_0002 ? array_update_80275 : array_update_80264[2];
  assign array_update_80277[3] = add_80123 == 32'h0000_0003 ? array_update_80275 : array_update_80264[3];
  assign array_update_80277[4] = add_80123 == 32'h0000_0004 ? array_update_80275 : array_update_80264[4];
  assign array_update_80277[5] = add_80123 == 32'h0000_0005 ? array_update_80275 : array_update_80264[5];
  assign array_update_80277[6] = add_80123 == 32'h0000_0006 ? array_update_80275 : array_update_80264[6];
  assign array_update_80277[7] = add_80123 == 32'h0000_0007 ? array_update_80275 : array_update_80264[7];
  assign array_update_80277[8] = add_80123 == 32'h0000_0008 ? array_update_80275 : array_update_80264[8];
  assign array_update_80277[9] = add_80123 == 32'h0000_0009 ? array_update_80275 : array_update_80264[9];
  assign array_index_80279 = array_update_72021[add_80276 > 32'h0000_0009 ? 4'h9 : add_80276[3:0]];
  assign array_index_80280 = array_update_80277[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_80284 = smul32b_32b_x_32b(array_index_80130[add_80276 > 32'h0000_0009 ? 4'h9 : add_80276[3:0]], array_index_80279[add_80261 > 32'h0000_0009 ? 4'h9 : add_80261[3:0]]);
  assign add_80286 = array_index_80280[add_80261 > 32'h0000_0009 ? 4'h9 : add_80261[3:0]] + smul_80284;
  assign array_update_80288[0] = add_80261 == 32'h0000_0000 ? add_80286 : array_index_80280[0];
  assign array_update_80288[1] = add_80261 == 32'h0000_0001 ? add_80286 : array_index_80280[1];
  assign array_update_80288[2] = add_80261 == 32'h0000_0002 ? add_80286 : array_index_80280[2];
  assign array_update_80288[3] = add_80261 == 32'h0000_0003 ? add_80286 : array_index_80280[3];
  assign array_update_80288[4] = add_80261 == 32'h0000_0004 ? add_80286 : array_index_80280[4];
  assign array_update_80288[5] = add_80261 == 32'h0000_0005 ? add_80286 : array_index_80280[5];
  assign array_update_80288[6] = add_80261 == 32'h0000_0006 ? add_80286 : array_index_80280[6];
  assign array_update_80288[7] = add_80261 == 32'h0000_0007 ? add_80286 : array_index_80280[7];
  assign array_update_80288[8] = add_80261 == 32'h0000_0008 ? add_80286 : array_index_80280[8];
  assign array_update_80288[9] = add_80261 == 32'h0000_0009 ? add_80286 : array_index_80280[9];
  assign add_80289 = add_80276 + 32'h0000_0001;
  assign array_update_80290[0] = add_80123 == 32'h0000_0000 ? array_update_80288 : array_update_80277[0];
  assign array_update_80290[1] = add_80123 == 32'h0000_0001 ? array_update_80288 : array_update_80277[1];
  assign array_update_80290[2] = add_80123 == 32'h0000_0002 ? array_update_80288 : array_update_80277[2];
  assign array_update_80290[3] = add_80123 == 32'h0000_0003 ? array_update_80288 : array_update_80277[3];
  assign array_update_80290[4] = add_80123 == 32'h0000_0004 ? array_update_80288 : array_update_80277[4];
  assign array_update_80290[5] = add_80123 == 32'h0000_0005 ? array_update_80288 : array_update_80277[5];
  assign array_update_80290[6] = add_80123 == 32'h0000_0006 ? array_update_80288 : array_update_80277[6];
  assign array_update_80290[7] = add_80123 == 32'h0000_0007 ? array_update_80288 : array_update_80277[7];
  assign array_update_80290[8] = add_80123 == 32'h0000_0008 ? array_update_80288 : array_update_80277[8];
  assign array_update_80290[9] = add_80123 == 32'h0000_0009 ? array_update_80288 : array_update_80277[9];
  assign array_index_80292 = array_update_72021[add_80289 > 32'h0000_0009 ? 4'h9 : add_80289[3:0]];
  assign array_index_80293 = array_update_80290[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_80297 = smul32b_32b_x_32b(array_index_80130[add_80289 > 32'h0000_0009 ? 4'h9 : add_80289[3:0]], array_index_80292[add_80261 > 32'h0000_0009 ? 4'h9 : add_80261[3:0]]);
  assign add_80299 = array_index_80293[add_80261 > 32'h0000_0009 ? 4'h9 : add_80261[3:0]] + smul_80297;
  assign array_update_80301[0] = add_80261 == 32'h0000_0000 ? add_80299 : array_index_80293[0];
  assign array_update_80301[1] = add_80261 == 32'h0000_0001 ? add_80299 : array_index_80293[1];
  assign array_update_80301[2] = add_80261 == 32'h0000_0002 ? add_80299 : array_index_80293[2];
  assign array_update_80301[3] = add_80261 == 32'h0000_0003 ? add_80299 : array_index_80293[3];
  assign array_update_80301[4] = add_80261 == 32'h0000_0004 ? add_80299 : array_index_80293[4];
  assign array_update_80301[5] = add_80261 == 32'h0000_0005 ? add_80299 : array_index_80293[5];
  assign array_update_80301[6] = add_80261 == 32'h0000_0006 ? add_80299 : array_index_80293[6];
  assign array_update_80301[7] = add_80261 == 32'h0000_0007 ? add_80299 : array_index_80293[7];
  assign array_update_80301[8] = add_80261 == 32'h0000_0008 ? add_80299 : array_index_80293[8];
  assign array_update_80301[9] = add_80261 == 32'h0000_0009 ? add_80299 : array_index_80293[9];
  assign add_80302 = add_80289 + 32'h0000_0001;
  assign array_update_80303[0] = add_80123 == 32'h0000_0000 ? array_update_80301 : array_update_80290[0];
  assign array_update_80303[1] = add_80123 == 32'h0000_0001 ? array_update_80301 : array_update_80290[1];
  assign array_update_80303[2] = add_80123 == 32'h0000_0002 ? array_update_80301 : array_update_80290[2];
  assign array_update_80303[3] = add_80123 == 32'h0000_0003 ? array_update_80301 : array_update_80290[3];
  assign array_update_80303[4] = add_80123 == 32'h0000_0004 ? array_update_80301 : array_update_80290[4];
  assign array_update_80303[5] = add_80123 == 32'h0000_0005 ? array_update_80301 : array_update_80290[5];
  assign array_update_80303[6] = add_80123 == 32'h0000_0006 ? array_update_80301 : array_update_80290[6];
  assign array_update_80303[7] = add_80123 == 32'h0000_0007 ? array_update_80301 : array_update_80290[7];
  assign array_update_80303[8] = add_80123 == 32'h0000_0008 ? array_update_80301 : array_update_80290[8];
  assign array_update_80303[9] = add_80123 == 32'h0000_0009 ? array_update_80301 : array_update_80290[9];
  assign array_index_80305 = array_update_72021[add_80302 > 32'h0000_0009 ? 4'h9 : add_80302[3:0]];
  assign array_index_80306 = array_update_80303[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_80310 = smul32b_32b_x_32b(array_index_80130[add_80302 > 32'h0000_0009 ? 4'h9 : add_80302[3:0]], array_index_80305[add_80261 > 32'h0000_0009 ? 4'h9 : add_80261[3:0]]);
  assign add_80312 = array_index_80306[add_80261 > 32'h0000_0009 ? 4'h9 : add_80261[3:0]] + smul_80310;
  assign array_update_80314[0] = add_80261 == 32'h0000_0000 ? add_80312 : array_index_80306[0];
  assign array_update_80314[1] = add_80261 == 32'h0000_0001 ? add_80312 : array_index_80306[1];
  assign array_update_80314[2] = add_80261 == 32'h0000_0002 ? add_80312 : array_index_80306[2];
  assign array_update_80314[3] = add_80261 == 32'h0000_0003 ? add_80312 : array_index_80306[3];
  assign array_update_80314[4] = add_80261 == 32'h0000_0004 ? add_80312 : array_index_80306[4];
  assign array_update_80314[5] = add_80261 == 32'h0000_0005 ? add_80312 : array_index_80306[5];
  assign array_update_80314[6] = add_80261 == 32'h0000_0006 ? add_80312 : array_index_80306[6];
  assign array_update_80314[7] = add_80261 == 32'h0000_0007 ? add_80312 : array_index_80306[7];
  assign array_update_80314[8] = add_80261 == 32'h0000_0008 ? add_80312 : array_index_80306[8];
  assign array_update_80314[9] = add_80261 == 32'h0000_0009 ? add_80312 : array_index_80306[9];
  assign add_80315 = add_80302 + 32'h0000_0001;
  assign array_update_80316[0] = add_80123 == 32'h0000_0000 ? array_update_80314 : array_update_80303[0];
  assign array_update_80316[1] = add_80123 == 32'h0000_0001 ? array_update_80314 : array_update_80303[1];
  assign array_update_80316[2] = add_80123 == 32'h0000_0002 ? array_update_80314 : array_update_80303[2];
  assign array_update_80316[3] = add_80123 == 32'h0000_0003 ? array_update_80314 : array_update_80303[3];
  assign array_update_80316[4] = add_80123 == 32'h0000_0004 ? array_update_80314 : array_update_80303[4];
  assign array_update_80316[5] = add_80123 == 32'h0000_0005 ? array_update_80314 : array_update_80303[5];
  assign array_update_80316[6] = add_80123 == 32'h0000_0006 ? array_update_80314 : array_update_80303[6];
  assign array_update_80316[7] = add_80123 == 32'h0000_0007 ? array_update_80314 : array_update_80303[7];
  assign array_update_80316[8] = add_80123 == 32'h0000_0008 ? array_update_80314 : array_update_80303[8];
  assign array_update_80316[9] = add_80123 == 32'h0000_0009 ? array_update_80314 : array_update_80303[9];
  assign array_index_80318 = array_update_72021[add_80315 > 32'h0000_0009 ? 4'h9 : add_80315[3:0]];
  assign array_index_80319 = array_update_80316[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_80323 = smul32b_32b_x_32b(array_index_80130[add_80315 > 32'h0000_0009 ? 4'h9 : add_80315[3:0]], array_index_80318[add_80261 > 32'h0000_0009 ? 4'h9 : add_80261[3:0]]);
  assign add_80325 = array_index_80319[add_80261 > 32'h0000_0009 ? 4'h9 : add_80261[3:0]] + smul_80323;
  assign array_update_80327[0] = add_80261 == 32'h0000_0000 ? add_80325 : array_index_80319[0];
  assign array_update_80327[1] = add_80261 == 32'h0000_0001 ? add_80325 : array_index_80319[1];
  assign array_update_80327[2] = add_80261 == 32'h0000_0002 ? add_80325 : array_index_80319[2];
  assign array_update_80327[3] = add_80261 == 32'h0000_0003 ? add_80325 : array_index_80319[3];
  assign array_update_80327[4] = add_80261 == 32'h0000_0004 ? add_80325 : array_index_80319[4];
  assign array_update_80327[5] = add_80261 == 32'h0000_0005 ? add_80325 : array_index_80319[5];
  assign array_update_80327[6] = add_80261 == 32'h0000_0006 ? add_80325 : array_index_80319[6];
  assign array_update_80327[7] = add_80261 == 32'h0000_0007 ? add_80325 : array_index_80319[7];
  assign array_update_80327[8] = add_80261 == 32'h0000_0008 ? add_80325 : array_index_80319[8];
  assign array_update_80327[9] = add_80261 == 32'h0000_0009 ? add_80325 : array_index_80319[9];
  assign add_80328 = add_80315 + 32'h0000_0001;
  assign array_update_80329[0] = add_80123 == 32'h0000_0000 ? array_update_80327 : array_update_80316[0];
  assign array_update_80329[1] = add_80123 == 32'h0000_0001 ? array_update_80327 : array_update_80316[1];
  assign array_update_80329[2] = add_80123 == 32'h0000_0002 ? array_update_80327 : array_update_80316[2];
  assign array_update_80329[3] = add_80123 == 32'h0000_0003 ? array_update_80327 : array_update_80316[3];
  assign array_update_80329[4] = add_80123 == 32'h0000_0004 ? array_update_80327 : array_update_80316[4];
  assign array_update_80329[5] = add_80123 == 32'h0000_0005 ? array_update_80327 : array_update_80316[5];
  assign array_update_80329[6] = add_80123 == 32'h0000_0006 ? array_update_80327 : array_update_80316[6];
  assign array_update_80329[7] = add_80123 == 32'h0000_0007 ? array_update_80327 : array_update_80316[7];
  assign array_update_80329[8] = add_80123 == 32'h0000_0008 ? array_update_80327 : array_update_80316[8];
  assign array_update_80329[9] = add_80123 == 32'h0000_0009 ? array_update_80327 : array_update_80316[9];
  assign array_index_80331 = array_update_72021[add_80328 > 32'h0000_0009 ? 4'h9 : add_80328[3:0]];
  assign array_index_80332 = array_update_80329[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_80336 = smul32b_32b_x_32b(array_index_80130[add_80328 > 32'h0000_0009 ? 4'h9 : add_80328[3:0]], array_index_80331[add_80261 > 32'h0000_0009 ? 4'h9 : add_80261[3:0]]);
  assign add_80338 = array_index_80332[add_80261 > 32'h0000_0009 ? 4'h9 : add_80261[3:0]] + smul_80336;
  assign array_update_80340[0] = add_80261 == 32'h0000_0000 ? add_80338 : array_index_80332[0];
  assign array_update_80340[1] = add_80261 == 32'h0000_0001 ? add_80338 : array_index_80332[1];
  assign array_update_80340[2] = add_80261 == 32'h0000_0002 ? add_80338 : array_index_80332[2];
  assign array_update_80340[3] = add_80261 == 32'h0000_0003 ? add_80338 : array_index_80332[3];
  assign array_update_80340[4] = add_80261 == 32'h0000_0004 ? add_80338 : array_index_80332[4];
  assign array_update_80340[5] = add_80261 == 32'h0000_0005 ? add_80338 : array_index_80332[5];
  assign array_update_80340[6] = add_80261 == 32'h0000_0006 ? add_80338 : array_index_80332[6];
  assign array_update_80340[7] = add_80261 == 32'h0000_0007 ? add_80338 : array_index_80332[7];
  assign array_update_80340[8] = add_80261 == 32'h0000_0008 ? add_80338 : array_index_80332[8];
  assign array_update_80340[9] = add_80261 == 32'h0000_0009 ? add_80338 : array_index_80332[9];
  assign add_80341 = add_80328 + 32'h0000_0001;
  assign array_update_80342[0] = add_80123 == 32'h0000_0000 ? array_update_80340 : array_update_80329[0];
  assign array_update_80342[1] = add_80123 == 32'h0000_0001 ? array_update_80340 : array_update_80329[1];
  assign array_update_80342[2] = add_80123 == 32'h0000_0002 ? array_update_80340 : array_update_80329[2];
  assign array_update_80342[3] = add_80123 == 32'h0000_0003 ? array_update_80340 : array_update_80329[3];
  assign array_update_80342[4] = add_80123 == 32'h0000_0004 ? array_update_80340 : array_update_80329[4];
  assign array_update_80342[5] = add_80123 == 32'h0000_0005 ? array_update_80340 : array_update_80329[5];
  assign array_update_80342[6] = add_80123 == 32'h0000_0006 ? array_update_80340 : array_update_80329[6];
  assign array_update_80342[7] = add_80123 == 32'h0000_0007 ? array_update_80340 : array_update_80329[7];
  assign array_update_80342[8] = add_80123 == 32'h0000_0008 ? array_update_80340 : array_update_80329[8];
  assign array_update_80342[9] = add_80123 == 32'h0000_0009 ? array_update_80340 : array_update_80329[9];
  assign array_index_80344 = array_update_72021[add_80341 > 32'h0000_0009 ? 4'h9 : add_80341[3:0]];
  assign array_index_80345 = array_update_80342[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_80349 = smul32b_32b_x_32b(array_index_80130[add_80341 > 32'h0000_0009 ? 4'h9 : add_80341[3:0]], array_index_80344[add_80261 > 32'h0000_0009 ? 4'h9 : add_80261[3:0]]);
  assign add_80351 = array_index_80345[add_80261 > 32'h0000_0009 ? 4'h9 : add_80261[3:0]] + smul_80349;
  assign array_update_80353[0] = add_80261 == 32'h0000_0000 ? add_80351 : array_index_80345[0];
  assign array_update_80353[1] = add_80261 == 32'h0000_0001 ? add_80351 : array_index_80345[1];
  assign array_update_80353[2] = add_80261 == 32'h0000_0002 ? add_80351 : array_index_80345[2];
  assign array_update_80353[3] = add_80261 == 32'h0000_0003 ? add_80351 : array_index_80345[3];
  assign array_update_80353[4] = add_80261 == 32'h0000_0004 ? add_80351 : array_index_80345[4];
  assign array_update_80353[5] = add_80261 == 32'h0000_0005 ? add_80351 : array_index_80345[5];
  assign array_update_80353[6] = add_80261 == 32'h0000_0006 ? add_80351 : array_index_80345[6];
  assign array_update_80353[7] = add_80261 == 32'h0000_0007 ? add_80351 : array_index_80345[7];
  assign array_update_80353[8] = add_80261 == 32'h0000_0008 ? add_80351 : array_index_80345[8];
  assign array_update_80353[9] = add_80261 == 32'h0000_0009 ? add_80351 : array_index_80345[9];
  assign add_80354 = add_80341 + 32'h0000_0001;
  assign array_update_80355[0] = add_80123 == 32'h0000_0000 ? array_update_80353 : array_update_80342[0];
  assign array_update_80355[1] = add_80123 == 32'h0000_0001 ? array_update_80353 : array_update_80342[1];
  assign array_update_80355[2] = add_80123 == 32'h0000_0002 ? array_update_80353 : array_update_80342[2];
  assign array_update_80355[3] = add_80123 == 32'h0000_0003 ? array_update_80353 : array_update_80342[3];
  assign array_update_80355[4] = add_80123 == 32'h0000_0004 ? array_update_80353 : array_update_80342[4];
  assign array_update_80355[5] = add_80123 == 32'h0000_0005 ? array_update_80353 : array_update_80342[5];
  assign array_update_80355[6] = add_80123 == 32'h0000_0006 ? array_update_80353 : array_update_80342[6];
  assign array_update_80355[7] = add_80123 == 32'h0000_0007 ? array_update_80353 : array_update_80342[7];
  assign array_update_80355[8] = add_80123 == 32'h0000_0008 ? array_update_80353 : array_update_80342[8];
  assign array_update_80355[9] = add_80123 == 32'h0000_0009 ? array_update_80353 : array_update_80342[9];
  assign array_index_80357 = array_update_72021[add_80354 > 32'h0000_0009 ? 4'h9 : add_80354[3:0]];
  assign array_index_80358 = array_update_80355[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_80362 = smul32b_32b_x_32b(array_index_80130[add_80354 > 32'h0000_0009 ? 4'h9 : add_80354[3:0]], array_index_80357[add_80261 > 32'h0000_0009 ? 4'h9 : add_80261[3:0]]);
  assign add_80364 = array_index_80358[add_80261 > 32'h0000_0009 ? 4'h9 : add_80261[3:0]] + smul_80362;
  assign array_update_80366[0] = add_80261 == 32'h0000_0000 ? add_80364 : array_index_80358[0];
  assign array_update_80366[1] = add_80261 == 32'h0000_0001 ? add_80364 : array_index_80358[1];
  assign array_update_80366[2] = add_80261 == 32'h0000_0002 ? add_80364 : array_index_80358[2];
  assign array_update_80366[3] = add_80261 == 32'h0000_0003 ? add_80364 : array_index_80358[3];
  assign array_update_80366[4] = add_80261 == 32'h0000_0004 ? add_80364 : array_index_80358[4];
  assign array_update_80366[5] = add_80261 == 32'h0000_0005 ? add_80364 : array_index_80358[5];
  assign array_update_80366[6] = add_80261 == 32'h0000_0006 ? add_80364 : array_index_80358[6];
  assign array_update_80366[7] = add_80261 == 32'h0000_0007 ? add_80364 : array_index_80358[7];
  assign array_update_80366[8] = add_80261 == 32'h0000_0008 ? add_80364 : array_index_80358[8];
  assign array_update_80366[9] = add_80261 == 32'h0000_0009 ? add_80364 : array_index_80358[9];
  assign add_80367 = add_80354 + 32'h0000_0001;
  assign array_update_80368[0] = add_80123 == 32'h0000_0000 ? array_update_80366 : array_update_80355[0];
  assign array_update_80368[1] = add_80123 == 32'h0000_0001 ? array_update_80366 : array_update_80355[1];
  assign array_update_80368[2] = add_80123 == 32'h0000_0002 ? array_update_80366 : array_update_80355[2];
  assign array_update_80368[3] = add_80123 == 32'h0000_0003 ? array_update_80366 : array_update_80355[3];
  assign array_update_80368[4] = add_80123 == 32'h0000_0004 ? array_update_80366 : array_update_80355[4];
  assign array_update_80368[5] = add_80123 == 32'h0000_0005 ? array_update_80366 : array_update_80355[5];
  assign array_update_80368[6] = add_80123 == 32'h0000_0006 ? array_update_80366 : array_update_80355[6];
  assign array_update_80368[7] = add_80123 == 32'h0000_0007 ? array_update_80366 : array_update_80355[7];
  assign array_update_80368[8] = add_80123 == 32'h0000_0008 ? array_update_80366 : array_update_80355[8];
  assign array_update_80368[9] = add_80123 == 32'h0000_0009 ? array_update_80366 : array_update_80355[9];
  assign array_index_80370 = array_update_72021[add_80367 > 32'h0000_0009 ? 4'h9 : add_80367[3:0]];
  assign array_index_80371 = array_update_80368[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_80375 = smul32b_32b_x_32b(array_index_80130[add_80367 > 32'h0000_0009 ? 4'h9 : add_80367[3:0]], array_index_80370[add_80261 > 32'h0000_0009 ? 4'h9 : add_80261[3:0]]);
  assign add_80377 = array_index_80371[add_80261 > 32'h0000_0009 ? 4'h9 : add_80261[3:0]] + smul_80375;
  assign array_update_80379[0] = add_80261 == 32'h0000_0000 ? add_80377 : array_index_80371[0];
  assign array_update_80379[1] = add_80261 == 32'h0000_0001 ? add_80377 : array_index_80371[1];
  assign array_update_80379[2] = add_80261 == 32'h0000_0002 ? add_80377 : array_index_80371[2];
  assign array_update_80379[3] = add_80261 == 32'h0000_0003 ? add_80377 : array_index_80371[3];
  assign array_update_80379[4] = add_80261 == 32'h0000_0004 ? add_80377 : array_index_80371[4];
  assign array_update_80379[5] = add_80261 == 32'h0000_0005 ? add_80377 : array_index_80371[5];
  assign array_update_80379[6] = add_80261 == 32'h0000_0006 ? add_80377 : array_index_80371[6];
  assign array_update_80379[7] = add_80261 == 32'h0000_0007 ? add_80377 : array_index_80371[7];
  assign array_update_80379[8] = add_80261 == 32'h0000_0008 ? add_80377 : array_index_80371[8];
  assign array_update_80379[9] = add_80261 == 32'h0000_0009 ? add_80377 : array_index_80371[9];
  assign add_80380 = add_80367 + 32'h0000_0001;
  assign array_update_80381[0] = add_80123 == 32'h0000_0000 ? array_update_80379 : array_update_80368[0];
  assign array_update_80381[1] = add_80123 == 32'h0000_0001 ? array_update_80379 : array_update_80368[1];
  assign array_update_80381[2] = add_80123 == 32'h0000_0002 ? array_update_80379 : array_update_80368[2];
  assign array_update_80381[3] = add_80123 == 32'h0000_0003 ? array_update_80379 : array_update_80368[3];
  assign array_update_80381[4] = add_80123 == 32'h0000_0004 ? array_update_80379 : array_update_80368[4];
  assign array_update_80381[5] = add_80123 == 32'h0000_0005 ? array_update_80379 : array_update_80368[5];
  assign array_update_80381[6] = add_80123 == 32'h0000_0006 ? array_update_80379 : array_update_80368[6];
  assign array_update_80381[7] = add_80123 == 32'h0000_0007 ? array_update_80379 : array_update_80368[7];
  assign array_update_80381[8] = add_80123 == 32'h0000_0008 ? array_update_80379 : array_update_80368[8];
  assign array_update_80381[9] = add_80123 == 32'h0000_0009 ? array_update_80379 : array_update_80368[9];
  assign array_index_80383 = array_update_72021[add_80380 > 32'h0000_0009 ? 4'h9 : add_80380[3:0]];
  assign array_index_80384 = array_update_80381[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_80388 = smul32b_32b_x_32b(array_index_80130[add_80380 > 32'h0000_0009 ? 4'h9 : add_80380[3:0]], array_index_80383[add_80261 > 32'h0000_0009 ? 4'h9 : add_80261[3:0]]);
  assign add_80390 = array_index_80384[add_80261 > 32'h0000_0009 ? 4'h9 : add_80261[3:0]] + smul_80388;
  assign array_update_80391[0] = add_80261 == 32'h0000_0000 ? add_80390 : array_index_80384[0];
  assign array_update_80391[1] = add_80261 == 32'h0000_0001 ? add_80390 : array_index_80384[1];
  assign array_update_80391[2] = add_80261 == 32'h0000_0002 ? add_80390 : array_index_80384[2];
  assign array_update_80391[3] = add_80261 == 32'h0000_0003 ? add_80390 : array_index_80384[3];
  assign array_update_80391[4] = add_80261 == 32'h0000_0004 ? add_80390 : array_index_80384[4];
  assign array_update_80391[5] = add_80261 == 32'h0000_0005 ? add_80390 : array_index_80384[5];
  assign array_update_80391[6] = add_80261 == 32'h0000_0006 ? add_80390 : array_index_80384[6];
  assign array_update_80391[7] = add_80261 == 32'h0000_0007 ? add_80390 : array_index_80384[7];
  assign array_update_80391[8] = add_80261 == 32'h0000_0008 ? add_80390 : array_index_80384[8];
  assign array_update_80391[9] = add_80261 == 32'h0000_0009 ? add_80390 : array_index_80384[9];
  assign array_update_80392[0] = add_80123 == 32'h0000_0000 ? array_update_80391 : array_update_80381[0];
  assign array_update_80392[1] = add_80123 == 32'h0000_0001 ? array_update_80391 : array_update_80381[1];
  assign array_update_80392[2] = add_80123 == 32'h0000_0002 ? array_update_80391 : array_update_80381[2];
  assign array_update_80392[3] = add_80123 == 32'h0000_0003 ? array_update_80391 : array_update_80381[3];
  assign array_update_80392[4] = add_80123 == 32'h0000_0004 ? array_update_80391 : array_update_80381[4];
  assign array_update_80392[5] = add_80123 == 32'h0000_0005 ? array_update_80391 : array_update_80381[5];
  assign array_update_80392[6] = add_80123 == 32'h0000_0006 ? array_update_80391 : array_update_80381[6];
  assign array_update_80392[7] = add_80123 == 32'h0000_0007 ? array_update_80391 : array_update_80381[7];
  assign array_update_80392[8] = add_80123 == 32'h0000_0008 ? array_update_80391 : array_update_80381[8];
  assign array_update_80392[9] = add_80123 == 32'h0000_0009 ? array_update_80391 : array_update_80381[9];
  assign array_index_80394 = array_update_80392[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign add_80396 = add_80261 + 32'h0000_0001;
  assign array_update_80397[0] = add_80396 == 32'h0000_0000 ? 32'h0000_0000 : array_index_80394[0];
  assign array_update_80397[1] = add_80396 == 32'h0000_0001 ? 32'h0000_0000 : array_index_80394[1];
  assign array_update_80397[2] = add_80396 == 32'h0000_0002 ? 32'h0000_0000 : array_index_80394[2];
  assign array_update_80397[3] = add_80396 == 32'h0000_0003 ? 32'h0000_0000 : array_index_80394[3];
  assign array_update_80397[4] = add_80396 == 32'h0000_0004 ? 32'h0000_0000 : array_index_80394[4];
  assign array_update_80397[5] = add_80396 == 32'h0000_0005 ? 32'h0000_0000 : array_index_80394[5];
  assign array_update_80397[6] = add_80396 == 32'h0000_0006 ? 32'h0000_0000 : array_index_80394[6];
  assign array_update_80397[7] = add_80396 == 32'h0000_0007 ? 32'h0000_0000 : array_index_80394[7];
  assign array_update_80397[8] = add_80396 == 32'h0000_0008 ? 32'h0000_0000 : array_index_80394[8];
  assign array_update_80397[9] = add_80396 == 32'h0000_0009 ? 32'h0000_0000 : array_index_80394[9];
  assign literal_80398 = 32'h0000_0000;
  assign array_update_80399[0] = add_80123 == 32'h0000_0000 ? array_update_80397 : array_update_80392[0];
  assign array_update_80399[1] = add_80123 == 32'h0000_0001 ? array_update_80397 : array_update_80392[1];
  assign array_update_80399[2] = add_80123 == 32'h0000_0002 ? array_update_80397 : array_update_80392[2];
  assign array_update_80399[3] = add_80123 == 32'h0000_0003 ? array_update_80397 : array_update_80392[3];
  assign array_update_80399[4] = add_80123 == 32'h0000_0004 ? array_update_80397 : array_update_80392[4];
  assign array_update_80399[5] = add_80123 == 32'h0000_0005 ? array_update_80397 : array_update_80392[5];
  assign array_update_80399[6] = add_80123 == 32'h0000_0006 ? array_update_80397 : array_update_80392[6];
  assign array_update_80399[7] = add_80123 == 32'h0000_0007 ? array_update_80397 : array_update_80392[7];
  assign array_update_80399[8] = add_80123 == 32'h0000_0008 ? array_update_80397 : array_update_80392[8];
  assign array_update_80399[9] = add_80123 == 32'h0000_0009 ? array_update_80397 : array_update_80392[9];
  assign array_index_80401 = array_update_72021[literal_80398 > 32'h0000_0009 ? 4'h9 : literal_80398[3:0]];
  assign array_index_80402 = array_update_80399[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_80406 = smul32b_32b_x_32b(array_index_80130[literal_80398 > 32'h0000_0009 ? 4'h9 : literal_80398[3:0]], array_index_80401[add_80396 > 32'h0000_0009 ? 4'h9 : add_80396[3:0]]);
  assign add_80408 = array_index_80402[add_80396 > 32'h0000_0009 ? 4'h9 : add_80396[3:0]] + smul_80406;
  assign array_update_80410[0] = add_80396 == 32'h0000_0000 ? add_80408 : array_index_80402[0];
  assign array_update_80410[1] = add_80396 == 32'h0000_0001 ? add_80408 : array_index_80402[1];
  assign array_update_80410[2] = add_80396 == 32'h0000_0002 ? add_80408 : array_index_80402[2];
  assign array_update_80410[3] = add_80396 == 32'h0000_0003 ? add_80408 : array_index_80402[3];
  assign array_update_80410[4] = add_80396 == 32'h0000_0004 ? add_80408 : array_index_80402[4];
  assign array_update_80410[5] = add_80396 == 32'h0000_0005 ? add_80408 : array_index_80402[5];
  assign array_update_80410[6] = add_80396 == 32'h0000_0006 ? add_80408 : array_index_80402[6];
  assign array_update_80410[7] = add_80396 == 32'h0000_0007 ? add_80408 : array_index_80402[7];
  assign array_update_80410[8] = add_80396 == 32'h0000_0008 ? add_80408 : array_index_80402[8];
  assign array_update_80410[9] = add_80396 == 32'h0000_0009 ? add_80408 : array_index_80402[9];
  assign add_80411 = literal_80398 + 32'h0000_0001;
  assign array_update_80412[0] = add_80123 == 32'h0000_0000 ? array_update_80410 : array_update_80399[0];
  assign array_update_80412[1] = add_80123 == 32'h0000_0001 ? array_update_80410 : array_update_80399[1];
  assign array_update_80412[2] = add_80123 == 32'h0000_0002 ? array_update_80410 : array_update_80399[2];
  assign array_update_80412[3] = add_80123 == 32'h0000_0003 ? array_update_80410 : array_update_80399[3];
  assign array_update_80412[4] = add_80123 == 32'h0000_0004 ? array_update_80410 : array_update_80399[4];
  assign array_update_80412[5] = add_80123 == 32'h0000_0005 ? array_update_80410 : array_update_80399[5];
  assign array_update_80412[6] = add_80123 == 32'h0000_0006 ? array_update_80410 : array_update_80399[6];
  assign array_update_80412[7] = add_80123 == 32'h0000_0007 ? array_update_80410 : array_update_80399[7];
  assign array_update_80412[8] = add_80123 == 32'h0000_0008 ? array_update_80410 : array_update_80399[8];
  assign array_update_80412[9] = add_80123 == 32'h0000_0009 ? array_update_80410 : array_update_80399[9];
  assign array_index_80414 = array_update_72021[add_80411 > 32'h0000_0009 ? 4'h9 : add_80411[3:0]];
  assign array_index_80415 = array_update_80412[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_80419 = smul32b_32b_x_32b(array_index_80130[add_80411 > 32'h0000_0009 ? 4'h9 : add_80411[3:0]], array_index_80414[add_80396 > 32'h0000_0009 ? 4'h9 : add_80396[3:0]]);
  assign add_80421 = array_index_80415[add_80396 > 32'h0000_0009 ? 4'h9 : add_80396[3:0]] + smul_80419;
  assign array_update_80423[0] = add_80396 == 32'h0000_0000 ? add_80421 : array_index_80415[0];
  assign array_update_80423[1] = add_80396 == 32'h0000_0001 ? add_80421 : array_index_80415[1];
  assign array_update_80423[2] = add_80396 == 32'h0000_0002 ? add_80421 : array_index_80415[2];
  assign array_update_80423[3] = add_80396 == 32'h0000_0003 ? add_80421 : array_index_80415[3];
  assign array_update_80423[4] = add_80396 == 32'h0000_0004 ? add_80421 : array_index_80415[4];
  assign array_update_80423[5] = add_80396 == 32'h0000_0005 ? add_80421 : array_index_80415[5];
  assign array_update_80423[6] = add_80396 == 32'h0000_0006 ? add_80421 : array_index_80415[6];
  assign array_update_80423[7] = add_80396 == 32'h0000_0007 ? add_80421 : array_index_80415[7];
  assign array_update_80423[8] = add_80396 == 32'h0000_0008 ? add_80421 : array_index_80415[8];
  assign array_update_80423[9] = add_80396 == 32'h0000_0009 ? add_80421 : array_index_80415[9];
  assign add_80424 = add_80411 + 32'h0000_0001;
  assign array_update_80425[0] = add_80123 == 32'h0000_0000 ? array_update_80423 : array_update_80412[0];
  assign array_update_80425[1] = add_80123 == 32'h0000_0001 ? array_update_80423 : array_update_80412[1];
  assign array_update_80425[2] = add_80123 == 32'h0000_0002 ? array_update_80423 : array_update_80412[2];
  assign array_update_80425[3] = add_80123 == 32'h0000_0003 ? array_update_80423 : array_update_80412[3];
  assign array_update_80425[4] = add_80123 == 32'h0000_0004 ? array_update_80423 : array_update_80412[4];
  assign array_update_80425[5] = add_80123 == 32'h0000_0005 ? array_update_80423 : array_update_80412[5];
  assign array_update_80425[6] = add_80123 == 32'h0000_0006 ? array_update_80423 : array_update_80412[6];
  assign array_update_80425[7] = add_80123 == 32'h0000_0007 ? array_update_80423 : array_update_80412[7];
  assign array_update_80425[8] = add_80123 == 32'h0000_0008 ? array_update_80423 : array_update_80412[8];
  assign array_update_80425[9] = add_80123 == 32'h0000_0009 ? array_update_80423 : array_update_80412[9];
  assign array_index_80427 = array_update_72021[add_80424 > 32'h0000_0009 ? 4'h9 : add_80424[3:0]];
  assign array_index_80428 = array_update_80425[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_80432 = smul32b_32b_x_32b(array_index_80130[add_80424 > 32'h0000_0009 ? 4'h9 : add_80424[3:0]], array_index_80427[add_80396 > 32'h0000_0009 ? 4'h9 : add_80396[3:0]]);
  assign add_80434 = array_index_80428[add_80396 > 32'h0000_0009 ? 4'h9 : add_80396[3:0]] + smul_80432;
  assign array_update_80436[0] = add_80396 == 32'h0000_0000 ? add_80434 : array_index_80428[0];
  assign array_update_80436[1] = add_80396 == 32'h0000_0001 ? add_80434 : array_index_80428[1];
  assign array_update_80436[2] = add_80396 == 32'h0000_0002 ? add_80434 : array_index_80428[2];
  assign array_update_80436[3] = add_80396 == 32'h0000_0003 ? add_80434 : array_index_80428[3];
  assign array_update_80436[4] = add_80396 == 32'h0000_0004 ? add_80434 : array_index_80428[4];
  assign array_update_80436[5] = add_80396 == 32'h0000_0005 ? add_80434 : array_index_80428[5];
  assign array_update_80436[6] = add_80396 == 32'h0000_0006 ? add_80434 : array_index_80428[6];
  assign array_update_80436[7] = add_80396 == 32'h0000_0007 ? add_80434 : array_index_80428[7];
  assign array_update_80436[8] = add_80396 == 32'h0000_0008 ? add_80434 : array_index_80428[8];
  assign array_update_80436[9] = add_80396 == 32'h0000_0009 ? add_80434 : array_index_80428[9];
  assign add_80437 = add_80424 + 32'h0000_0001;
  assign array_update_80438[0] = add_80123 == 32'h0000_0000 ? array_update_80436 : array_update_80425[0];
  assign array_update_80438[1] = add_80123 == 32'h0000_0001 ? array_update_80436 : array_update_80425[1];
  assign array_update_80438[2] = add_80123 == 32'h0000_0002 ? array_update_80436 : array_update_80425[2];
  assign array_update_80438[3] = add_80123 == 32'h0000_0003 ? array_update_80436 : array_update_80425[3];
  assign array_update_80438[4] = add_80123 == 32'h0000_0004 ? array_update_80436 : array_update_80425[4];
  assign array_update_80438[5] = add_80123 == 32'h0000_0005 ? array_update_80436 : array_update_80425[5];
  assign array_update_80438[6] = add_80123 == 32'h0000_0006 ? array_update_80436 : array_update_80425[6];
  assign array_update_80438[7] = add_80123 == 32'h0000_0007 ? array_update_80436 : array_update_80425[7];
  assign array_update_80438[8] = add_80123 == 32'h0000_0008 ? array_update_80436 : array_update_80425[8];
  assign array_update_80438[9] = add_80123 == 32'h0000_0009 ? array_update_80436 : array_update_80425[9];
  assign array_index_80440 = array_update_72021[add_80437 > 32'h0000_0009 ? 4'h9 : add_80437[3:0]];
  assign array_index_80441 = array_update_80438[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_80445 = smul32b_32b_x_32b(array_index_80130[add_80437 > 32'h0000_0009 ? 4'h9 : add_80437[3:0]], array_index_80440[add_80396 > 32'h0000_0009 ? 4'h9 : add_80396[3:0]]);
  assign add_80447 = array_index_80441[add_80396 > 32'h0000_0009 ? 4'h9 : add_80396[3:0]] + smul_80445;
  assign array_update_80449[0] = add_80396 == 32'h0000_0000 ? add_80447 : array_index_80441[0];
  assign array_update_80449[1] = add_80396 == 32'h0000_0001 ? add_80447 : array_index_80441[1];
  assign array_update_80449[2] = add_80396 == 32'h0000_0002 ? add_80447 : array_index_80441[2];
  assign array_update_80449[3] = add_80396 == 32'h0000_0003 ? add_80447 : array_index_80441[3];
  assign array_update_80449[4] = add_80396 == 32'h0000_0004 ? add_80447 : array_index_80441[4];
  assign array_update_80449[5] = add_80396 == 32'h0000_0005 ? add_80447 : array_index_80441[5];
  assign array_update_80449[6] = add_80396 == 32'h0000_0006 ? add_80447 : array_index_80441[6];
  assign array_update_80449[7] = add_80396 == 32'h0000_0007 ? add_80447 : array_index_80441[7];
  assign array_update_80449[8] = add_80396 == 32'h0000_0008 ? add_80447 : array_index_80441[8];
  assign array_update_80449[9] = add_80396 == 32'h0000_0009 ? add_80447 : array_index_80441[9];
  assign add_80450 = add_80437 + 32'h0000_0001;
  assign array_update_80451[0] = add_80123 == 32'h0000_0000 ? array_update_80449 : array_update_80438[0];
  assign array_update_80451[1] = add_80123 == 32'h0000_0001 ? array_update_80449 : array_update_80438[1];
  assign array_update_80451[2] = add_80123 == 32'h0000_0002 ? array_update_80449 : array_update_80438[2];
  assign array_update_80451[3] = add_80123 == 32'h0000_0003 ? array_update_80449 : array_update_80438[3];
  assign array_update_80451[4] = add_80123 == 32'h0000_0004 ? array_update_80449 : array_update_80438[4];
  assign array_update_80451[5] = add_80123 == 32'h0000_0005 ? array_update_80449 : array_update_80438[5];
  assign array_update_80451[6] = add_80123 == 32'h0000_0006 ? array_update_80449 : array_update_80438[6];
  assign array_update_80451[7] = add_80123 == 32'h0000_0007 ? array_update_80449 : array_update_80438[7];
  assign array_update_80451[8] = add_80123 == 32'h0000_0008 ? array_update_80449 : array_update_80438[8];
  assign array_update_80451[9] = add_80123 == 32'h0000_0009 ? array_update_80449 : array_update_80438[9];
  assign array_index_80453 = array_update_72021[add_80450 > 32'h0000_0009 ? 4'h9 : add_80450[3:0]];
  assign array_index_80454 = array_update_80451[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_80458 = smul32b_32b_x_32b(array_index_80130[add_80450 > 32'h0000_0009 ? 4'h9 : add_80450[3:0]], array_index_80453[add_80396 > 32'h0000_0009 ? 4'h9 : add_80396[3:0]]);
  assign add_80460 = array_index_80454[add_80396 > 32'h0000_0009 ? 4'h9 : add_80396[3:0]] + smul_80458;
  assign array_update_80462[0] = add_80396 == 32'h0000_0000 ? add_80460 : array_index_80454[0];
  assign array_update_80462[1] = add_80396 == 32'h0000_0001 ? add_80460 : array_index_80454[1];
  assign array_update_80462[2] = add_80396 == 32'h0000_0002 ? add_80460 : array_index_80454[2];
  assign array_update_80462[3] = add_80396 == 32'h0000_0003 ? add_80460 : array_index_80454[3];
  assign array_update_80462[4] = add_80396 == 32'h0000_0004 ? add_80460 : array_index_80454[4];
  assign array_update_80462[5] = add_80396 == 32'h0000_0005 ? add_80460 : array_index_80454[5];
  assign array_update_80462[6] = add_80396 == 32'h0000_0006 ? add_80460 : array_index_80454[6];
  assign array_update_80462[7] = add_80396 == 32'h0000_0007 ? add_80460 : array_index_80454[7];
  assign array_update_80462[8] = add_80396 == 32'h0000_0008 ? add_80460 : array_index_80454[8];
  assign array_update_80462[9] = add_80396 == 32'h0000_0009 ? add_80460 : array_index_80454[9];
  assign add_80463 = add_80450 + 32'h0000_0001;
  assign array_update_80464[0] = add_80123 == 32'h0000_0000 ? array_update_80462 : array_update_80451[0];
  assign array_update_80464[1] = add_80123 == 32'h0000_0001 ? array_update_80462 : array_update_80451[1];
  assign array_update_80464[2] = add_80123 == 32'h0000_0002 ? array_update_80462 : array_update_80451[2];
  assign array_update_80464[3] = add_80123 == 32'h0000_0003 ? array_update_80462 : array_update_80451[3];
  assign array_update_80464[4] = add_80123 == 32'h0000_0004 ? array_update_80462 : array_update_80451[4];
  assign array_update_80464[5] = add_80123 == 32'h0000_0005 ? array_update_80462 : array_update_80451[5];
  assign array_update_80464[6] = add_80123 == 32'h0000_0006 ? array_update_80462 : array_update_80451[6];
  assign array_update_80464[7] = add_80123 == 32'h0000_0007 ? array_update_80462 : array_update_80451[7];
  assign array_update_80464[8] = add_80123 == 32'h0000_0008 ? array_update_80462 : array_update_80451[8];
  assign array_update_80464[9] = add_80123 == 32'h0000_0009 ? array_update_80462 : array_update_80451[9];
  assign array_index_80466 = array_update_72021[add_80463 > 32'h0000_0009 ? 4'h9 : add_80463[3:0]];
  assign array_index_80467 = array_update_80464[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_80471 = smul32b_32b_x_32b(array_index_80130[add_80463 > 32'h0000_0009 ? 4'h9 : add_80463[3:0]], array_index_80466[add_80396 > 32'h0000_0009 ? 4'h9 : add_80396[3:0]]);
  assign add_80473 = array_index_80467[add_80396 > 32'h0000_0009 ? 4'h9 : add_80396[3:0]] + smul_80471;
  assign array_update_80475[0] = add_80396 == 32'h0000_0000 ? add_80473 : array_index_80467[0];
  assign array_update_80475[1] = add_80396 == 32'h0000_0001 ? add_80473 : array_index_80467[1];
  assign array_update_80475[2] = add_80396 == 32'h0000_0002 ? add_80473 : array_index_80467[2];
  assign array_update_80475[3] = add_80396 == 32'h0000_0003 ? add_80473 : array_index_80467[3];
  assign array_update_80475[4] = add_80396 == 32'h0000_0004 ? add_80473 : array_index_80467[4];
  assign array_update_80475[5] = add_80396 == 32'h0000_0005 ? add_80473 : array_index_80467[5];
  assign array_update_80475[6] = add_80396 == 32'h0000_0006 ? add_80473 : array_index_80467[6];
  assign array_update_80475[7] = add_80396 == 32'h0000_0007 ? add_80473 : array_index_80467[7];
  assign array_update_80475[8] = add_80396 == 32'h0000_0008 ? add_80473 : array_index_80467[8];
  assign array_update_80475[9] = add_80396 == 32'h0000_0009 ? add_80473 : array_index_80467[9];
  assign add_80476 = add_80463 + 32'h0000_0001;
  assign array_update_80477[0] = add_80123 == 32'h0000_0000 ? array_update_80475 : array_update_80464[0];
  assign array_update_80477[1] = add_80123 == 32'h0000_0001 ? array_update_80475 : array_update_80464[1];
  assign array_update_80477[2] = add_80123 == 32'h0000_0002 ? array_update_80475 : array_update_80464[2];
  assign array_update_80477[3] = add_80123 == 32'h0000_0003 ? array_update_80475 : array_update_80464[3];
  assign array_update_80477[4] = add_80123 == 32'h0000_0004 ? array_update_80475 : array_update_80464[4];
  assign array_update_80477[5] = add_80123 == 32'h0000_0005 ? array_update_80475 : array_update_80464[5];
  assign array_update_80477[6] = add_80123 == 32'h0000_0006 ? array_update_80475 : array_update_80464[6];
  assign array_update_80477[7] = add_80123 == 32'h0000_0007 ? array_update_80475 : array_update_80464[7];
  assign array_update_80477[8] = add_80123 == 32'h0000_0008 ? array_update_80475 : array_update_80464[8];
  assign array_update_80477[9] = add_80123 == 32'h0000_0009 ? array_update_80475 : array_update_80464[9];
  assign array_index_80479 = array_update_72021[add_80476 > 32'h0000_0009 ? 4'h9 : add_80476[3:0]];
  assign array_index_80480 = array_update_80477[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_80484 = smul32b_32b_x_32b(array_index_80130[add_80476 > 32'h0000_0009 ? 4'h9 : add_80476[3:0]], array_index_80479[add_80396 > 32'h0000_0009 ? 4'h9 : add_80396[3:0]]);
  assign add_80486 = array_index_80480[add_80396 > 32'h0000_0009 ? 4'h9 : add_80396[3:0]] + smul_80484;
  assign array_update_80488[0] = add_80396 == 32'h0000_0000 ? add_80486 : array_index_80480[0];
  assign array_update_80488[1] = add_80396 == 32'h0000_0001 ? add_80486 : array_index_80480[1];
  assign array_update_80488[2] = add_80396 == 32'h0000_0002 ? add_80486 : array_index_80480[2];
  assign array_update_80488[3] = add_80396 == 32'h0000_0003 ? add_80486 : array_index_80480[3];
  assign array_update_80488[4] = add_80396 == 32'h0000_0004 ? add_80486 : array_index_80480[4];
  assign array_update_80488[5] = add_80396 == 32'h0000_0005 ? add_80486 : array_index_80480[5];
  assign array_update_80488[6] = add_80396 == 32'h0000_0006 ? add_80486 : array_index_80480[6];
  assign array_update_80488[7] = add_80396 == 32'h0000_0007 ? add_80486 : array_index_80480[7];
  assign array_update_80488[8] = add_80396 == 32'h0000_0008 ? add_80486 : array_index_80480[8];
  assign array_update_80488[9] = add_80396 == 32'h0000_0009 ? add_80486 : array_index_80480[9];
  assign add_80489 = add_80476 + 32'h0000_0001;
  assign array_update_80490[0] = add_80123 == 32'h0000_0000 ? array_update_80488 : array_update_80477[0];
  assign array_update_80490[1] = add_80123 == 32'h0000_0001 ? array_update_80488 : array_update_80477[1];
  assign array_update_80490[2] = add_80123 == 32'h0000_0002 ? array_update_80488 : array_update_80477[2];
  assign array_update_80490[3] = add_80123 == 32'h0000_0003 ? array_update_80488 : array_update_80477[3];
  assign array_update_80490[4] = add_80123 == 32'h0000_0004 ? array_update_80488 : array_update_80477[4];
  assign array_update_80490[5] = add_80123 == 32'h0000_0005 ? array_update_80488 : array_update_80477[5];
  assign array_update_80490[6] = add_80123 == 32'h0000_0006 ? array_update_80488 : array_update_80477[6];
  assign array_update_80490[7] = add_80123 == 32'h0000_0007 ? array_update_80488 : array_update_80477[7];
  assign array_update_80490[8] = add_80123 == 32'h0000_0008 ? array_update_80488 : array_update_80477[8];
  assign array_update_80490[9] = add_80123 == 32'h0000_0009 ? array_update_80488 : array_update_80477[9];
  assign array_index_80492 = array_update_72021[add_80489 > 32'h0000_0009 ? 4'h9 : add_80489[3:0]];
  assign array_index_80493 = array_update_80490[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_80497 = smul32b_32b_x_32b(array_index_80130[add_80489 > 32'h0000_0009 ? 4'h9 : add_80489[3:0]], array_index_80492[add_80396 > 32'h0000_0009 ? 4'h9 : add_80396[3:0]]);
  assign add_80499 = array_index_80493[add_80396 > 32'h0000_0009 ? 4'h9 : add_80396[3:0]] + smul_80497;
  assign array_update_80501[0] = add_80396 == 32'h0000_0000 ? add_80499 : array_index_80493[0];
  assign array_update_80501[1] = add_80396 == 32'h0000_0001 ? add_80499 : array_index_80493[1];
  assign array_update_80501[2] = add_80396 == 32'h0000_0002 ? add_80499 : array_index_80493[2];
  assign array_update_80501[3] = add_80396 == 32'h0000_0003 ? add_80499 : array_index_80493[3];
  assign array_update_80501[4] = add_80396 == 32'h0000_0004 ? add_80499 : array_index_80493[4];
  assign array_update_80501[5] = add_80396 == 32'h0000_0005 ? add_80499 : array_index_80493[5];
  assign array_update_80501[6] = add_80396 == 32'h0000_0006 ? add_80499 : array_index_80493[6];
  assign array_update_80501[7] = add_80396 == 32'h0000_0007 ? add_80499 : array_index_80493[7];
  assign array_update_80501[8] = add_80396 == 32'h0000_0008 ? add_80499 : array_index_80493[8];
  assign array_update_80501[9] = add_80396 == 32'h0000_0009 ? add_80499 : array_index_80493[9];
  assign add_80502 = add_80489 + 32'h0000_0001;
  assign array_update_80503[0] = add_80123 == 32'h0000_0000 ? array_update_80501 : array_update_80490[0];
  assign array_update_80503[1] = add_80123 == 32'h0000_0001 ? array_update_80501 : array_update_80490[1];
  assign array_update_80503[2] = add_80123 == 32'h0000_0002 ? array_update_80501 : array_update_80490[2];
  assign array_update_80503[3] = add_80123 == 32'h0000_0003 ? array_update_80501 : array_update_80490[3];
  assign array_update_80503[4] = add_80123 == 32'h0000_0004 ? array_update_80501 : array_update_80490[4];
  assign array_update_80503[5] = add_80123 == 32'h0000_0005 ? array_update_80501 : array_update_80490[5];
  assign array_update_80503[6] = add_80123 == 32'h0000_0006 ? array_update_80501 : array_update_80490[6];
  assign array_update_80503[7] = add_80123 == 32'h0000_0007 ? array_update_80501 : array_update_80490[7];
  assign array_update_80503[8] = add_80123 == 32'h0000_0008 ? array_update_80501 : array_update_80490[8];
  assign array_update_80503[9] = add_80123 == 32'h0000_0009 ? array_update_80501 : array_update_80490[9];
  assign array_index_80505 = array_update_72021[add_80502 > 32'h0000_0009 ? 4'h9 : add_80502[3:0]];
  assign array_index_80506 = array_update_80503[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_80510 = smul32b_32b_x_32b(array_index_80130[add_80502 > 32'h0000_0009 ? 4'h9 : add_80502[3:0]], array_index_80505[add_80396 > 32'h0000_0009 ? 4'h9 : add_80396[3:0]]);
  assign add_80512 = array_index_80506[add_80396 > 32'h0000_0009 ? 4'h9 : add_80396[3:0]] + smul_80510;
  assign array_update_80514[0] = add_80396 == 32'h0000_0000 ? add_80512 : array_index_80506[0];
  assign array_update_80514[1] = add_80396 == 32'h0000_0001 ? add_80512 : array_index_80506[1];
  assign array_update_80514[2] = add_80396 == 32'h0000_0002 ? add_80512 : array_index_80506[2];
  assign array_update_80514[3] = add_80396 == 32'h0000_0003 ? add_80512 : array_index_80506[3];
  assign array_update_80514[4] = add_80396 == 32'h0000_0004 ? add_80512 : array_index_80506[4];
  assign array_update_80514[5] = add_80396 == 32'h0000_0005 ? add_80512 : array_index_80506[5];
  assign array_update_80514[6] = add_80396 == 32'h0000_0006 ? add_80512 : array_index_80506[6];
  assign array_update_80514[7] = add_80396 == 32'h0000_0007 ? add_80512 : array_index_80506[7];
  assign array_update_80514[8] = add_80396 == 32'h0000_0008 ? add_80512 : array_index_80506[8];
  assign array_update_80514[9] = add_80396 == 32'h0000_0009 ? add_80512 : array_index_80506[9];
  assign add_80515 = add_80502 + 32'h0000_0001;
  assign array_update_80516[0] = add_80123 == 32'h0000_0000 ? array_update_80514 : array_update_80503[0];
  assign array_update_80516[1] = add_80123 == 32'h0000_0001 ? array_update_80514 : array_update_80503[1];
  assign array_update_80516[2] = add_80123 == 32'h0000_0002 ? array_update_80514 : array_update_80503[2];
  assign array_update_80516[3] = add_80123 == 32'h0000_0003 ? array_update_80514 : array_update_80503[3];
  assign array_update_80516[4] = add_80123 == 32'h0000_0004 ? array_update_80514 : array_update_80503[4];
  assign array_update_80516[5] = add_80123 == 32'h0000_0005 ? array_update_80514 : array_update_80503[5];
  assign array_update_80516[6] = add_80123 == 32'h0000_0006 ? array_update_80514 : array_update_80503[6];
  assign array_update_80516[7] = add_80123 == 32'h0000_0007 ? array_update_80514 : array_update_80503[7];
  assign array_update_80516[8] = add_80123 == 32'h0000_0008 ? array_update_80514 : array_update_80503[8];
  assign array_update_80516[9] = add_80123 == 32'h0000_0009 ? array_update_80514 : array_update_80503[9];
  assign array_index_80518 = array_update_72021[add_80515 > 32'h0000_0009 ? 4'h9 : add_80515[3:0]];
  assign array_index_80519 = array_update_80516[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_80523 = smul32b_32b_x_32b(array_index_80130[add_80515 > 32'h0000_0009 ? 4'h9 : add_80515[3:0]], array_index_80518[add_80396 > 32'h0000_0009 ? 4'h9 : add_80396[3:0]]);
  assign add_80525 = array_index_80519[add_80396 > 32'h0000_0009 ? 4'h9 : add_80396[3:0]] + smul_80523;
  assign array_update_80526[0] = add_80396 == 32'h0000_0000 ? add_80525 : array_index_80519[0];
  assign array_update_80526[1] = add_80396 == 32'h0000_0001 ? add_80525 : array_index_80519[1];
  assign array_update_80526[2] = add_80396 == 32'h0000_0002 ? add_80525 : array_index_80519[2];
  assign array_update_80526[3] = add_80396 == 32'h0000_0003 ? add_80525 : array_index_80519[3];
  assign array_update_80526[4] = add_80396 == 32'h0000_0004 ? add_80525 : array_index_80519[4];
  assign array_update_80526[5] = add_80396 == 32'h0000_0005 ? add_80525 : array_index_80519[5];
  assign array_update_80526[6] = add_80396 == 32'h0000_0006 ? add_80525 : array_index_80519[6];
  assign array_update_80526[7] = add_80396 == 32'h0000_0007 ? add_80525 : array_index_80519[7];
  assign array_update_80526[8] = add_80396 == 32'h0000_0008 ? add_80525 : array_index_80519[8];
  assign array_update_80526[9] = add_80396 == 32'h0000_0009 ? add_80525 : array_index_80519[9];
  assign array_update_80527[0] = add_80123 == 32'h0000_0000 ? array_update_80526 : array_update_80516[0];
  assign array_update_80527[1] = add_80123 == 32'h0000_0001 ? array_update_80526 : array_update_80516[1];
  assign array_update_80527[2] = add_80123 == 32'h0000_0002 ? array_update_80526 : array_update_80516[2];
  assign array_update_80527[3] = add_80123 == 32'h0000_0003 ? array_update_80526 : array_update_80516[3];
  assign array_update_80527[4] = add_80123 == 32'h0000_0004 ? array_update_80526 : array_update_80516[4];
  assign array_update_80527[5] = add_80123 == 32'h0000_0005 ? array_update_80526 : array_update_80516[5];
  assign array_update_80527[6] = add_80123 == 32'h0000_0006 ? array_update_80526 : array_update_80516[6];
  assign array_update_80527[7] = add_80123 == 32'h0000_0007 ? array_update_80526 : array_update_80516[7];
  assign array_update_80527[8] = add_80123 == 32'h0000_0008 ? array_update_80526 : array_update_80516[8];
  assign array_update_80527[9] = add_80123 == 32'h0000_0009 ? array_update_80526 : array_update_80516[9];
  assign array_index_80529 = array_update_80527[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign add_80531 = add_80396 + 32'h0000_0001;
  assign array_update_80532[0] = add_80531 == 32'h0000_0000 ? 32'h0000_0000 : array_index_80529[0];
  assign array_update_80532[1] = add_80531 == 32'h0000_0001 ? 32'h0000_0000 : array_index_80529[1];
  assign array_update_80532[2] = add_80531 == 32'h0000_0002 ? 32'h0000_0000 : array_index_80529[2];
  assign array_update_80532[3] = add_80531 == 32'h0000_0003 ? 32'h0000_0000 : array_index_80529[3];
  assign array_update_80532[4] = add_80531 == 32'h0000_0004 ? 32'h0000_0000 : array_index_80529[4];
  assign array_update_80532[5] = add_80531 == 32'h0000_0005 ? 32'h0000_0000 : array_index_80529[5];
  assign array_update_80532[6] = add_80531 == 32'h0000_0006 ? 32'h0000_0000 : array_index_80529[6];
  assign array_update_80532[7] = add_80531 == 32'h0000_0007 ? 32'h0000_0000 : array_index_80529[7];
  assign array_update_80532[8] = add_80531 == 32'h0000_0008 ? 32'h0000_0000 : array_index_80529[8];
  assign array_update_80532[9] = add_80531 == 32'h0000_0009 ? 32'h0000_0000 : array_index_80529[9];
  assign literal_80533 = 32'h0000_0000;
  assign array_update_80534[0] = add_80123 == 32'h0000_0000 ? array_update_80532 : array_update_80527[0];
  assign array_update_80534[1] = add_80123 == 32'h0000_0001 ? array_update_80532 : array_update_80527[1];
  assign array_update_80534[2] = add_80123 == 32'h0000_0002 ? array_update_80532 : array_update_80527[2];
  assign array_update_80534[3] = add_80123 == 32'h0000_0003 ? array_update_80532 : array_update_80527[3];
  assign array_update_80534[4] = add_80123 == 32'h0000_0004 ? array_update_80532 : array_update_80527[4];
  assign array_update_80534[5] = add_80123 == 32'h0000_0005 ? array_update_80532 : array_update_80527[5];
  assign array_update_80534[6] = add_80123 == 32'h0000_0006 ? array_update_80532 : array_update_80527[6];
  assign array_update_80534[7] = add_80123 == 32'h0000_0007 ? array_update_80532 : array_update_80527[7];
  assign array_update_80534[8] = add_80123 == 32'h0000_0008 ? array_update_80532 : array_update_80527[8];
  assign array_update_80534[9] = add_80123 == 32'h0000_0009 ? array_update_80532 : array_update_80527[9];
  assign array_index_80536 = array_update_72021[literal_80533 > 32'h0000_0009 ? 4'h9 : literal_80533[3:0]];
  assign array_index_80537 = array_update_80534[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_80541 = smul32b_32b_x_32b(array_index_80130[literal_80533 > 32'h0000_0009 ? 4'h9 : literal_80533[3:0]], array_index_80536[add_80531 > 32'h0000_0009 ? 4'h9 : add_80531[3:0]]);
  assign add_80543 = array_index_80537[add_80531 > 32'h0000_0009 ? 4'h9 : add_80531[3:0]] + smul_80541;
  assign array_update_80545[0] = add_80531 == 32'h0000_0000 ? add_80543 : array_index_80537[0];
  assign array_update_80545[1] = add_80531 == 32'h0000_0001 ? add_80543 : array_index_80537[1];
  assign array_update_80545[2] = add_80531 == 32'h0000_0002 ? add_80543 : array_index_80537[2];
  assign array_update_80545[3] = add_80531 == 32'h0000_0003 ? add_80543 : array_index_80537[3];
  assign array_update_80545[4] = add_80531 == 32'h0000_0004 ? add_80543 : array_index_80537[4];
  assign array_update_80545[5] = add_80531 == 32'h0000_0005 ? add_80543 : array_index_80537[5];
  assign array_update_80545[6] = add_80531 == 32'h0000_0006 ? add_80543 : array_index_80537[6];
  assign array_update_80545[7] = add_80531 == 32'h0000_0007 ? add_80543 : array_index_80537[7];
  assign array_update_80545[8] = add_80531 == 32'h0000_0008 ? add_80543 : array_index_80537[8];
  assign array_update_80545[9] = add_80531 == 32'h0000_0009 ? add_80543 : array_index_80537[9];
  assign add_80546 = literal_80533 + 32'h0000_0001;
  assign array_update_80547[0] = add_80123 == 32'h0000_0000 ? array_update_80545 : array_update_80534[0];
  assign array_update_80547[1] = add_80123 == 32'h0000_0001 ? array_update_80545 : array_update_80534[1];
  assign array_update_80547[2] = add_80123 == 32'h0000_0002 ? array_update_80545 : array_update_80534[2];
  assign array_update_80547[3] = add_80123 == 32'h0000_0003 ? array_update_80545 : array_update_80534[3];
  assign array_update_80547[4] = add_80123 == 32'h0000_0004 ? array_update_80545 : array_update_80534[4];
  assign array_update_80547[5] = add_80123 == 32'h0000_0005 ? array_update_80545 : array_update_80534[5];
  assign array_update_80547[6] = add_80123 == 32'h0000_0006 ? array_update_80545 : array_update_80534[6];
  assign array_update_80547[7] = add_80123 == 32'h0000_0007 ? array_update_80545 : array_update_80534[7];
  assign array_update_80547[8] = add_80123 == 32'h0000_0008 ? array_update_80545 : array_update_80534[8];
  assign array_update_80547[9] = add_80123 == 32'h0000_0009 ? array_update_80545 : array_update_80534[9];
  assign array_index_80549 = array_update_72021[add_80546 > 32'h0000_0009 ? 4'h9 : add_80546[3:0]];
  assign array_index_80550 = array_update_80547[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_80554 = smul32b_32b_x_32b(array_index_80130[add_80546 > 32'h0000_0009 ? 4'h9 : add_80546[3:0]], array_index_80549[add_80531 > 32'h0000_0009 ? 4'h9 : add_80531[3:0]]);
  assign add_80556 = array_index_80550[add_80531 > 32'h0000_0009 ? 4'h9 : add_80531[3:0]] + smul_80554;
  assign array_update_80558[0] = add_80531 == 32'h0000_0000 ? add_80556 : array_index_80550[0];
  assign array_update_80558[1] = add_80531 == 32'h0000_0001 ? add_80556 : array_index_80550[1];
  assign array_update_80558[2] = add_80531 == 32'h0000_0002 ? add_80556 : array_index_80550[2];
  assign array_update_80558[3] = add_80531 == 32'h0000_0003 ? add_80556 : array_index_80550[3];
  assign array_update_80558[4] = add_80531 == 32'h0000_0004 ? add_80556 : array_index_80550[4];
  assign array_update_80558[5] = add_80531 == 32'h0000_0005 ? add_80556 : array_index_80550[5];
  assign array_update_80558[6] = add_80531 == 32'h0000_0006 ? add_80556 : array_index_80550[6];
  assign array_update_80558[7] = add_80531 == 32'h0000_0007 ? add_80556 : array_index_80550[7];
  assign array_update_80558[8] = add_80531 == 32'h0000_0008 ? add_80556 : array_index_80550[8];
  assign array_update_80558[9] = add_80531 == 32'h0000_0009 ? add_80556 : array_index_80550[9];
  assign add_80559 = add_80546 + 32'h0000_0001;
  assign array_update_80560[0] = add_80123 == 32'h0000_0000 ? array_update_80558 : array_update_80547[0];
  assign array_update_80560[1] = add_80123 == 32'h0000_0001 ? array_update_80558 : array_update_80547[1];
  assign array_update_80560[2] = add_80123 == 32'h0000_0002 ? array_update_80558 : array_update_80547[2];
  assign array_update_80560[3] = add_80123 == 32'h0000_0003 ? array_update_80558 : array_update_80547[3];
  assign array_update_80560[4] = add_80123 == 32'h0000_0004 ? array_update_80558 : array_update_80547[4];
  assign array_update_80560[5] = add_80123 == 32'h0000_0005 ? array_update_80558 : array_update_80547[5];
  assign array_update_80560[6] = add_80123 == 32'h0000_0006 ? array_update_80558 : array_update_80547[6];
  assign array_update_80560[7] = add_80123 == 32'h0000_0007 ? array_update_80558 : array_update_80547[7];
  assign array_update_80560[8] = add_80123 == 32'h0000_0008 ? array_update_80558 : array_update_80547[8];
  assign array_update_80560[9] = add_80123 == 32'h0000_0009 ? array_update_80558 : array_update_80547[9];
  assign array_index_80562 = array_update_72021[add_80559 > 32'h0000_0009 ? 4'h9 : add_80559[3:0]];
  assign array_index_80563 = array_update_80560[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_80567 = smul32b_32b_x_32b(array_index_80130[add_80559 > 32'h0000_0009 ? 4'h9 : add_80559[3:0]], array_index_80562[add_80531 > 32'h0000_0009 ? 4'h9 : add_80531[3:0]]);
  assign add_80569 = array_index_80563[add_80531 > 32'h0000_0009 ? 4'h9 : add_80531[3:0]] + smul_80567;
  assign array_update_80571[0] = add_80531 == 32'h0000_0000 ? add_80569 : array_index_80563[0];
  assign array_update_80571[1] = add_80531 == 32'h0000_0001 ? add_80569 : array_index_80563[1];
  assign array_update_80571[2] = add_80531 == 32'h0000_0002 ? add_80569 : array_index_80563[2];
  assign array_update_80571[3] = add_80531 == 32'h0000_0003 ? add_80569 : array_index_80563[3];
  assign array_update_80571[4] = add_80531 == 32'h0000_0004 ? add_80569 : array_index_80563[4];
  assign array_update_80571[5] = add_80531 == 32'h0000_0005 ? add_80569 : array_index_80563[5];
  assign array_update_80571[6] = add_80531 == 32'h0000_0006 ? add_80569 : array_index_80563[6];
  assign array_update_80571[7] = add_80531 == 32'h0000_0007 ? add_80569 : array_index_80563[7];
  assign array_update_80571[8] = add_80531 == 32'h0000_0008 ? add_80569 : array_index_80563[8];
  assign array_update_80571[9] = add_80531 == 32'h0000_0009 ? add_80569 : array_index_80563[9];
  assign add_80572 = add_80559 + 32'h0000_0001;
  assign array_update_80573[0] = add_80123 == 32'h0000_0000 ? array_update_80571 : array_update_80560[0];
  assign array_update_80573[1] = add_80123 == 32'h0000_0001 ? array_update_80571 : array_update_80560[1];
  assign array_update_80573[2] = add_80123 == 32'h0000_0002 ? array_update_80571 : array_update_80560[2];
  assign array_update_80573[3] = add_80123 == 32'h0000_0003 ? array_update_80571 : array_update_80560[3];
  assign array_update_80573[4] = add_80123 == 32'h0000_0004 ? array_update_80571 : array_update_80560[4];
  assign array_update_80573[5] = add_80123 == 32'h0000_0005 ? array_update_80571 : array_update_80560[5];
  assign array_update_80573[6] = add_80123 == 32'h0000_0006 ? array_update_80571 : array_update_80560[6];
  assign array_update_80573[7] = add_80123 == 32'h0000_0007 ? array_update_80571 : array_update_80560[7];
  assign array_update_80573[8] = add_80123 == 32'h0000_0008 ? array_update_80571 : array_update_80560[8];
  assign array_update_80573[9] = add_80123 == 32'h0000_0009 ? array_update_80571 : array_update_80560[9];
  assign array_index_80575 = array_update_72021[add_80572 > 32'h0000_0009 ? 4'h9 : add_80572[3:0]];
  assign array_index_80576 = array_update_80573[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_80580 = smul32b_32b_x_32b(array_index_80130[add_80572 > 32'h0000_0009 ? 4'h9 : add_80572[3:0]], array_index_80575[add_80531 > 32'h0000_0009 ? 4'h9 : add_80531[3:0]]);
  assign add_80582 = array_index_80576[add_80531 > 32'h0000_0009 ? 4'h9 : add_80531[3:0]] + smul_80580;
  assign array_update_80584[0] = add_80531 == 32'h0000_0000 ? add_80582 : array_index_80576[0];
  assign array_update_80584[1] = add_80531 == 32'h0000_0001 ? add_80582 : array_index_80576[1];
  assign array_update_80584[2] = add_80531 == 32'h0000_0002 ? add_80582 : array_index_80576[2];
  assign array_update_80584[3] = add_80531 == 32'h0000_0003 ? add_80582 : array_index_80576[3];
  assign array_update_80584[4] = add_80531 == 32'h0000_0004 ? add_80582 : array_index_80576[4];
  assign array_update_80584[5] = add_80531 == 32'h0000_0005 ? add_80582 : array_index_80576[5];
  assign array_update_80584[6] = add_80531 == 32'h0000_0006 ? add_80582 : array_index_80576[6];
  assign array_update_80584[7] = add_80531 == 32'h0000_0007 ? add_80582 : array_index_80576[7];
  assign array_update_80584[8] = add_80531 == 32'h0000_0008 ? add_80582 : array_index_80576[8];
  assign array_update_80584[9] = add_80531 == 32'h0000_0009 ? add_80582 : array_index_80576[9];
  assign add_80585 = add_80572 + 32'h0000_0001;
  assign array_update_80586[0] = add_80123 == 32'h0000_0000 ? array_update_80584 : array_update_80573[0];
  assign array_update_80586[1] = add_80123 == 32'h0000_0001 ? array_update_80584 : array_update_80573[1];
  assign array_update_80586[2] = add_80123 == 32'h0000_0002 ? array_update_80584 : array_update_80573[2];
  assign array_update_80586[3] = add_80123 == 32'h0000_0003 ? array_update_80584 : array_update_80573[3];
  assign array_update_80586[4] = add_80123 == 32'h0000_0004 ? array_update_80584 : array_update_80573[4];
  assign array_update_80586[5] = add_80123 == 32'h0000_0005 ? array_update_80584 : array_update_80573[5];
  assign array_update_80586[6] = add_80123 == 32'h0000_0006 ? array_update_80584 : array_update_80573[6];
  assign array_update_80586[7] = add_80123 == 32'h0000_0007 ? array_update_80584 : array_update_80573[7];
  assign array_update_80586[8] = add_80123 == 32'h0000_0008 ? array_update_80584 : array_update_80573[8];
  assign array_update_80586[9] = add_80123 == 32'h0000_0009 ? array_update_80584 : array_update_80573[9];
  assign array_index_80588 = array_update_72021[add_80585 > 32'h0000_0009 ? 4'h9 : add_80585[3:0]];
  assign array_index_80589 = array_update_80586[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_80593 = smul32b_32b_x_32b(array_index_80130[add_80585 > 32'h0000_0009 ? 4'h9 : add_80585[3:0]], array_index_80588[add_80531 > 32'h0000_0009 ? 4'h9 : add_80531[3:0]]);
  assign add_80595 = array_index_80589[add_80531 > 32'h0000_0009 ? 4'h9 : add_80531[3:0]] + smul_80593;
  assign array_update_80597[0] = add_80531 == 32'h0000_0000 ? add_80595 : array_index_80589[0];
  assign array_update_80597[1] = add_80531 == 32'h0000_0001 ? add_80595 : array_index_80589[1];
  assign array_update_80597[2] = add_80531 == 32'h0000_0002 ? add_80595 : array_index_80589[2];
  assign array_update_80597[3] = add_80531 == 32'h0000_0003 ? add_80595 : array_index_80589[3];
  assign array_update_80597[4] = add_80531 == 32'h0000_0004 ? add_80595 : array_index_80589[4];
  assign array_update_80597[5] = add_80531 == 32'h0000_0005 ? add_80595 : array_index_80589[5];
  assign array_update_80597[6] = add_80531 == 32'h0000_0006 ? add_80595 : array_index_80589[6];
  assign array_update_80597[7] = add_80531 == 32'h0000_0007 ? add_80595 : array_index_80589[7];
  assign array_update_80597[8] = add_80531 == 32'h0000_0008 ? add_80595 : array_index_80589[8];
  assign array_update_80597[9] = add_80531 == 32'h0000_0009 ? add_80595 : array_index_80589[9];
  assign add_80598 = add_80585 + 32'h0000_0001;
  assign array_update_80599[0] = add_80123 == 32'h0000_0000 ? array_update_80597 : array_update_80586[0];
  assign array_update_80599[1] = add_80123 == 32'h0000_0001 ? array_update_80597 : array_update_80586[1];
  assign array_update_80599[2] = add_80123 == 32'h0000_0002 ? array_update_80597 : array_update_80586[2];
  assign array_update_80599[3] = add_80123 == 32'h0000_0003 ? array_update_80597 : array_update_80586[3];
  assign array_update_80599[4] = add_80123 == 32'h0000_0004 ? array_update_80597 : array_update_80586[4];
  assign array_update_80599[5] = add_80123 == 32'h0000_0005 ? array_update_80597 : array_update_80586[5];
  assign array_update_80599[6] = add_80123 == 32'h0000_0006 ? array_update_80597 : array_update_80586[6];
  assign array_update_80599[7] = add_80123 == 32'h0000_0007 ? array_update_80597 : array_update_80586[7];
  assign array_update_80599[8] = add_80123 == 32'h0000_0008 ? array_update_80597 : array_update_80586[8];
  assign array_update_80599[9] = add_80123 == 32'h0000_0009 ? array_update_80597 : array_update_80586[9];
  assign array_index_80601 = array_update_72021[add_80598 > 32'h0000_0009 ? 4'h9 : add_80598[3:0]];
  assign array_index_80602 = array_update_80599[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_80606 = smul32b_32b_x_32b(array_index_80130[add_80598 > 32'h0000_0009 ? 4'h9 : add_80598[3:0]], array_index_80601[add_80531 > 32'h0000_0009 ? 4'h9 : add_80531[3:0]]);
  assign add_80608 = array_index_80602[add_80531 > 32'h0000_0009 ? 4'h9 : add_80531[3:0]] + smul_80606;
  assign array_update_80610[0] = add_80531 == 32'h0000_0000 ? add_80608 : array_index_80602[0];
  assign array_update_80610[1] = add_80531 == 32'h0000_0001 ? add_80608 : array_index_80602[1];
  assign array_update_80610[2] = add_80531 == 32'h0000_0002 ? add_80608 : array_index_80602[2];
  assign array_update_80610[3] = add_80531 == 32'h0000_0003 ? add_80608 : array_index_80602[3];
  assign array_update_80610[4] = add_80531 == 32'h0000_0004 ? add_80608 : array_index_80602[4];
  assign array_update_80610[5] = add_80531 == 32'h0000_0005 ? add_80608 : array_index_80602[5];
  assign array_update_80610[6] = add_80531 == 32'h0000_0006 ? add_80608 : array_index_80602[6];
  assign array_update_80610[7] = add_80531 == 32'h0000_0007 ? add_80608 : array_index_80602[7];
  assign array_update_80610[8] = add_80531 == 32'h0000_0008 ? add_80608 : array_index_80602[8];
  assign array_update_80610[9] = add_80531 == 32'h0000_0009 ? add_80608 : array_index_80602[9];
  assign add_80611 = add_80598 + 32'h0000_0001;
  assign array_update_80612[0] = add_80123 == 32'h0000_0000 ? array_update_80610 : array_update_80599[0];
  assign array_update_80612[1] = add_80123 == 32'h0000_0001 ? array_update_80610 : array_update_80599[1];
  assign array_update_80612[2] = add_80123 == 32'h0000_0002 ? array_update_80610 : array_update_80599[2];
  assign array_update_80612[3] = add_80123 == 32'h0000_0003 ? array_update_80610 : array_update_80599[3];
  assign array_update_80612[4] = add_80123 == 32'h0000_0004 ? array_update_80610 : array_update_80599[4];
  assign array_update_80612[5] = add_80123 == 32'h0000_0005 ? array_update_80610 : array_update_80599[5];
  assign array_update_80612[6] = add_80123 == 32'h0000_0006 ? array_update_80610 : array_update_80599[6];
  assign array_update_80612[7] = add_80123 == 32'h0000_0007 ? array_update_80610 : array_update_80599[7];
  assign array_update_80612[8] = add_80123 == 32'h0000_0008 ? array_update_80610 : array_update_80599[8];
  assign array_update_80612[9] = add_80123 == 32'h0000_0009 ? array_update_80610 : array_update_80599[9];
  assign array_index_80614 = array_update_72021[add_80611 > 32'h0000_0009 ? 4'h9 : add_80611[3:0]];
  assign array_index_80615 = array_update_80612[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_80619 = smul32b_32b_x_32b(array_index_80130[add_80611 > 32'h0000_0009 ? 4'h9 : add_80611[3:0]], array_index_80614[add_80531 > 32'h0000_0009 ? 4'h9 : add_80531[3:0]]);
  assign add_80621 = array_index_80615[add_80531 > 32'h0000_0009 ? 4'h9 : add_80531[3:0]] + smul_80619;
  assign array_update_80623[0] = add_80531 == 32'h0000_0000 ? add_80621 : array_index_80615[0];
  assign array_update_80623[1] = add_80531 == 32'h0000_0001 ? add_80621 : array_index_80615[1];
  assign array_update_80623[2] = add_80531 == 32'h0000_0002 ? add_80621 : array_index_80615[2];
  assign array_update_80623[3] = add_80531 == 32'h0000_0003 ? add_80621 : array_index_80615[3];
  assign array_update_80623[4] = add_80531 == 32'h0000_0004 ? add_80621 : array_index_80615[4];
  assign array_update_80623[5] = add_80531 == 32'h0000_0005 ? add_80621 : array_index_80615[5];
  assign array_update_80623[6] = add_80531 == 32'h0000_0006 ? add_80621 : array_index_80615[6];
  assign array_update_80623[7] = add_80531 == 32'h0000_0007 ? add_80621 : array_index_80615[7];
  assign array_update_80623[8] = add_80531 == 32'h0000_0008 ? add_80621 : array_index_80615[8];
  assign array_update_80623[9] = add_80531 == 32'h0000_0009 ? add_80621 : array_index_80615[9];
  assign add_80624 = add_80611 + 32'h0000_0001;
  assign array_update_80625[0] = add_80123 == 32'h0000_0000 ? array_update_80623 : array_update_80612[0];
  assign array_update_80625[1] = add_80123 == 32'h0000_0001 ? array_update_80623 : array_update_80612[1];
  assign array_update_80625[2] = add_80123 == 32'h0000_0002 ? array_update_80623 : array_update_80612[2];
  assign array_update_80625[3] = add_80123 == 32'h0000_0003 ? array_update_80623 : array_update_80612[3];
  assign array_update_80625[4] = add_80123 == 32'h0000_0004 ? array_update_80623 : array_update_80612[4];
  assign array_update_80625[5] = add_80123 == 32'h0000_0005 ? array_update_80623 : array_update_80612[5];
  assign array_update_80625[6] = add_80123 == 32'h0000_0006 ? array_update_80623 : array_update_80612[6];
  assign array_update_80625[7] = add_80123 == 32'h0000_0007 ? array_update_80623 : array_update_80612[7];
  assign array_update_80625[8] = add_80123 == 32'h0000_0008 ? array_update_80623 : array_update_80612[8];
  assign array_update_80625[9] = add_80123 == 32'h0000_0009 ? array_update_80623 : array_update_80612[9];
  assign array_index_80627 = array_update_72021[add_80624 > 32'h0000_0009 ? 4'h9 : add_80624[3:0]];
  assign array_index_80628 = array_update_80625[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_80632 = smul32b_32b_x_32b(array_index_80130[add_80624 > 32'h0000_0009 ? 4'h9 : add_80624[3:0]], array_index_80627[add_80531 > 32'h0000_0009 ? 4'h9 : add_80531[3:0]]);
  assign add_80634 = array_index_80628[add_80531 > 32'h0000_0009 ? 4'h9 : add_80531[3:0]] + smul_80632;
  assign array_update_80636[0] = add_80531 == 32'h0000_0000 ? add_80634 : array_index_80628[0];
  assign array_update_80636[1] = add_80531 == 32'h0000_0001 ? add_80634 : array_index_80628[1];
  assign array_update_80636[2] = add_80531 == 32'h0000_0002 ? add_80634 : array_index_80628[2];
  assign array_update_80636[3] = add_80531 == 32'h0000_0003 ? add_80634 : array_index_80628[3];
  assign array_update_80636[4] = add_80531 == 32'h0000_0004 ? add_80634 : array_index_80628[4];
  assign array_update_80636[5] = add_80531 == 32'h0000_0005 ? add_80634 : array_index_80628[5];
  assign array_update_80636[6] = add_80531 == 32'h0000_0006 ? add_80634 : array_index_80628[6];
  assign array_update_80636[7] = add_80531 == 32'h0000_0007 ? add_80634 : array_index_80628[7];
  assign array_update_80636[8] = add_80531 == 32'h0000_0008 ? add_80634 : array_index_80628[8];
  assign array_update_80636[9] = add_80531 == 32'h0000_0009 ? add_80634 : array_index_80628[9];
  assign add_80637 = add_80624 + 32'h0000_0001;
  assign array_update_80638[0] = add_80123 == 32'h0000_0000 ? array_update_80636 : array_update_80625[0];
  assign array_update_80638[1] = add_80123 == 32'h0000_0001 ? array_update_80636 : array_update_80625[1];
  assign array_update_80638[2] = add_80123 == 32'h0000_0002 ? array_update_80636 : array_update_80625[2];
  assign array_update_80638[3] = add_80123 == 32'h0000_0003 ? array_update_80636 : array_update_80625[3];
  assign array_update_80638[4] = add_80123 == 32'h0000_0004 ? array_update_80636 : array_update_80625[4];
  assign array_update_80638[5] = add_80123 == 32'h0000_0005 ? array_update_80636 : array_update_80625[5];
  assign array_update_80638[6] = add_80123 == 32'h0000_0006 ? array_update_80636 : array_update_80625[6];
  assign array_update_80638[7] = add_80123 == 32'h0000_0007 ? array_update_80636 : array_update_80625[7];
  assign array_update_80638[8] = add_80123 == 32'h0000_0008 ? array_update_80636 : array_update_80625[8];
  assign array_update_80638[9] = add_80123 == 32'h0000_0009 ? array_update_80636 : array_update_80625[9];
  assign array_index_80640 = array_update_72021[add_80637 > 32'h0000_0009 ? 4'h9 : add_80637[3:0]];
  assign array_index_80641 = array_update_80638[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_80645 = smul32b_32b_x_32b(array_index_80130[add_80637 > 32'h0000_0009 ? 4'h9 : add_80637[3:0]], array_index_80640[add_80531 > 32'h0000_0009 ? 4'h9 : add_80531[3:0]]);
  assign add_80647 = array_index_80641[add_80531 > 32'h0000_0009 ? 4'h9 : add_80531[3:0]] + smul_80645;
  assign array_update_80649[0] = add_80531 == 32'h0000_0000 ? add_80647 : array_index_80641[0];
  assign array_update_80649[1] = add_80531 == 32'h0000_0001 ? add_80647 : array_index_80641[1];
  assign array_update_80649[2] = add_80531 == 32'h0000_0002 ? add_80647 : array_index_80641[2];
  assign array_update_80649[3] = add_80531 == 32'h0000_0003 ? add_80647 : array_index_80641[3];
  assign array_update_80649[4] = add_80531 == 32'h0000_0004 ? add_80647 : array_index_80641[4];
  assign array_update_80649[5] = add_80531 == 32'h0000_0005 ? add_80647 : array_index_80641[5];
  assign array_update_80649[6] = add_80531 == 32'h0000_0006 ? add_80647 : array_index_80641[6];
  assign array_update_80649[7] = add_80531 == 32'h0000_0007 ? add_80647 : array_index_80641[7];
  assign array_update_80649[8] = add_80531 == 32'h0000_0008 ? add_80647 : array_index_80641[8];
  assign array_update_80649[9] = add_80531 == 32'h0000_0009 ? add_80647 : array_index_80641[9];
  assign add_80650 = add_80637 + 32'h0000_0001;
  assign array_update_80651[0] = add_80123 == 32'h0000_0000 ? array_update_80649 : array_update_80638[0];
  assign array_update_80651[1] = add_80123 == 32'h0000_0001 ? array_update_80649 : array_update_80638[1];
  assign array_update_80651[2] = add_80123 == 32'h0000_0002 ? array_update_80649 : array_update_80638[2];
  assign array_update_80651[3] = add_80123 == 32'h0000_0003 ? array_update_80649 : array_update_80638[3];
  assign array_update_80651[4] = add_80123 == 32'h0000_0004 ? array_update_80649 : array_update_80638[4];
  assign array_update_80651[5] = add_80123 == 32'h0000_0005 ? array_update_80649 : array_update_80638[5];
  assign array_update_80651[6] = add_80123 == 32'h0000_0006 ? array_update_80649 : array_update_80638[6];
  assign array_update_80651[7] = add_80123 == 32'h0000_0007 ? array_update_80649 : array_update_80638[7];
  assign array_update_80651[8] = add_80123 == 32'h0000_0008 ? array_update_80649 : array_update_80638[8];
  assign array_update_80651[9] = add_80123 == 32'h0000_0009 ? array_update_80649 : array_update_80638[9];
  assign array_index_80653 = array_update_72021[add_80650 > 32'h0000_0009 ? 4'h9 : add_80650[3:0]];
  assign array_index_80654 = array_update_80651[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_80658 = smul32b_32b_x_32b(array_index_80130[add_80650 > 32'h0000_0009 ? 4'h9 : add_80650[3:0]], array_index_80653[add_80531 > 32'h0000_0009 ? 4'h9 : add_80531[3:0]]);
  assign add_80660 = array_index_80654[add_80531 > 32'h0000_0009 ? 4'h9 : add_80531[3:0]] + smul_80658;
  assign array_update_80661[0] = add_80531 == 32'h0000_0000 ? add_80660 : array_index_80654[0];
  assign array_update_80661[1] = add_80531 == 32'h0000_0001 ? add_80660 : array_index_80654[1];
  assign array_update_80661[2] = add_80531 == 32'h0000_0002 ? add_80660 : array_index_80654[2];
  assign array_update_80661[3] = add_80531 == 32'h0000_0003 ? add_80660 : array_index_80654[3];
  assign array_update_80661[4] = add_80531 == 32'h0000_0004 ? add_80660 : array_index_80654[4];
  assign array_update_80661[5] = add_80531 == 32'h0000_0005 ? add_80660 : array_index_80654[5];
  assign array_update_80661[6] = add_80531 == 32'h0000_0006 ? add_80660 : array_index_80654[6];
  assign array_update_80661[7] = add_80531 == 32'h0000_0007 ? add_80660 : array_index_80654[7];
  assign array_update_80661[8] = add_80531 == 32'h0000_0008 ? add_80660 : array_index_80654[8];
  assign array_update_80661[9] = add_80531 == 32'h0000_0009 ? add_80660 : array_index_80654[9];
  assign array_update_80662[0] = add_80123 == 32'h0000_0000 ? array_update_80661 : array_update_80651[0];
  assign array_update_80662[1] = add_80123 == 32'h0000_0001 ? array_update_80661 : array_update_80651[1];
  assign array_update_80662[2] = add_80123 == 32'h0000_0002 ? array_update_80661 : array_update_80651[2];
  assign array_update_80662[3] = add_80123 == 32'h0000_0003 ? array_update_80661 : array_update_80651[3];
  assign array_update_80662[4] = add_80123 == 32'h0000_0004 ? array_update_80661 : array_update_80651[4];
  assign array_update_80662[5] = add_80123 == 32'h0000_0005 ? array_update_80661 : array_update_80651[5];
  assign array_update_80662[6] = add_80123 == 32'h0000_0006 ? array_update_80661 : array_update_80651[6];
  assign array_update_80662[7] = add_80123 == 32'h0000_0007 ? array_update_80661 : array_update_80651[7];
  assign array_update_80662[8] = add_80123 == 32'h0000_0008 ? array_update_80661 : array_update_80651[8];
  assign array_update_80662[9] = add_80123 == 32'h0000_0009 ? array_update_80661 : array_update_80651[9];
  assign array_index_80664 = array_update_80662[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign add_80666 = add_80531 + 32'h0000_0001;
  assign array_update_80667[0] = add_80666 == 32'h0000_0000 ? 32'h0000_0000 : array_index_80664[0];
  assign array_update_80667[1] = add_80666 == 32'h0000_0001 ? 32'h0000_0000 : array_index_80664[1];
  assign array_update_80667[2] = add_80666 == 32'h0000_0002 ? 32'h0000_0000 : array_index_80664[2];
  assign array_update_80667[3] = add_80666 == 32'h0000_0003 ? 32'h0000_0000 : array_index_80664[3];
  assign array_update_80667[4] = add_80666 == 32'h0000_0004 ? 32'h0000_0000 : array_index_80664[4];
  assign array_update_80667[5] = add_80666 == 32'h0000_0005 ? 32'h0000_0000 : array_index_80664[5];
  assign array_update_80667[6] = add_80666 == 32'h0000_0006 ? 32'h0000_0000 : array_index_80664[6];
  assign array_update_80667[7] = add_80666 == 32'h0000_0007 ? 32'h0000_0000 : array_index_80664[7];
  assign array_update_80667[8] = add_80666 == 32'h0000_0008 ? 32'h0000_0000 : array_index_80664[8];
  assign array_update_80667[9] = add_80666 == 32'h0000_0009 ? 32'h0000_0000 : array_index_80664[9];
  assign literal_80668 = 32'h0000_0000;
  assign array_update_80669[0] = add_80123 == 32'h0000_0000 ? array_update_80667 : array_update_80662[0];
  assign array_update_80669[1] = add_80123 == 32'h0000_0001 ? array_update_80667 : array_update_80662[1];
  assign array_update_80669[2] = add_80123 == 32'h0000_0002 ? array_update_80667 : array_update_80662[2];
  assign array_update_80669[3] = add_80123 == 32'h0000_0003 ? array_update_80667 : array_update_80662[3];
  assign array_update_80669[4] = add_80123 == 32'h0000_0004 ? array_update_80667 : array_update_80662[4];
  assign array_update_80669[5] = add_80123 == 32'h0000_0005 ? array_update_80667 : array_update_80662[5];
  assign array_update_80669[6] = add_80123 == 32'h0000_0006 ? array_update_80667 : array_update_80662[6];
  assign array_update_80669[7] = add_80123 == 32'h0000_0007 ? array_update_80667 : array_update_80662[7];
  assign array_update_80669[8] = add_80123 == 32'h0000_0008 ? array_update_80667 : array_update_80662[8];
  assign array_update_80669[9] = add_80123 == 32'h0000_0009 ? array_update_80667 : array_update_80662[9];
  assign array_index_80671 = array_update_72021[literal_80668 > 32'h0000_0009 ? 4'h9 : literal_80668[3:0]];
  assign array_index_80672 = array_update_80669[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_80676 = smul32b_32b_x_32b(array_index_80130[literal_80668 > 32'h0000_0009 ? 4'h9 : literal_80668[3:0]], array_index_80671[add_80666 > 32'h0000_0009 ? 4'h9 : add_80666[3:0]]);
  assign add_80678 = array_index_80672[add_80666 > 32'h0000_0009 ? 4'h9 : add_80666[3:0]] + smul_80676;
  assign array_update_80680[0] = add_80666 == 32'h0000_0000 ? add_80678 : array_index_80672[0];
  assign array_update_80680[1] = add_80666 == 32'h0000_0001 ? add_80678 : array_index_80672[1];
  assign array_update_80680[2] = add_80666 == 32'h0000_0002 ? add_80678 : array_index_80672[2];
  assign array_update_80680[3] = add_80666 == 32'h0000_0003 ? add_80678 : array_index_80672[3];
  assign array_update_80680[4] = add_80666 == 32'h0000_0004 ? add_80678 : array_index_80672[4];
  assign array_update_80680[5] = add_80666 == 32'h0000_0005 ? add_80678 : array_index_80672[5];
  assign array_update_80680[6] = add_80666 == 32'h0000_0006 ? add_80678 : array_index_80672[6];
  assign array_update_80680[7] = add_80666 == 32'h0000_0007 ? add_80678 : array_index_80672[7];
  assign array_update_80680[8] = add_80666 == 32'h0000_0008 ? add_80678 : array_index_80672[8];
  assign array_update_80680[9] = add_80666 == 32'h0000_0009 ? add_80678 : array_index_80672[9];
  assign add_80681 = literal_80668 + 32'h0000_0001;
  assign array_update_80682[0] = add_80123 == 32'h0000_0000 ? array_update_80680 : array_update_80669[0];
  assign array_update_80682[1] = add_80123 == 32'h0000_0001 ? array_update_80680 : array_update_80669[1];
  assign array_update_80682[2] = add_80123 == 32'h0000_0002 ? array_update_80680 : array_update_80669[2];
  assign array_update_80682[3] = add_80123 == 32'h0000_0003 ? array_update_80680 : array_update_80669[3];
  assign array_update_80682[4] = add_80123 == 32'h0000_0004 ? array_update_80680 : array_update_80669[4];
  assign array_update_80682[5] = add_80123 == 32'h0000_0005 ? array_update_80680 : array_update_80669[5];
  assign array_update_80682[6] = add_80123 == 32'h0000_0006 ? array_update_80680 : array_update_80669[6];
  assign array_update_80682[7] = add_80123 == 32'h0000_0007 ? array_update_80680 : array_update_80669[7];
  assign array_update_80682[8] = add_80123 == 32'h0000_0008 ? array_update_80680 : array_update_80669[8];
  assign array_update_80682[9] = add_80123 == 32'h0000_0009 ? array_update_80680 : array_update_80669[9];
  assign array_index_80684 = array_update_72021[add_80681 > 32'h0000_0009 ? 4'h9 : add_80681[3:0]];
  assign array_index_80685 = array_update_80682[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_80689 = smul32b_32b_x_32b(array_index_80130[add_80681 > 32'h0000_0009 ? 4'h9 : add_80681[3:0]], array_index_80684[add_80666 > 32'h0000_0009 ? 4'h9 : add_80666[3:0]]);
  assign add_80691 = array_index_80685[add_80666 > 32'h0000_0009 ? 4'h9 : add_80666[3:0]] + smul_80689;
  assign array_update_80693[0] = add_80666 == 32'h0000_0000 ? add_80691 : array_index_80685[0];
  assign array_update_80693[1] = add_80666 == 32'h0000_0001 ? add_80691 : array_index_80685[1];
  assign array_update_80693[2] = add_80666 == 32'h0000_0002 ? add_80691 : array_index_80685[2];
  assign array_update_80693[3] = add_80666 == 32'h0000_0003 ? add_80691 : array_index_80685[3];
  assign array_update_80693[4] = add_80666 == 32'h0000_0004 ? add_80691 : array_index_80685[4];
  assign array_update_80693[5] = add_80666 == 32'h0000_0005 ? add_80691 : array_index_80685[5];
  assign array_update_80693[6] = add_80666 == 32'h0000_0006 ? add_80691 : array_index_80685[6];
  assign array_update_80693[7] = add_80666 == 32'h0000_0007 ? add_80691 : array_index_80685[7];
  assign array_update_80693[8] = add_80666 == 32'h0000_0008 ? add_80691 : array_index_80685[8];
  assign array_update_80693[9] = add_80666 == 32'h0000_0009 ? add_80691 : array_index_80685[9];
  assign add_80694 = add_80681 + 32'h0000_0001;
  assign array_update_80695[0] = add_80123 == 32'h0000_0000 ? array_update_80693 : array_update_80682[0];
  assign array_update_80695[1] = add_80123 == 32'h0000_0001 ? array_update_80693 : array_update_80682[1];
  assign array_update_80695[2] = add_80123 == 32'h0000_0002 ? array_update_80693 : array_update_80682[2];
  assign array_update_80695[3] = add_80123 == 32'h0000_0003 ? array_update_80693 : array_update_80682[3];
  assign array_update_80695[4] = add_80123 == 32'h0000_0004 ? array_update_80693 : array_update_80682[4];
  assign array_update_80695[5] = add_80123 == 32'h0000_0005 ? array_update_80693 : array_update_80682[5];
  assign array_update_80695[6] = add_80123 == 32'h0000_0006 ? array_update_80693 : array_update_80682[6];
  assign array_update_80695[7] = add_80123 == 32'h0000_0007 ? array_update_80693 : array_update_80682[7];
  assign array_update_80695[8] = add_80123 == 32'h0000_0008 ? array_update_80693 : array_update_80682[8];
  assign array_update_80695[9] = add_80123 == 32'h0000_0009 ? array_update_80693 : array_update_80682[9];
  assign array_index_80697 = array_update_72021[add_80694 > 32'h0000_0009 ? 4'h9 : add_80694[3:0]];
  assign array_index_80698 = array_update_80695[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_80702 = smul32b_32b_x_32b(array_index_80130[add_80694 > 32'h0000_0009 ? 4'h9 : add_80694[3:0]], array_index_80697[add_80666 > 32'h0000_0009 ? 4'h9 : add_80666[3:0]]);
  assign add_80704 = array_index_80698[add_80666 > 32'h0000_0009 ? 4'h9 : add_80666[3:0]] + smul_80702;
  assign array_update_80706[0] = add_80666 == 32'h0000_0000 ? add_80704 : array_index_80698[0];
  assign array_update_80706[1] = add_80666 == 32'h0000_0001 ? add_80704 : array_index_80698[1];
  assign array_update_80706[2] = add_80666 == 32'h0000_0002 ? add_80704 : array_index_80698[2];
  assign array_update_80706[3] = add_80666 == 32'h0000_0003 ? add_80704 : array_index_80698[3];
  assign array_update_80706[4] = add_80666 == 32'h0000_0004 ? add_80704 : array_index_80698[4];
  assign array_update_80706[5] = add_80666 == 32'h0000_0005 ? add_80704 : array_index_80698[5];
  assign array_update_80706[6] = add_80666 == 32'h0000_0006 ? add_80704 : array_index_80698[6];
  assign array_update_80706[7] = add_80666 == 32'h0000_0007 ? add_80704 : array_index_80698[7];
  assign array_update_80706[8] = add_80666 == 32'h0000_0008 ? add_80704 : array_index_80698[8];
  assign array_update_80706[9] = add_80666 == 32'h0000_0009 ? add_80704 : array_index_80698[9];
  assign add_80707 = add_80694 + 32'h0000_0001;
  assign array_update_80708[0] = add_80123 == 32'h0000_0000 ? array_update_80706 : array_update_80695[0];
  assign array_update_80708[1] = add_80123 == 32'h0000_0001 ? array_update_80706 : array_update_80695[1];
  assign array_update_80708[2] = add_80123 == 32'h0000_0002 ? array_update_80706 : array_update_80695[2];
  assign array_update_80708[3] = add_80123 == 32'h0000_0003 ? array_update_80706 : array_update_80695[3];
  assign array_update_80708[4] = add_80123 == 32'h0000_0004 ? array_update_80706 : array_update_80695[4];
  assign array_update_80708[5] = add_80123 == 32'h0000_0005 ? array_update_80706 : array_update_80695[5];
  assign array_update_80708[6] = add_80123 == 32'h0000_0006 ? array_update_80706 : array_update_80695[6];
  assign array_update_80708[7] = add_80123 == 32'h0000_0007 ? array_update_80706 : array_update_80695[7];
  assign array_update_80708[8] = add_80123 == 32'h0000_0008 ? array_update_80706 : array_update_80695[8];
  assign array_update_80708[9] = add_80123 == 32'h0000_0009 ? array_update_80706 : array_update_80695[9];
  assign array_index_80710 = array_update_72021[add_80707 > 32'h0000_0009 ? 4'h9 : add_80707[3:0]];
  assign array_index_80711 = array_update_80708[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_80715 = smul32b_32b_x_32b(array_index_80130[add_80707 > 32'h0000_0009 ? 4'h9 : add_80707[3:0]], array_index_80710[add_80666 > 32'h0000_0009 ? 4'h9 : add_80666[3:0]]);
  assign add_80717 = array_index_80711[add_80666 > 32'h0000_0009 ? 4'h9 : add_80666[3:0]] + smul_80715;
  assign array_update_80719[0] = add_80666 == 32'h0000_0000 ? add_80717 : array_index_80711[0];
  assign array_update_80719[1] = add_80666 == 32'h0000_0001 ? add_80717 : array_index_80711[1];
  assign array_update_80719[2] = add_80666 == 32'h0000_0002 ? add_80717 : array_index_80711[2];
  assign array_update_80719[3] = add_80666 == 32'h0000_0003 ? add_80717 : array_index_80711[3];
  assign array_update_80719[4] = add_80666 == 32'h0000_0004 ? add_80717 : array_index_80711[4];
  assign array_update_80719[5] = add_80666 == 32'h0000_0005 ? add_80717 : array_index_80711[5];
  assign array_update_80719[6] = add_80666 == 32'h0000_0006 ? add_80717 : array_index_80711[6];
  assign array_update_80719[7] = add_80666 == 32'h0000_0007 ? add_80717 : array_index_80711[7];
  assign array_update_80719[8] = add_80666 == 32'h0000_0008 ? add_80717 : array_index_80711[8];
  assign array_update_80719[9] = add_80666 == 32'h0000_0009 ? add_80717 : array_index_80711[9];
  assign add_80720 = add_80707 + 32'h0000_0001;
  assign array_update_80721[0] = add_80123 == 32'h0000_0000 ? array_update_80719 : array_update_80708[0];
  assign array_update_80721[1] = add_80123 == 32'h0000_0001 ? array_update_80719 : array_update_80708[1];
  assign array_update_80721[2] = add_80123 == 32'h0000_0002 ? array_update_80719 : array_update_80708[2];
  assign array_update_80721[3] = add_80123 == 32'h0000_0003 ? array_update_80719 : array_update_80708[3];
  assign array_update_80721[4] = add_80123 == 32'h0000_0004 ? array_update_80719 : array_update_80708[4];
  assign array_update_80721[5] = add_80123 == 32'h0000_0005 ? array_update_80719 : array_update_80708[5];
  assign array_update_80721[6] = add_80123 == 32'h0000_0006 ? array_update_80719 : array_update_80708[6];
  assign array_update_80721[7] = add_80123 == 32'h0000_0007 ? array_update_80719 : array_update_80708[7];
  assign array_update_80721[8] = add_80123 == 32'h0000_0008 ? array_update_80719 : array_update_80708[8];
  assign array_update_80721[9] = add_80123 == 32'h0000_0009 ? array_update_80719 : array_update_80708[9];
  assign array_index_80723 = array_update_72021[add_80720 > 32'h0000_0009 ? 4'h9 : add_80720[3:0]];
  assign array_index_80724 = array_update_80721[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_80728 = smul32b_32b_x_32b(array_index_80130[add_80720 > 32'h0000_0009 ? 4'h9 : add_80720[3:0]], array_index_80723[add_80666 > 32'h0000_0009 ? 4'h9 : add_80666[3:0]]);
  assign add_80730 = array_index_80724[add_80666 > 32'h0000_0009 ? 4'h9 : add_80666[3:0]] + smul_80728;
  assign array_update_80732[0] = add_80666 == 32'h0000_0000 ? add_80730 : array_index_80724[0];
  assign array_update_80732[1] = add_80666 == 32'h0000_0001 ? add_80730 : array_index_80724[1];
  assign array_update_80732[2] = add_80666 == 32'h0000_0002 ? add_80730 : array_index_80724[2];
  assign array_update_80732[3] = add_80666 == 32'h0000_0003 ? add_80730 : array_index_80724[3];
  assign array_update_80732[4] = add_80666 == 32'h0000_0004 ? add_80730 : array_index_80724[4];
  assign array_update_80732[5] = add_80666 == 32'h0000_0005 ? add_80730 : array_index_80724[5];
  assign array_update_80732[6] = add_80666 == 32'h0000_0006 ? add_80730 : array_index_80724[6];
  assign array_update_80732[7] = add_80666 == 32'h0000_0007 ? add_80730 : array_index_80724[7];
  assign array_update_80732[8] = add_80666 == 32'h0000_0008 ? add_80730 : array_index_80724[8];
  assign array_update_80732[9] = add_80666 == 32'h0000_0009 ? add_80730 : array_index_80724[9];
  assign add_80733 = add_80720 + 32'h0000_0001;
  assign array_update_80734[0] = add_80123 == 32'h0000_0000 ? array_update_80732 : array_update_80721[0];
  assign array_update_80734[1] = add_80123 == 32'h0000_0001 ? array_update_80732 : array_update_80721[1];
  assign array_update_80734[2] = add_80123 == 32'h0000_0002 ? array_update_80732 : array_update_80721[2];
  assign array_update_80734[3] = add_80123 == 32'h0000_0003 ? array_update_80732 : array_update_80721[3];
  assign array_update_80734[4] = add_80123 == 32'h0000_0004 ? array_update_80732 : array_update_80721[4];
  assign array_update_80734[5] = add_80123 == 32'h0000_0005 ? array_update_80732 : array_update_80721[5];
  assign array_update_80734[6] = add_80123 == 32'h0000_0006 ? array_update_80732 : array_update_80721[6];
  assign array_update_80734[7] = add_80123 == 32'h0000_0007 ? array_update_80732 : array_update_80721[7];
  assign array_update_80734[8] = add_80123 == 32'h0000_0008 ? array_update_80732 : array_update_80721[8];
  assign array_update_80734[9] = add_80123 == 32'h0000_0009 ? array_update_80732 : array_update_80721[9];
  assign array_index_80736 = array_update_72021[add_80733 > 32'h0000_0009 ? 4'h9 : add_80733[3:0]];
  assign array_index_80737 = array_update_80734[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_80741 = smul32b_32b_x_32b(array_index_80130[add_80733 > 32'h0000_0009 ? 4'h9 : add_80733[3:0]], array_index_80736[add_80666 > 32'h0000_0009 ? 4'h9 : add_80666[3:0]]);
  assign add_80743 = array_index_80737[add_80666 > 32'h0000_0009 ? 4'h9 : add_80666[3:0]] + smul_80741;
  assign array_update_80745[0] = add_80666 == 32'h0000_0000 ? add_80743 : array_index_80737[0];
  assign array_update_80745[1] = add_80666 == 32'h0000_0001 ? add_80743 : array_index_80737[1];
  assign array_update_80745[2] = add_80666 == 32'h0000_0002 ? add_80743 : array_index_80737[2];
  assign array_update_80745[3] = add_80666 == 32'h0000_0003 ? add_80743 : array_index_80737[3];
  assign array_update_80745[4] = add_80666 == 32'h0000_0004 ? add_80743 : array_index_80737[4];
  assign array_update_80745[5] = add_80666 == 32'h0000_0005 ? add_80743 : array_index_80737[5];
  assign array_update_80745[6] = add_80666 == 32'h0000_0006 ? add_80743 : array_index_80737[6];
  assign array_update_80745[7] = add_80666 == 32'h0000_0007 ? add_80743 : array_index_80737[7];
  assign array_update_80745[8] = add_80666 == 32'h0000_0008 ? add_80743 : array_index_80737[8];
  assign array_update_80745[9] = add_80666 == 32'h0000_0009 ? add_80743 : array_index_80737[9];
  assign add_80746 = add_80733 + 32'h0000_0001;
  assign array_update_80747[0] = add_80123 == 32'h0000_0000 ? array_update_80745 : array_update_80734[0];
  assign array_update_80747[1] = add_80123 == 32'h0000_0001 ? array_update_80745 : array_update_80734[1];
  assign array_update_80747[2] = add_80123 == 32'h0000_0002 ? array_update_80745 : array_update_80734[2];
  assign array_update_80747[3] = add_80123 == 32'h0000_0003 ? array_update_80745 : array_update_80734[3];
  assign array_update_80747[4] = add_80123 == 32'h0000_0004 ? array_update_80745 : array_update_80734[4];
  assign array_update_80747[5] = add_80123 == 32'h0000_0005 ? array_update_80745 : array_update_80734[5];
  assign array_update_80747[6] = add_80123 == 32'h0000_0006 ? array_update_80745 : array_update_80734[6];
  assign array_update_80747[7] = add_80123 == 32'h0000_0007 ? array_update_80745 : array_update_80734[7];
  assign array_update_80747[8] = add_80123 == 32'h0000_0008 ? array_update_80745 : array_update_80734[8];
  assign array_update_80747[9] = add_80123 == 32'h0000_0009 ? array_update_80745 : array_update_80734[9];
  assign array_index_80749 = array_update_72021[add_80746 > 32'h0000_0009 ? 4'h9 : add_80746[3:0]];
  assign array_index_80750 = array_update_80747[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_80754 = smul32b_32b_x_32b(array_index_80130[add_80746 > 32'h0000_0009 ? 4'h9 : add_80746[3:0]], array_index_80749[add_80666 > 32'h0000_0009 ? 4'h9 : add_80666[3:0]]);
  assign add_80756 = array_index_80750[add_80666 > 32'h0000_0009 ? 4'h9 : add_80666[3:0]] + smul_80754;
  assign array_update_80758[0] = add_80666 == 32'h0000_0000 ? add_80756 : array_index_80750[0];
  assign array_update_80758[1] = add_80666 == 32'h0000_0001 ? add_80756 : array_index_80750[1];
  assign array_update_80758[2] = add_80666 == 32'h0000_0002 ? add_80756 : array_index_80750[2];
  assign array_update_80758[3] = add_80666 == 32'h0000_0003 ? add_80756 : array_index_80750[3];
  assign array_update_80758[4] = add_80666 == 32'h0000_0004 ? add_80756 : array_index_80750[4];
  assign array_update_80758[5] = add_80666 == 32'h0000_0005 ? add_80756 : array_index_80750[5];
  assign array_update_80758[6] = add_80666 == 32'h0000_0006 ? add_80756 : array_index_80750[6];
  assign array_update_80758[7] = add_80666 == 32'h0000_0007 ? add_80756 : array_index_80750[7];
  assign array_update_80758[8] = add_80666 == 32'h0000_0008 ? add_80756 : array_index_80750[8];
  assign array_update_80758[9] = add_80666 == 32'h0000_0009 ? add_80756 : array_index_80750[9];
  assign add_80759 = add_80746 + 32'h0000_0001;
  assign array_update_80760[0] = add_80123 == 32'h0000_0000 ? array_update_80758 : array_update_80747[0];
  assign array_update_80760[1] = add_80123 == 32'h0000_0001 ? array_update_80758 : array_update_80747[1];
  assign array_update_80760[2] = add_80123 == 32'h0000_0002 ? array_update_80758 : array_update_80747[2];
  assign array_update_80760[3] = add_80123 == 32'h0000_0003 ? array_update_80758 : array_update_80747[3];
  assign array_update_80760[4] = add_80123 == 32'h0000_0004 ? array_update_80758 : array_update_80747[4];
  assign array_update_80760[5] = add_80123 == 32'h0000_0005 ? array_update_80758 : array_update_80747[5];
  assign array_update_80760[6] = add_80123 == 32'h0000_0006 ? array_update_80758 : array_update_80747[6];
  assign array_update_80760[7] = add_80123 == 32'h0000_0007 ? array_update_80758 : array_update_80747[7];
  assign array_update_80760[8] = add_80123 == 32'h0000_0008 ? array_update_80758 : array_update_80747[8];
  assign array_update_80760[9] = add_80123 == 32'h0000_0009 ? array_update_80758 : array_update_80747[9];
  assign array_index_80762 = array_update_72021[add_80759 > 32'h0000_0009 ? 4'h9 : add_80759[3:0]];
  assign array_index_80763 = array_update_80760[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_80767 = smul32b_32b_x_32b(array_index_80130[add_80759 > 32'h0000_0009 ? 4'h9 : add_80759[3:0]], array_index_80762[add_80666 > 32'h0000_0009 ? 4'h9 : add_80666[3:0]]);
  assign add_80769 = array_index_80763[add_80666 > 32'h0000_0009 ? 4'h9 : add_80666[3:0]] + smul_80767;
  assign array_update_80771[0] = add_80666 == 32'h0000_0000 ? add_80769 : array_index_80763[0];
  assign array_update_80771[1] = add_80666 == 32'h0000_0001 ? add_80769 : array_index_80763[1];
  assign array_update_80771[2] = add_80666 == 32'h0000_0002 ? add_80769 : array_index_80763[2];
  assign array_update_80771[3] = add_80666 == 32'h0000_0003 ? add_80769 : array_index_80763[3];
  assign array_update_80771[4] = add_80666 == 32'h0000_0004 ? add_80769 : array_index_80763[4];
  assign array_update_80771[5] = add_80666 == 32'h0000_0005 ? add_80769 : array_index_80763[5];
  assign array_update_80771[6] = add_80666 == 32'h0000_0006 ? add_80769 : array_index_80763[6];
  assign array_update_80771[7] = add_80666 == 32'h0000_0007 ? add_80769 : array_index_80763[7];
  assign array_update_80771[8] = add_80666 == 32'h0000_0008 ? add_80769 : array_index_80763[8];
  assign array_update_80771[9] = add_80666 == 32'h0000_0009 ? add_80769 : array_index_80763[9];
  assign add_80772 = add_80759 + 32'h0000_0001;
  assign array_update_80773[0] = add_80123 == 32'h0000_0000 ? array_update_80771 : array_update_80760[0];
  assign array_update_80773[1] = add_80123 == 32'h0000_0001 ? array_update_80771 : array_update_80760[1];
  assign array_update_80773[2] = add_80123 == 32'h0000_0002 ? array_update_80771 : array_update_80760[2];
  assign array_update_80773[3] = add_80123 == 32'h0000_0003 ? array_update_80771 : array_update_80760[3];
  assign array_update_80773[4] = add_80123 == 32'h0000_0004 ? array_update_80771 : array_update_80760[4];
  assign array_update_80773[5] = add_80123 == 32'h0000_0005 ? array_update_80771 : array_update_80760[5];
  assign array_update_80773[6] = add_80123 == 32'h0000_0006 ? array_update_80771 : array_update_80760[6];
  assign array_update_80773[7] = add_80123 == 32'h0000_0007 ? array_update_80771 : array_update_80760[7];
  assign array_update_80773[8] = add_80123 == 32'h0000_0008 ? array_update_80771 : array_update_80760[8];
  assign array_update_80773[9] = add_80123 == 32'h0000_0009 ? array_update_80771 : array_update_80760[9];
  assign array_index_80775 = array_update_72021[add_80772 > 32'h0000_0009 ? 4'h9 : add_80772[3:0]];
  assign array_index_80776 = array_update_80773[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_80780 = smul32b_32b_x_32b(array_index_80130[add_80772 > 32'h0000_0009 ? 4'h9 : add_80772[3:0]], array_index_80775[add_80666 > 32'h0000_0009 ? 4'h9 : add_80666[3:0]]);
  assign add_80782 = array_index_80776[add_80666 > 32'h0000_0009 ? 4'h9 : add_80666[3:0]] + smul_80780;
  assign array_update_80784[0] = add_80666 == 32'h0000_0000 ? add_80782 : array_index_80776[0];
  assign array_update_80784[1] = add_80666 == 32'h0000_0001 ? add_80782 : array_index_80776[1];
  assign array_update_80784[2] = add_80666 == 32'h0000_0002 ? add_80782 : array_index_80776[2];
  assign array_update_80784[3] = add_80666 == 32'h0000_0003 ? add_80782 : array_index_80776[3];
  assign array_update_80784[4] = add_80666 == 32'h0000_0004 ? add_80782 : array_index_80776[4];
  assign array_update_80784[5] = add_80666 == 32'h0000_0005 ? add_80782 : array_index_80776[5];
  assign array_update_80784[6] = add_80666 == 32'h0000_0006 ? add_80782 : array_index_80776[6];
  assign array_update_80784[7] = add_80666 == 32'h0000_0007 ? add_80782 : array_index_80776[7];
  assign array_update_80784[8] = add_80666 == 32'h0000_0008 ? add_80782 : array_index_80776[8];
  assign array_update_80784[9] = add_80666 == 32'h0000_0009 ? add_80782 : array_index_80776[9];
  assign add_80785 = add_80772 + 32'h0000_0001;
  assign array_update_80786[0] = add_80123 == 32'h0000_0000 ? array_update_80784 : array_update_80773[0];
  assign array_update_80786[1] = add_80123 == 32'h0000_0001 ? array_update_80784 : array_update_80773[1];
  assign array_update_80786[2] = add_80123 == 32'h0000_0002 ? array_update_80784 : array_update_80773[2];
  assign array_update_80786[3] = add_80123 == 32'h0000_0003 ? array_update_80784 : array_update_80773[3];
  assign array_update_80786[4] = add_80123 == 32'h0000_0004 ? array_update_80784 : array_update_80773[4];
  assign array_update_80786[5] = add_80123 == 32'h0000_0005 ? array_update_80784 : array_update_80773[5];
  assign array_update_80786[6] = add_80123 == 32'h0000_0006 ? array_update_80784 : array_update_80773[6];
  assign array_update_80786[7] = add_80123 == 32'h0000_0007 ? array_update_80784 : array_update_80773[7];
  assign array_update_80786[8] = add_80123 == 32'h0000_0008 ? array_update_80784 : array_update_80773[8];
  assign array_update_80786[9] = add_80123 == 32'h0000_0009 ? array_update_80784 : array_update_80773[9];
  assign array_index_80788 = array_update_72021[add_80785 > 32'h0000_0009 ? 4'h9 : add_80785[3:0]];
  assign array_index_80789 = array_update_80786[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_80793 = smul32b_32b_x_32b(array_index_80130[add_80785 > 32'h0000_0009 ? 4'h9 : add_80785[3:0]], array_index_80788[add_80666 > 32'h0000_0009 ? 4'h9 : add_80666[3:0]]);
  assign add_80795 = array_index_80789[add_80666 > 32'h0000_0009 ? 4'h9 : add_80666[3:0]] + smul_80793;
  assign array_update_80796[0] = add_80666 == 32'h0000_0000 ? add_80795 : array_index_80789[0];
  assign array_update_80796[1] = add_80666 == 32'h0000_0001 ? add_80795 : array_index_80789[1];
  assign array_update_80796[2] = add_80666 == 32'h0000_0002 ? add_80795 : array_index_80789[2];
  assign array_update_80796[3] = add_80666 == 32'h0000_0003 ? add_80795 : array_index_80789[3];
  assign array_update_80796[4] = add_80666 == 32'h0000_0004 ? add_80795 : array_index_80789[4];
  assign array_update_80796[5] = add_80666 == 32'h0000_0005 ? add_80795 : array_index_80789[5];
  assign array_update_80796[6] = add_80666 == 32'h0000_0006 ? add_80795 : array_index_80789[6];
  assign array_update_80796[7] = add_80666 == 32'h0000_0007 ? add_80795 : array_index_80789[7];
  assign array_update_80796[8] = add_80666 == 32'h0000_0008 ? add_80795 : array_index_80789[8];
  assign array_update_80796[9] = add_80666 == 32'h0000_0009 ? add_80795 : array_index_80789[9];
  assign array_update_80797[0] = add_80123 == 32'h0000_0000 ? array_update_80796 : array_update_80786[0];
  assign array_update_80797[1] = add_80123 == 32'h0000_0001 ? array_update_80796 : array_update_80786[1];
  assign array_update_80797[2] = add_80123 == 32'h0000_0002 ? array_update_80796 : array_update_80786[2];
  assign array_update_80797[3] = add_80123 == 32'h0000_0003 ? array_update_80796 : array_update_80786[3];
  assign array_update_80797[4] = add_80123 == 32'h0000_0004 ? array_update_80796 : array_update_80786[4];
  assign array_update_80797[5] = add_80123 == 32'h0000_0005 ? array_update_80796 : array_update_80786[5];
  assign array_update_80797[6] = add_80123 == 32'h0000_0006 ? array_update_80796 : array_update_80786[6];
  assign array_update_80797[7] = add_80123 == 32'h0000_0007 ? array_update_80796 : array_update_80786[7];
  assign array_update_80797[8] = add_80123 == 32'h0000_0008 ? array_update_80796 : array_update_80786[8];
  assign array_update_80797[9] = add_80123 == 32'h0000_0009 ? array_update_80796 : array_update_80786[9];
  assign array_index_80799 = array_update_80797[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign add_80801 = add_80666 + 32'h0000_0001;
  assign array_update_80802[0] = add_80801 == 32'h0000_0000 ? 32'h0000_0000 : array_index_80799[0];
  assign array_update_80802[1] = add_80801 == 32'h0000_0001 ? 32'h0000_0000 : array_index_80799[1];
  assign array_update_80802[2] = add_80801 == 32'h0000_0002 ? 32'h0000_0000 : array_index_80799[2];
  assign array_update_80802[3] = add_80801 == 32'h0000_0003 ? 32'h0000_0000 : array_index_80799[3];
  assign array_update_80802[4] = add_80801 == 32'h0000_0004 ? 32'h0000_0000 : array_index_80799[4];
  assign array_update_80802[5] = add_80801 == 32'h0000_0005 ? 32'h0000_0000 : array_index_80799[5];
  assign array_update_80802[6] = add_80801 == 32'h0000_0006 ? 32'h0000_0000 : array_index_80799[6];
  assign array_update_80802[7] = add_80801 == 32'h0000_0007 ? 32'h0000_0000 : array_index_80799[7];
  assign array_update_80802[8] = add_80801 == 32'h0000_0008 ? 32'h0000_0000 : array_index_80799[8];
  assign array_update_80802[9] = add_80801 == 32'h0000_0009 ? 32'h0000_0000 : array_index_80799[9];
  assign literal_80803 = 32'h0000_0000;
  assign array_update_80804[0] = add_80123 == 32'h0000_0000 ? array_update_80802 : array_update_80797[0];
  assign array_update_80804[1] = add_80123 == 32'h0000_0001 ? array_update_80802 : array_update_80797[1];
  assign array_update_80804[2] = add_80123 == 32'h0000_0002 ? array_update_80802 : array_update_80797[2];
  assign array_update_80804[3] = add_80123 == 32'h0000_0003 ? array_update_80802 : array_update_80797[3];
  assign array_update_80804[4] = add_80123 == 32'h0000_0004 ? array_update_80802 : array_update_80797[4];
  assign array_update_80804[5] = add_80123 == 32'h0000_0005 ? array_update_80802 : array_update_80797[5];
  assign array_update_80804[6] = add_80123 == 32'h0000_0006 ? array_update_80802 : array_update_80797[6];
  assign array_update_80804[7] = add_80123 == 32'h0000_0007 ? array_update_80802 : array_update_80797[7];
  assign array_update_80804[8] = add_80123 == 32'h0000_0008 ? array_update_80802 : array_update_80797[8];
  assign array_update_80804[9] = add_80123 == 32'h0000_0009 ? array_update_80802 : array_update_80797[9];
  assign array_index_80806 = array_update_72021[literal_80803 > 32'h0000_0009 ? 4'h9 : literal_80803[3:0]];
  assign array_index_80807 = array_update_80804[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_80811 = smul32b_32b_x_32b(array_index_80130[literal_80803 > 32'h0000_0009 ? 4'h9 : literal_80803[3:0]], array_index_80806[add_80801 > 32'h0000_0009 ? 4'h9 : add_80801[3:0]]);
  assign add_80813 = array_index_80807[add_80801 > 32'h0000_0009 ? 4'h9 : add_80801[3:0]] + smul_80811;
  assign array_update_80815[0] = add_80801 == 32'h0000_0000 ? add_80813 : array_index_80807[0];
  assign array_update_80815[1] = add_80801 == 32'h0000_0001 ? add_80813 : array_index_80807[1];
  assign array_update_80815[2] = add_80801 == 32'h0000_0002 ? add_80813 : array_index_80807[2];
  assign array_update_80815[3] = add_80801 == 32'h0000_0003 ? add_80813 : array_index_80807[3];
  assign array_update_80815[4] = add_80801 == 32'h0000_0004 ? add_80813 : array_index_80807[4];
  assign array_update_80815[5] = add_80801 == 32'h0000_0005 ? add_80813 : array_index_80807[5];
  assign array_update_80815[6] = add_80801 == 32'h0000_0006 ? add_80813 : array_index_80807[6];
  assign array_update_80815[7] = add_80801 == 32'h0000_0007 ? add_80813 : array_index_80807[7];
  assign array_update_80815[8] = add_80801 == 32'h0000_0008 ? add_80813 : array_index_80807[8];
  assign array_update_80815[9] = add_80801 == 32'h0000_0009 ? add_80813 : array_index_80807[9];
  assign add_80816 = literal_80803 + 32'h0000_0001;
  assign array_update_80817[0] = add_80123 == 32'h0000_0000 ? array_update_80815 : array_update_80804[0];
  assign array_update_80817[1] = add_80123 == 32'h0000_0001 ? array_update_80815 : array_update_80804[1];
  assign array_update_80817[2] = add_80123 == 32'h0000_0002 ? array_update_80815 : array_update_80804[2];
  assign array_update_80817[3] = add_80123 == 32'h0000_0003 ? array_update_80815 : array_update_80804[3];
  assign array_update_80817[4] = add_80123 == 32'h0000_0004 ? array_update_80815 : array_update_80804[4];
  assign array_update_80817[5] = add_80123 == 32'h0000_0005 ? array_update_80815 : array_update_80804[5];
  assign array_update_80817[6] = add_80123 == 32'h0000_0006 ? array_update_80815 : array_update_80804[6];
  assign array_update_80817[7] = add_80123 == 32'h0000_0007 ? array_update_80815 : array_update_80804[7];
  assign array_update_80817[8] = add_80123 == 32'h0000_0008 ? array_update_80815 : array_update_80804[8];
  assign array_update_80817[9] = add_80123 == 32'h0000_0009 ? array_update_80815 : array_update_80804[9];
  assign array_index_80819 = array_update_72021[add_80816 > 32'h0000_0009 ? 4'h9 : add_80816[3:0]];
  assign array_index_80820 = array_update_80817[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_80824 = smul32b_32b_x_32b(array_index_80130[add_80816 > 32'h0000_0009 ? 4'h9 : add_80816[3:0]], array_index_80819[add_80801 > 32'h0000_0009 ? 4'h9 : add_80801[3:0]]);
  assign add_80826 = array_index_80820[add_80801 > 32'h0000_0009 ? 4'h9 : add_80801[3:0]] + smul_80824;
  assign array_update_80828[0] = add_80801 == 32'h0000_0000 ? add_80826 : array_index_80820[0];
  assign array_update_80828[1] = add_80801 == 32'h0000_0001 ? add_80826 : array_index_80820[1];
  assign array_update_80828[2] = add_80801 == 32'h0000_0002 ? add_80826 : array_index_80820[2];
  assign array_update_80828[3] = add_80801 == 32'h0000_0003 ? add_80826 : array_index_80820[3];
  assign array_update_80828[4] = add_80801 == 32'h0000_0004 ? add_80826 : array_index_80820[4];
  assign array_update_80828[5] = add_80801 == 32'h0000_0005 ? add_80826 : array_index_80820[5];
  assign array_update_80828[6] = add_80801 == 32'h0000_0006 ? add_80826 : array_index_80820[6];
  assign array_update_80828[7] = add_80801 == 32'h0000_0007 ? add_80826 : array_index_80820[7];
  assign array_update_80828[8] = add_80801 == 32'h0000_0008 ? add_80826 : array_index_80820[8];
  assign array_update_80828[9] = add_80801 == 32'h0000_0009 ? add_80826 : array_index_80820[9];
  assign add_80829 = add_80816 + 32'h0000_0001;
  assign array_update_80830[0] = add_80123 == 32'h0000_0000 ? array_update_80828 : array_update_80817[0];
  assign array_update_80830[1] = add_80123 == 32'h0000_0001 ? array_update_80828 : array_update_80817[1];
  assign array_update_80830[2] = add_80123 == 32'h0000_0002 ? array_update_80828 : array_update_80817[2];
  assign array_update_80830[3] = add_80123 == 32'h0000_0003 ? array_update_80828 : array_update_80817[3];
  assign array_update_80830[4] = add_80123 == 32'h0000_0004 ? array_update_80828 : array_update_80817[4];
  assign array_update_80830[5] = add_80123 == 32'h0000_0005 ? array_update_80828 : array_update_80817[5];
  assign array_update_80830[6] = add_80123 == 32'h0000_0006 ? array_update_80828 : array_update_80817[6];
  assign array_update_80830[7] = add_80123 == 32'h0000_0007 ? array_update_80828 : array_update_80817[7];
  assign array_update_80830[8] = add_80123 == 32'h0000_0008 ? array_update_80828 : array_update_80817[8];
  assign array_update_80830[9] = add_80123 == 32'h0000_0009 ? array_update_80828 : array_update_80817[9];
  assign array_index_80832 = array_update_72021[add_80829 > 32'h0000_0009 ? 4'h9 : add_80829[3:0]];
  assign array_index_80833 = array_update_80830[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_80837 = smul32b_32b_x_32b(array_index_80130[add_80829 > 32'h0000_0009 ? 4'h9 : add_80829[3:0]], array_index_80832[add_80801 > 32'h0000_0009 ? 4'h9 : add_80801[3:0]]);
  assign add_80839 = array_index_80833[add_80801 > 32'h0000_0009 ? 4'h9 : add_80801[3:0]] + smul_80837;
  assign array_update_80841[0] = add_80801 == 32'h0000_0000 ? add_80839 : array_index_80833[0];
  assign array_update_80841[1] = add_80801 == 32'h0000_0001 ? add_80839 : array_index_80833[1];
  assign array_update_80841[2] = add_80801 == 32'h0000_0002 ? add_80839 : array_index_80833[2];
  assign array_update_80841[3] = add_80801 == 32'h0000_0003 ? add_80839 : array_index_80833[3];
  assign array_update_80841[4] = add_80801 == 32'h0000_0004 ? add_80839 : array_index_80833[4];
  assign array_update_80841[5] = add_80801 == 32'h0000_0005 ? add_80839 : array_index_80833[5];
  assign array_update_80841[6] = add_80801 == 32'h0000_0006 ? add_80839 : array_index_80833[6];
  assign array_update_80841[7] = add_80801 == 32'h0000_0007 ? add_80839 : array_index_80833[7];
  assign array_update_80841[8] = add_80801 == 32'h0000_0008 ? add_80839 : array_index_80833[8];
  assign array_update_80841[9] = add_80801 == 32'h0000_0009 ? add_80839 : array_index_80833[9];
  assign add_80842 = add_80829 + 32'h0000_0001;
  assign array_update_80843[0] = add_80123 == 32'h0000_0000 ? array_update_80841 : array_update_80830[0];
  assign array_update_80843[1] = add_80123 == 32'h0000_0001 ? array_update_80841 : array_update_80830[1];
  assign array_update_80843[2] = add_80123 == 32'h0000_0002 ? array_update_80841 : array_update_80830[2];
  assign array_update_80843[3] = add_80123 == 32'h0000_0003 ? array_update_80841 : array_update_80830[3];
  assign array_update_80843[4] = add_80123 == 32'h0000_0004 ? array_update_80841 : array_update_80830[4];
  assign array_update_80843[5] = add_80123 == 32'h0000_0005 ? array_update_80841 : array_update_80830[5];
  assign array_update_80843[6] = add_80123 == 32'h0000_0006 ? array_update_80841 : array_update_80830[6];
  assign array_update_80843[7] = add_80123 == 32'h0000_0007 ? array_update_80841 : array_update_80830[7];
  assign array_update_80843[8] = add_80123 == 32'h0000_0008 ? array_update_80841 : array_update_80830[8];
  assign array_update_80843[9] = add_80123 == 32'h0000_0009 ? array_update_80841 : array_update_80830[9];
  assign array_index_80845 = array_update_72021[add_80842 > 32'h0000_0009 ? 4'h9 : add_80842[3:0]];
  assign array_index_80846 = array_update_80843[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_80850 = smul32b_32b_x_32b(array_index_80130[add_80842 > 32'h0000_0009 ? 4'h9 : add_80842[3:0]], array_index_80845[add_80801 > 32'h0000_0009 ? 4'h9 : add_80801[3:0]]);
  assign add_80852 = array_index_80846[add_80801 > 32'h0000_0009 ? 4'h9 : add_80801[3:0]] + smul_80850;
  assign array_update_80854[0] = add_80801 == 32'h0000_0000 ? add_80852 : array_index_80846[0];
  assign array_update_80854[1] = add_80801 == 32'h0000_0001 ? add_80852 : array_index_80846[1];
  assign array_update_80854[2] = add_80801 == 32'h0000_0002 ? add_80852 : array_index_80846[2];
  assign array_update_80854[3] = add_80801 == 32'h0000_0003 ? add_80852 : array_index_80846[3];
  assign array_update_80854[4] = add_80801 == 32'h0000_0004 ? add_80852 : array_index_80846[4];
  assign array_update_80854[5] = add_80801 == 32'h0000_0005 ? add_80852 : array_index_80846[5];
  assign array_update_80854[6] = add_80801 == 32'h0000_0006 ? add_80852 : array_index_80846[6];
  assign array_update_80854[7] = add_80801 == 32'h0000_0007 ? add_80852 : array_index_80846[7];
  assign array_update_80854[8] = add_80801 == 32'h0000_0008 ? add_80852 : array_index_80846[8];
  assign array_update_80854[9] = add_80801 == 32'h0000_0009 ? add_80852 : array_index_80846[9];
  assign add_80855 = add_80842 + 32'h0000_0001;
  assign array_update_80856[0] = add_80123 == 32'h0000_0000 ? array_update_80854 : array_update_80843[0];
  assign array_update_80856[1] = add_80123 == 32'h0000_0001 ? array_update_80854 : array_update_80843[1];
  assign array_update_80856[2] = add_80123 == 32'h0000_0002 ? array_update_80854 : array_update_80843[2];
  assign array_update_80856[3] = add_80123 == 32'h0000_0003 ? array_update_80854 : array_update_80843[3];
  assign array_update_80856[4] = add_80123 == 32'h0000_0004 ? array_update_80854 : array_update_80843[4];
  assign array_update_80856[5] = add_80123 == 32'h0000_0005 ? array_update_80854 : array_update_80843[5];
  assign array_update_80856[6] = add_80123 == 32'h0000_0006 ? array_update_80854 : array_update_80843[6];
  assign array_update_80856[7] = add_80123 == 32'h0000_0007 ? array_update_80854 : array_update_80843[7];
  assign array_update_80856[8] = add_80123 == 32'h0000_0008 ? array_update_80854 : array_update_80843[8];
  assign array_update_80856[9] = add_80123 == 32'h0000_0009 ? array_update_80854 : array_update_80843[9];
  assign array_index_80858 = array_update_72021[add_80855 > 32'h0000_0009 ? 4'h9 : add_80855[3:0]];
  assign array_index_80859 = array_update_80856[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_80863 = smul32b_32b_x_32b(array_index_80130[add_80855 > 32'h0000_0009 ? 4'h9 : add_80855[3:0]], array_index_80858[add_80801 > 32'h0000_0009 ? 4'h9 : add_80801[3:0]]);
  assign add_80865 = array_index_80859[add_80801 > 32'h0000_0009 ? 4'h9 : add_80801[3:0]] + smul_80863;
  assign array_update_80867[0] = add_80801 == 32'h0000_0000 ? add_80865 : array_index_80859[0];
  assign array_update_80867[1] = add_80801 == 32'h0000_0001 ? add_80865 : array_index_80859[1];
  assign array_update_80867[2] = add_80801 == 32'h0000_0002 ? add_80865 : array_index_80859[2];
  assign array_update_80867[3] = add_80801 == 32'h0000_0003 ? add_80865 : array_index_80859[3];
  assign array_update_80867[4] = add_80801 == 32'h0000_0004 ? add_80865 : array_index_80859[4];
  assign array_update_80867[5] = add_80801 == 32'h0000_0005 ? add_80865 : array_index_80859[5];
  assign array_update_80867[6] = add_80801 == 32'h0000_0006 ? add_80865 : array_index_80859[6];
  assign array_update_80867[7] = add_80801 == 32'h0000_0007 ? add_80865 : array_index_80859[7];
  assign array_update_80867[8] = add_80801 == 32'h0000_0008 ? add_80865 : array_index_80859[8];
  assign array_update_80867[9] = add_80801 == 32'h0000_0009 ? add_80865 : array_index_80859[9];
  assign add_80868 = add_80855 + 32'h0000_0001;
  assign array_update_80869[0] = add_80123 == 32'h0000_0000 ? array_update_80867 : array_update_80856[0];
  assign array_update_80869[1] = add_80123 == 32'h0000_0001 ? array_update_80867 : array_update_80856[1];
  assign array_update_80869[2] = add_80123 == 32'h0000_0002 ? array_update_80867 : array_update_80856[2];
  assign array_update_80869[3] = add_80123 == 32'h0000_0003 ? array_update_80867 : array_update_80856[3];
  assign array_update_80869[4] = add_80123 == 32'h0000_0004 ? array_update_80867 : array_update_80856[4];
  assign array_update_80869[5] = add_80123 == 32'h0000_0005 ? array_update_80867 : array_update_80856[5];
  assign array_update_80869[6] = add_80123 == 32'h0000_0006 ? array_update_80867 : array_update_80856[6];
  assign array_update_80869[7] = add_80123 == 32'h0000_0007 ? array_update_80867 : array_update_80856[7];
  assign array_update_80869[8] = add_80123 == 32'h0000_0008 ? array_update_80867 : array_update_80856[8];
  assign array_update_80869[9] = add_80123 == 32'h0000_0009 ? array_update_80867 : array_update_80856[9];
  assign array_index_80871 = array_update_72021[add_80868 > 32'h0000_0009 ? 4'h9 : add_80868[3:0]];
  assign array_index_80872 = array_update_80869[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_80876 = smul32b_32b_x_32b(array_index_80130[add_80868 > 32'h0000_0009 ? 4'h9 : add_80868[3:0]], array_index_80871[add_80801 > 32'h0000_0009 ? 4'h9 : add_80801[3:0]]);
  assign add_80878 = array_index_80872[add_80801 > 32'h0000_0009 ? 4'h9 : add_80801[3:0]] + smul_80876;
  assign array_update_80880[0] = add_80801 == 32'h0000_0000 ? add_80878 : array_index_80872[0];
  assign array_update_80880[1] = add_80801 == 32'h0000_0001 ? add_80878 : array_index_80872[1];
  assign array_update_80880[2] = add_80801 == 32'h0000_0002 ? add_80878 : array_index_80872[2];
  assign array_update_80880[3] = add_80801 == 32'h0000_0003 ? add_80878 : array_index_80872[3];
  assign array_update_80880[4] = add_80801 == 32'h0000_0004 ? add_80878 : array_index_80872[4];
  assign array_update_80880[5] = add_80801 == 32'h0000_0005 ? add_80878 : array_index_80872[5];
  assign array_update_80880[6] = add_80801 == 32'h0000_0006 ? add_80878 : array_index_80872[6];
  assign array_update_80880[7] = add_80801 == 32'h0000_0007 ? add_80878 : array_index_80872[7];
  assign array_update_80880[8] = add_80801 == 32'h0000_0008 ? add_80878 : array_index_80872[8];
  assign array_update_80880[9] = add_80801 == 32'h0000_0009 ? add_80878 : array_index_80872[9];
  assign add_80881 = add_80868 + 32'h0000_0001;
  assign array_update_80882[0] = add_80123 == 32'h0000_0000 ? array_update_80880 : array_update_80869[0];
  assign array_update_80882[1] = add_80123 == 32'h0000_0001 ? array_update_80880 : array_update_80869[1];
  assign array_update_80882[2] = add_80123 == 32'h0000_0002 ? array_update_80880 : array_update_80869[2];
  assign array_update_80882[3] = add_80123 == 32'h0000_0003 ? array_update_80880 : array_update_80869[3];
  assign array_update_80882[4] = add_80123 == 32'h0000_0004 ? array_update_80880 : array_update_80869[4];
  assign array_update_80882[5] = add_80123 == 32'h0000_0005 ? array_update_80880 : array_update_80869[5];
  assign array_update_80882[6] = add_80123 == 32'h0000_0006 ? array_update_80880 : array_update_80869[6];
  assign array_update_80882[7] = add_80123 == 32'h0000_0007 ? array_update_80880 : array_update_80869[7];
  assign array_update_80882[8] = add_80123 == 32'h0000_0008 ? array_update_80880 : array_update_80869[8];
  assign array_update_80882[9] = add_80123 == 32'h0000_0009 ? array_update_80880 : array_update_80869[9];
  assign array_index_80884 = array_update_72021[add_80881 > 32'h0000_0009 ? 4'h9 : add_80881[3:0]];
  assign array_index_80885 = array_update_80882[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_80889 = smul32b_32b_x_32b(array_index_80130[add_80881 > 32'h0000_0009 ? 4'h9 : add_80881[3:0]], array_index_80884[add_80801 > 32'h0000_0009 ? 4'h9 : add_80801[3:0]]);
  assign add_80891 = array_index_80885[add_80801 > 32'h0000_0009 ? 4'h9 : add_80801[3:0]] + smul_80889;
  assign array_update_80893[0] = add_80801 == 32'h0000_0000 ? add_80891 : array_index_80885[0];
  assign array_update_80893[1] = add_80801 == 32'h0000_0001 ? add_80891 : array_index_80885[1];
  assign array_update_80893[2] = add_80801 == 32'h0000_0002 ? add_80891 : array_index_80885[2];
  assign array_update_80893[3] = add_80801 == 32'h0000_0003 ? add_80891 : array_index_80885[3];
  assign array_update_80893[4] = add_80801 == 32'h0000_0004 ? add_80891 : array_index_80885[4];
  assign array_update_80893[5] = add_80801 == 32'h0000_0005 ? add_80891 : array_index_80885[5];
  assign array_update_80893[6] = add_80801 == 32'h0000_0006 ? add_80891 : array_index_80885[6];
  assign array_update_80893[7] = add_80801 == 32'h0000_0007 ? add_80891 : array_index_80885[7];
  assign array_update_80893[8] = add_80801 == 32'h0000_0008 ? add_80891 : array_index_80885[8];
  assign array_update_80893[9] = add_80801 == 32'h0000_0009 ? add_80891 : array_index_80885[9];
  assign add_80894 = add_80881 + 32'h0000_0001;
  assign array_update_80895[0] = add_80123 == 32'h0000_0000 ? array_update_80893 : array_update_80882[0];
  assign array_update_80895[1] = add_80123 == 32'h0000_0001 ? array_update_80893 : array_update_80882[1];
  assign array_update_80895[2] = add_80123 == 32'h0000_0002 ? array_update_80893 : array_update_80882[2];
  assign array_update_80895[3] = add_80123 == 32'h0000_0003 ? array_update_80893 : array_update_80882[3];
  assign array_update_80895[4] = add_80123 == 32'h0000_0004 ? array_update_80893 : array_update_80882[4];
  assign array_update_80895[5] = add_80123 == 32'h0000_0005 ? array_update_80893 : array_update_80882[5];
  assign array_update_80895[6] = add_80123 == 32'h0000_0006 ? array_update_80893 : array_update_80882[6];
  assign array_update_80895[7] = add_80123 == 32'h0000_0007 ? array_update_80893 : array_update_80882[7];
  assign array_update_80895[8] = add_80123 == 32'h0000_0008 ? array_update_80893 : array_update_80882[8];
  assign array_update_80895[9] = add_80123 == 32'h0000_0009 ? array_update_80893 : array_update_80882[9];
  assign array_index_80897 = array_update_72021[add_80894 > 32'h0000_0009 ? 4'h9 : add_80894[3:0]];
  assign array_index_80898 = array_update_80895[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_80902 = smul32b_32b_x_32b(array_index_80130[add_80894 > 32'h0000_0009 ? 4'h9 : add_80894[3:0]], array_index_80897[add_80801 > 32'h0000_0009 ? 4'h9 : add_80801[3:0]]);
  assign add_80904 = array_index_80898[add_80801 > 32'h0000_0009 ? 4'h9 : add_80801[3:0]] + smul_80902;
  assign array_update_80906[0] = add_80801 == 32'h0000_0000 ? add_80904 : array_index_80898[0];
  assign array_update_80906[1] = add_80801 == 32'h0000_0001 ? add_80904 : array_index_80898[1];
  assign array_update_80906[2] = add_80801 == 32'h0000_0002 ? add_80904 : array_index_80898[2];
  assign array_update_80906[3] = add_80801 == 32'h0000_0003 ? add_80904 : array_index_80898[3];
  assign array_update_80906[4] = add_80801 == 32'h0000_0004 ? add_80904 : array_index_80898[4];
  assign array_update_80906[5] = add_80801 == 32'h0000_0005 ? add_80904 : array_index_80898[5];
  assign array_update_80906[6] = add_80801 == 32'h0000_0006 ? add_80904 : array_index_80898[6];
  assign array_update_80906[7] = add_80801 == 32'h0000_0007 ? add_80904 : array_index_80898[7];
  assign array_update_80906[8] = add_80801 == 32'h0000_0008 ? add_80904 : array_index_80898[8];
  assign array_update_80906[9] = add_80801 == 32'h0000_0009 ? add_80904 : array_index_80898[9];
  assign add_80907 = add_80894 + 32'h0000_0001;
  assign array_update_80908[0] = add_80123 == 32'h0000_0000 ? array_update_80906 : array_update_80895[0];
  assign array_update_80908[1] = add_80123 == 32'h0000_0001 ? array_update_80906 : array_update_80895[1];
  assign array_update_80908[2] = add_80123 == 32'h0000_0002 ? array_update_80906 : array_update_80895[2];
  assign array_update_80908[3] = add_80123 == 32'h0000_0003 ? array_update_80906 : array_update_80895[3];
  assign array_update_80908[4] = add_80123 == 32'h0000_0004 ? array_update_80906 : array_update_80895[4];
  assign array_update_80908[5] = add_80123 == 32'h0000_0005 ? array_update_80906 : array_update_80895[5];
  assign array_update_80908[6] = add_80123 == 32'h0000_0006 ? array_update_80906 : array_update_80895[6];
  assign array_update_80908[7] = add_80123 == 32'h0000_0007 ? array_update_80906 : array_update_80895[7];
  assign array_update_80908[8] = add_80123 == 32'h0000_0008 ? array_update_80906 : array_update_80895[8];
  assign array_update_80908[9] = add_80123 == 32'h0000_0009 ? array_update_80906 : array_update_80895[9];
  assign array_index_80910 = array_update_72021[add_80907 > 32'h0000_0009 ? 4'h9 : add_80907[3:0]];
  assign array_index_80911 = array_update_80908[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_80915 = smul32b_32b_x_32b(array_index_80130[add_80907 > 32'h0000_0009 ? 4'h9 : add_80907[3:0]], array_index_80910[add_80801 > 32'h0000_0009 ? 4'h9 : add_80801[3:0]]);
  assign add_80917 = array_index_80911[add_80801 > 32'h0000_0009 ? 4'h9 : add_80801[3:0]] + smul_80915;
  assign array_update_80919[0] = add_80801 == 32'h0000_0000 ? add_80917 : array_index_80911[0];
  assign array_update_80919[1] = add_80801 == 32'h0000_0001 ? add_80917 : array_index_80911[1];
  assign array_update_80919[2] = add_80801 == 32'h0000_0002 ? add_80917 : array_index_80911[2];
  assign array_update_80919[3] = add_80801 == 32'h0000_0003 ? add_80917 : array_index_80911[3];
  assign array_update_80919[4] = add_80801 == 32'h0000_0004 ? add_80917 : array_index_80911[4];
  assign array_update_80919[5] = add_80801 == 32'h0000_0005 ? add_80917 : array_index_80911[5];
  assign array_update_80919[6] = add_80801 == 32'h0000_0006 ? add_80917 : array_index_80911[6];
  assign array_update_80919[7] = add_80801 == 32'h0000_0007 ? add_80917 : array_index_80911[7];
  assign array_update_80919[8] = add_80801 == 32'h0000_0008 ? add_80917 : array_index_80911[8];
  assign array_update_80919[9] = add_80801 == 32'h0000_0009 ? add_80917 : array_index_80911[9];
  assign add_80920 = add_80907 + 32'h0000_0001;
  assign array_update_80921[0] = add_80123 == 32'h0000_0000 ? array_update_80919 : array_update_80908[0];
  assign array_update_80921[1] = add_80123 == 32'h0000_0001 ? array_update_80919 : array_update_80908[1];
  assign array_update_80921[2] = add_80123 == 32'h0000_0002 ? array_update_80919 : array_update_80908[2];
  assign array_update_80921[3] = add_80123 == 32'h0000_0003 ? array_update_80919 : array_update_80908[3];
  assign array_update_80921[4] = add_80123 == 32'h0000_0004 ? array_update_80919 : array_update_80908[4];
  assign array_update_80921[5] = add_80123 == 32'h0000_0005 ? array_update_80919 : array_update_80908[5];
  assign array_update_80921[6] = add_80123 == 32'h0000_0006 ? array_update_80919 : array_update_80908[6];
  assign array_update_80921[7] = add_80123 == 32'h0000_0007 ? array_update_80919 : array_update_80908[7];
  assign array_update_80921[8] = add_80123 == 32'h0000_0008 ? array_update_80919 : array_update_80908[8];
  assign array_update_80921[9] = add_80123 == 32'h0000_0009 ? array_update_80919 : array_update_80908[9];
  assign array_index_80923 = array_update_72021[add_80920 > 32'h0000_0009 ? 4'h9 : add_80920[3:0]];
  assign array_index_80924 = array_update_80921[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_80928 = smul32b_32b_x_32b(array_index_80130[add_80920 > 32'h0000_0009 ? 4'h9 : add_80920[3:0]], array_index_80923[add_80801 > 32'h0000_0009 ? 4'h9 : add_80801[3:0]]);
  assign add_80930 = array_index_80924[add_80801 > 32'h0000_0009 ? 4'h9 : add_80801[3:0]] + smul_80928;
  assign array_update_80931[0] = add_80801 == 32'h0000_0000 ? add_80930 : array_index_80924[0];
  assign array_update_80931[1] = add_80801 == 32'h0000_0001 ? add_80930 : array_index_80924[1];
  assign array_update_80931[2] = add_80801 == 32'h0000_0002 ? add_80930 : array_index_80924[2];
  assign array_update_80931[3] = add_80801 == 32'h0000_0003 ? add_80930 : array_index_80924[3];
  assign array_update_80931[4] = add_80801 == 32'h0000_0004 ? add_80930 : array_index_80924[4];
  assign array_update_80931[5] = add_80801 == 32'h0000_0005 ? add_80930 : array_index_80924[5];
  assign array_update_80931[6] = add_80801 == 32'h0000_0006 ? add_80930 : array_index_80924[6];
  assign array_update_80931[7] = add_80801 == 32'h0000_0007 ? add_80930 : array_index_80924[7];
  assign array_update_80931[8] = add_80801 == 32'h0000_0008 ? add_80930 : array_index_80924[8];
  assign array_update_80931[9] = add_80801 == 32'h0000_0009 ? add_80930 : array_index_80924[9];
  assign array_update_80932[0] = add_80123 == 32'h0000_0000 ? array_update_80931 : array_update_80921[0];
  assign array_update_80932[1] = add_80123 == 32'h0000_0001 ? array_update_80931 : array_update_80921[1];
  assign array_update_80932[2] = add_80123 == 32'h0000_0002 ? array_update_80931 : array_update_80921[2];
  assign array_update_80932[3] = add_80123 == 32'h0000_0003 ? array_update_80931 : array_update_80921[3];
  assign array_update_80932[4] = add_80123 == 32'h0000_0004 ? array_update_80931 : array_update_80921[4];
  assign array_update_80932[5] = add_80123 == 32'h0000_0005 ? array_update_80931 : array_update_80921[5];
  assign array_update_80932[6] = add_80123 == 32'h0000_0006 ? array_update_80931 : array_update_80921[6];
  assign array_update_80932[7] = add_80123 == 32'h0000_0007 ? array_update_80931 : array_update_80921[7];
  assign array_update_80932[8] = add_80123 == 32'h0000_0008 ? array_update_80931 : array_update_80921[8];
  assign array_update_80932[9] = add_80123 == 32'h0000_0009 ? array_update_80931 : array_update_80921[9];
  assign array_index_80934 = array_update_80932[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign add_80936 = add_80801 + 32'h0000_0001;
  assign array_update_80937[0] = add_80936 == 32'h0000_0000 ? 32'h0000_0000 : array_index_80934[0];
  assign array_update_80937[1] = add_80936 == 32'h0000_0001 ? 32'h0000_0000 : array_index_80934[1];
  assign array_update_80937[2] = add_80936 == 32'h0000_0002 ? 32'h0000_0000 : array_index_80934[2];
  assign array_update_80937[3] = add_80936 == 32'h0000_0003 ? 32'h0000_0000 : array_index_80934[3];
  assign array_update_80937[4] = add_80936 == 32'h0000_0004 ? 32'h0000_0000 : array_index_80934[4];
  assign array_update_80937[5] = add_80936 == 32'h0000_0005 ? 32'h0000_0000 : array_index_80934[5];
  assign array_update_80937[6] = add_80936 == 32'h0000_0006 ? 32'h0000_0000 : array_index_80934[6];
  assign array_update_80937[7] = add_80936 == 32'h0000_0007 ? 32'h0000_0000 : array_index_80934[7];
  assign array_update_80937[8] = add_80936 == 32'h0000_0008 ? 32'h0000_0000 : array_index_80934[8];
  assign array_update_80937[9] = add_80936 == 32'h0000_0009 ? 32'h0000_0000 : array_index_80934[9];
  assign literal_80938 = 32'h0000_0000;
  assign array_update_80939[0] = add_80123 == 32'h0000_0000 ? array_update_80937 : array_update_80932[0];
  assign array_update_80939[1] = add_80123 == 32'h0000_0001 ? array_update_80937 : array_update_80932[1];
  assign array_update_80939[2] = add_80123 == 32'h0000_0002 ? array_update_80937 : array_update_80932[2];
  assign array_update_80939[3] = add_80123 == 32'h0000_0003 ? array_update_80937 : array_update_80932[3];
  assign array_update_80939[4] = add_80123 == 32'h0000_0004 ? array_update_80937 : array_update_80932[4];
  assign array_update_80939[5] = add_80123 == 32'h0000_0005 ? array_update_80937 : array_update_80932[5];
  assign array_update_80939[6] = add_80123 == 32'h0000_0006 ? array_update_80937 : array_update_80932[6];
  assign array_update_80939[7] = add_80123 == 32'h0000_0007 ? array_update_80937 : array_update_80932[7];
  assign array_update_80939[8] = add_80123 == 32'h0000_0008 ? array_update_80937 : array_update_80932[8];
  assign array_update_80939[9] = add_80123 == 32'h0000_0009 ? array_update_80937 : array_update_80932[9];
  assign array_index_80941 = array_update_72021[literal_80938 > 32'h0000_0009 ? 4'h9 : literal_80938[3:0]];
  assign array_index_80942 = array_update_80939[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_80946 = smul32b_32b_x_32b(array_index_80130[literal_80938 > 32'h0000_0009 ? 4'h9 : literal_80938[3:0]], array_index_80941[add_80936 > 32'h0000_0009 ? 4'h9 : add_80936[3:0]]);
  assign add_80948 = array_index_80942[add_80936 > 32'h0000_0009 ? 4'h9 : add_80936[3:0]] + smul_80946;
  assign array_update_80950[0] = add_80936 == 32'h0000_0000 ? add_80948 : array_index_80942[0];
  assign array_update_80950[1] = add_80936 == 32'h0000_0001 ? add_80948 : array_index_80942[1];
  assign array_update_80950[2] = add_80936 == 32'h0000_0002 ? add_80948 : array_index_80942[2];
  assign array_update_80950[3] = add_80936 == 32'h0000_0003 ? add_80948 : array_index_80942[3];
  assign array_update_80950[4] = add_80936 == 32'h0000_0004 ? add_80948 : array_index_80942[4];
  assign array_update_80950[5] = add_80936 == 32'h0000_0005 ? add_80948 : array_index_80942[5];
  assign array_update_80950[6] = add_80936 == 32'h0000_0006 ? add_80948 : array_index_80942[6];
  assign array_update_80950[7] = add_80936 == 32'h0000_0007 ? add_80948 : array_index_80942[7];
  assign array_update_80950[8] = add_80936 == 32'h0000_0008 ? add_80948 : array_index_80942[8];
  assign array_update_80950[9] = add_80936 == 32'h0000_0009 ? add_80948 : array_index_80942[9];
  assign add_80951 = literal_80938 + 32'h0000_0001;
  assign array_update_80952[0] = add_80123 == 32'h0000_0000 ? array_update_80950 : array_update_80939[0];
  assign array_update_80952[1] = add_80123 == 32'h0000_0001 ? array_update_80950 : array_update_80939[1];
  assign array_update_80952[2] = add_80123 == 32'h0000_0002 ? array_update_80950 : array_update_80939[2];
  assign array_update_80952[3] = add_80123 == 32'h0000_0003 ? array_update_80950 : array_update_80939[3];
  assign array_update_80952[4] = add_80123 == 32'h0000_0004 ? array_update_80950 : array_update_80939[4];
  assign array_update_80952[5] = add_80123 == 32'h0000_0005 ? array_update_80950 : array_update_80939[5];
  assign array_update_80952[6] = add_80123 == 32'h0000_0006 ? array_update_80950 : array_update_80939[6];
  assign array_update_80952[7] = add_80123 == 32'h0000_0007 ? array_update_80950 : array_update_80939[7];
  assign array_update_80952[8] = add_80123 == 32'h0000_0008 ? array_update_80950 : array_update_80939[8];
  assign array_update_80952[9] = add_80123 == 32'h0000_0009 ? array_update_80950 : array_update_80939[9];
  assign array_index_80954 = array_update_72021[add_80951 > 32'h0000_0009 ? 4'h9 : add_80951[3:0]];
  assign array_index_80955 = array_update_80952[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_80959 = smul32b_32b_x_32b(array_index_80130[add_80951 > 32'h0000_0009 ? 4'h9 : add_80951[3:0]], array_index_80954[add_80936 > 32'h0000_0009 ? 4'h9 : add_80936[3:0]]);
  assign add_80961 = array_index_80955[add_80936 > 32'h0000_0009 ? 4'h9 : add_80936[3:0]] + smul_80959;
  assign array_update_80963[0] = add_80936 == 32'h0000_0000 ? add_80961 : array_index_80955[0];
  assign array_update_80963[1] = add_80936 == 32'h0000_0001 ? add_80961 : array_index_80955[1];
  assign array_update_80963[2] = add_80936 == 32'h0000_0002 ? add_80961 : array_index_80955[2];
  assign array_update_80963[3] = add_80936 == 32'h0000_0003 ? add_80961 : array_index_80955[3];
  assign array_update_80963[4] = add_80936 == 32'h0000_0004 ? add_80961 : array_index_80955[4];
  assign array_update_80963[5] = add_80936 == 32'h0000_0005 ? add_80961 : array_index_80955[5];
  assign array_update_80963[6] = add_80936 == 32'h0000_0006 ? add_80961 : array_index_80955[6];
  assign array_update_80963[7] = add_80936 == 32'h0000_0007 ? add_80961 : array_index_80955[7];
  assign array_update_80963[8] = add_80936 == 32'h0000_0008 ? add_80961 : array_index_80955[8];
  assign array_update_80963[9] = add_80936 == 32'h0000_0009 ? add_80961 : array_index_80955[9];
  assign add_80964 = add_80951 + 32'h0000_0001;
  assign array_update_80965[0] = add_80123 == 32'h0000_0000 ? array_update_80963 : array_update_80952[0];
  assign array_update_80965[1] = add_80123 == 32'h0000_0001 ? array_update_80963 : array_update_80952[1];
  assign array_update_80965[2] = add_80123 == 32'h0000_0002 ? array_update_80963 : array_update_80952[2];
  assign array_update_80965[3] = add_80123 == 32'h0000_0003 ? array_update_80963 : array_update_80952[3];
  assign array_update_80965[4] = add_80123 == 32'h0000_0004 ? array_update_80963 : array_update_80952[4];
  assign array_update_80965[5] = add_80123 == 32'h0000_0005 ? array_update_80963 : array_update_80952[5];
  assign array_update_80965[6] = add_80123 == 32'h0000_0006 ? array_update_80963 : array_update_80952[6];
  assign array_update_80965[7] = add_80123 == 32'h0000_0007 ? array_update_80963 : array_update_80952[7];
  assign array_update_80965[8] = add_80123 == 32'h0000_0008 ? array_update_80963 : array_update_80952[8];
  assign array_update_80965[9] = add_80123 == 32'h0000_0009 ? array_update_80963 : array_update_80952[9];
  assign array_index_80967 = array_update_72021[add_80964 > 32'h0000_0009 ? 4'h9 : add_80964[3:0]];
  assign array_index_80968 = array_update_80965[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_80972 = smul32b_32b_x_32b(array_index_80130[add_80964 > 32'h0000_0009 ? 4'h9 : add_80964[3:0]], array_index_80967[add_80936 > 32'h0000_0009 ? 4'h9 : add_80936[3:0]]);
  assign add_80974 = array_index_80968[add_80936 > 32'h0000_0009 ? 4'h9 : add_80936[3:0]] + smul_80972;
  assign array_update_80976[0] = add_80936 == 32'h0000_0000 ? add_80974 : array_index_80968[0];
  assign array_update_80976[1] = add_80936 == 32'h0000_0001 ? add_80974 : array_index_80968[1];
  assign array_update_80976[2] = add_80936 == 32'h0000_0002 ? add_80974 : array_index_80968[2];
  assign array_update_80976[3] = add_80936 == 32'h0000_0003 ? add_80974 : array_index_80968[3];
  assign array_update_80976[4] = add_80936 == 32'h0000_0004 ? add_80974 : array_index_80968[4];
  assign array_update_80976[5] = add_80936 == 32'h0000_0005 ? add_80974 : array_index_80968[5];
  assign array_update_80976[6] = add_80936 == 32'h0000_0006 ? add_80974 : array_index_80968[6];
  assign array_update_80976[7] = add_80936 == 32'h0000_0007 ? add_80974 : array_index_80968[7];
  assign array_update_80976[8] = add_80936 == 32'h0000_0008 ? add_80974 : array_index_80968[8];
  assign array_update_80976[9] = add_80936 == 32'h0000_0009 ? add_80974 : array_index_80968[9];
  assign add_80977 = add_80964 + 32'h0000_0001;
  assign array_update_80978[0] = add_80123 == 32'h0000_0000 ? array_update_80976 : array_update_80965[0];
  assign array_update_80978[1] = add_80123 == 32'h0000_0001 ? array_update_80976 : array_update_80965[1];
  assign array_update_80978[2] = add_80123 == 32'h0000_0002 ? array_update_80976 : array_update_80965[2];
  assign array_update_80978[3] = add_80123 == 32'h0000_0003 ? array_update_80976 : array_update_80965[3];
  assign array_update_80978[4] = add_80123 == 32'h0000_0004 ? array_update_80976 : array_update_80965[4];
  assign array_update_80978[5] = add_80123 == 32'h0000_0005 ? array_update_80976 : array_update_80965[5];
  assign array_update_80978[6] = add_80123 == 32'h0000_0006 ? array_update_80976 : array_update_80965[6];
  assign array_update_80978[7] = add_80123 == 32'h0000_0007 ? array_update_80976 : array_update_80965[7];
  assign array_update_80978[8] = add_80123 == 32'h0000_0008 ? array_update_80976 : array_update_80965[8];
  assign array_update_80978[9] = add_80123 == 32'h0000_0009 ? array_update_80976 : array_update_80965[9];
  assign array_index_80980 = array_update_72021[add_80977 > 32'h0000_0009 ? 4'h9 : add_80977[3:0]];
  assign array_index_80981 = array_update_80978[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_80985 = smul32b_32b_x_32b(array_index_80130[add_80977 > 32'h0000_0009 ? 4'h9 : add_80977[3:0]], array_index_80980[add_80936 > 32'h0000_0009 ? 4'h9 : add_80936[3:0]]);
  assign add_80987 = array_index_80981[add_80936 > 32'h0000_0009 ? 4'h9 : add_80936[3:0]] + smul_80985;
  assign array_update_80989[0] = add_80936 == 32'h0000_0000 ? add_80987 : array_index_80981[0];
  assign array_update_80989[1] = add_80936 == 32'h0000_0001 ? add_80987 : array_index_80981[1];
  assign array_update_80989[2] = add_80936 == 32'h0000_0002 ? add_80987 : array_index_80981[2];
  assign array_update_80989[3] = add_80936 == 32'h0000_0003 ? add_80987 : array_index_80981[3];
  assign array_update_80989[4] = add_80936 == 32'h0000_0004 ? add_80987 : array_index_80981[4];
  assign array_update_80989[5] = add_80936 == 32'h0000_0005 ? add_80987 : array_index_80981[5];
  assign array_update_80989[6] = add_80936 == 32'h0000_0006 ? add_80987 : array_index_80981[6];
  assign array_update_80989[7] = add_80936 == 32'h0000_0007 ? add_80987 : array_index_80981[7];
  assign array_update_80989[8] = add_80936 == 32'h0000_0008 ? add_80987 : array_index_80981[8];
  assign array_update_80989[9] = add_80936 == 32'h0000_0009 ? add_80987 : array_index_80981[9];
  assign add_80990 = add_80977 + 32'h0000_0001;
  assign array_update_80991[0] = add_80123 == 32'h0000_0000 ? array_update_80989 : array_update_80978[0];
  assign array_update_80991[1] = add_80123 == 32'h0000_0001 ? array_update_80989 : array_update_80978[1];
  assign array_update_80991[2] = add_80123 == 32'h0000_0002 ? array_update_80989 : array_update_80978[2];
  assign array_update_80991[3] = add_80123 == 32'h0000_0003 ? array_update_80989 : array_update_80978[3];
  assign array_update_80991[4] = add_80123 == 32'h0000_0004 ? array_update_80989 : array_update_80978[4];
  assign array_update_80991[5] = add_80123 == 32'h0000_0005 ? array_update_80989 : array_update_80978[5];
  assign array_update_80991[6] = add_80123 == 32'h0000_0006 ? array_update_80989 : array_update_80978[6];
  assign array_update_80991[7] = add_80123 == 32'h0000_0007 ? array_update_80989 : array_update_80978[7];
  assign array_update_80991[8] = add_80123 == 32'h0000_0008 ? array_update_80989 : array_update_80978[8];
  assign array_update_80991[9] = add_80123 == 32'h0000_0009 ? array_update_80989 : array_update_80978[9];
  assign array_index_80993 = array_update_72021[add_80990 > 32'h0000_0009 ? 4'h9 : add_80990[3:0]];
  assign array_index_80994 = array_update_80991[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_80998 = smul32b_32b_x_32b(array_index_80130[add_80990 > 32'h0000_0009 ? 4'h9 : add_80990[3:0]], array_index_80993[add_80936 > 32'h0000_0009 ? 4'h9 : add_80936[3:0]]);
  assign add_81000 = array_index_80994[add_80936 > 32'h0000_0009 ? 4'h9 : add_80936[3:0]] + smul_80998;
  assign array_update_81002[0] = add_80936 == 32'h0000_0000 ? add_81000 : array_index_80994[0];
  assign array_update_81002[1] = add_80936 == 32'h0000_0001 ? add_81000 : array_index_80994[1];
  assign array_update_81002[2] = add_80936 == 32'h0000_0002 ? add_81000 : array_index_80994[2];
  assign array_update_81002[3] = add_80936 == 32'h0000_0003 ? add_81000 : array_index_80994[3];
  assign array_update_81002[4] = add_80936 == 32'h0000_0004 ? add_81000 : array_index_80994[4];
  assign array_update_81002[5] = add_80936 == 32'h0000_0005 ? add_81000 : array_index_80994[5];
  assign array_update_81002[6] = add_80936 == 32'h0000_0006 ? add_81000 : array_index_80994[6];
  assign array_update_81002[7] = add_80936 == 32'h0000_0007 ? add_81000 : array_index_80994[7];
  assign array_update_81002[8] = add_80936 == 32'h0000_0008 ? add_81000 : array_index_80994[8];
  assign array_update_81002[9] = add_80936 == 32'h0000_0009 ? add_81000 : array_index_80994[9];
  assign add_81003 = add_80990 + 32'h0000_0001;
  assign array_update_81004[0] = add_80123 == 32'h0000_0000 ? array_update_81002 : array_update_80991[0];
  assign array_update_81004[1] = add_80123 == 32'h0000_0001 ? array_update_81002 : array_update_80991[1];
  assign array_update_81004[2] = add_80123 == 32'h0000_0002 ? array_update_81002 : array_update_80991[2];
  assign array_update_81004[3] = add_80123 == 32'h0000_0003 ? array_update_81002 : array_update_80991[3];
  assign array_update_81004[4] = add_80123 == 32'h0000_0004 ? array_update_81002 : array_update_80991[4];
  assign array_update_81004[5] = add_80123 == 32'h0000_0005 ? array_update_81002 : array_update_80991[5];
  assign array_update_81004[6] = add_80123 == 32'h0000_0006 ? array_update_81002 : array_update_80991[6];
  assign array_update_81004[7] = add_80123 == 32'h0000_0007 ? array_update_81002 : array_update_80991[7];
  assign array_update_81004[8] = add_80123 == 32'h0000_0008 ? array_update_81002 : array_update_80991[8];
  assign array_update_81004[9] = add_80123 == 32'h0000_0009 ? array_update_81002 : array_update_80991[9];
  assign array_index_81006 = array_update_72021[add_81003 > 32'h0000_0009 ? 4'h9 : add_81003[3:0]];
  assign array_index_81007 = array_update_81004[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_81011 = smul32b_32b_x_32b(array_index_80130[add_81003 > 32'h0000_0009 ? 4'h9 : add_81003[3:0]], array_index_81006[add_80936 > 32'h0000_0009 ? 4'h9 : add_80936[3:0]]);
  assign add_81013 = array_index_81007[add_80936 > 32'h0000_0009 ? 4'h9 : add_80936[3:0]] + smul_81011;
  assign array_update_81015[0] = add_80936 == 32'h0000_0000 ? add_81013 : array_index_81007[0];
  assign array_update_81015[1] = add_80936 == 32'h0000_0001 ? add_81013 : array_index_81007[1];
  assign array_update_81015[2] = add_80936 == 32'h0000_0002 ? add_81013 : array_index_81007[2];
  assign array_update_81015[3] = add_80936 == 32'h0000_0003 ? add_81013 : array_index_81007[3];
  assign array_update_81015[4] = add_80936 == 32'h0000_0004 ? add_81013 : array_index_81007[4];
  assign array_update_81015[5] = add_80936 == 32'h0000_0005 ? add_81013 : array_index_81007[5];
  assign array_update_81015[6] = add_80936 == 32'h0000_0006 ? add_81013 : array_index_81007[6];
  assign array_update_81015[7] = add_80936 == 32'h0000_0007 ? add_81013 : array_index_81007[7];
  assign array_update_81015[8] = add_80936 == 32'h0000_0008 ? add_81013 : array_index_81007[8];
  assign array_update_81015[9] = add_80936 == 32'h0000_0009 ? add_81013 : array_index_81007[9];
  assign add_81016 = add_81003 + 32'h0000_0001;
  assign array_update_81017[0] = add_80123 == 32'h0000_0000 ? array_update_81015 : array_update_81004[0];
  assign array_update_81017[1] = add_80123 == 32'h0000_0001 ? array_update_81015 : array_update_81004[1];
  assign array_update_81017[2] = add_80123 == 32'h0000_0002 ? array_update_81015 : array_update_81004[2];
  assign array_update_81017[3] = add_80123 == 32'h0000_0003 ? array_update_81015 : array_update_81004[3];
  assign array_update_81017[4] = add_80123 == 32'h0000_0004 ? array_update_81015 : array_update_81004[4];
  assign array_update_81017[5] = add_80123 == 32'h0000_0005 ? array_update_81015 : array_update_81004[5];
  assign array_update_81017[6] = add_80123 == 32'h0000_0006 ? array_update_81015 : array_update_81004[6];
  assign array_update_81017[7] = add_80123 == 32'h0000_0007 ? array_update_81015 : array_update_81004[7];
  assign array_update_81017[8] = add_80123 == 32'h0000_0008 ? array_update_81015 : array_update_81004[8];
  assign array_update_81017[9] = add_80123 == 32'h0000_0009 ? array_update_81015 : array_update_81004[9];
  assign array_index_81019 = array_update_72021[add_81016 > 32'h0000_0009 ? 4'h9 : add_81016[3:0]];
  assign array_index_81020 = array_update_81017[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_81024 = smul32b_32b_x_32b(array_index_80130[add_81016 > 32'h0000_0009 ? 4'h9 : add_81016[3:0]], array_index_81019[add_80936 > 32'h0000_0009 ? 4'h9 : add_80936[3:0]]);
  assign add_81026 = array_index_81020[add_80936 > 32'h0000_0009 ? 4'h9 : add_80936[3:0]] + smul_81024;
  assign array_update_81028[0] = add_80936 == 32'h0000_0000 ? add_81026 : array_index_81020[0];
  assign array_update_81028[1] = add_80936 == 32'h0000_0001 ? add_81026 : array_index_81020[1];
  assign array_update_81028[2] = add_80936 == 32'h0000_0002 ? add_81026 : array_index_81020[2];
  assign array_update_81028[3] = add_80936 == 32'h0000_0003 ? add_81026 : array_index_81020[3];
  assign array_update_81028[4] = add_80936 == 32'h0000_0004 ? add_81026 : array_index_81020[4];
  assign array_update_81028[5] = add_80936 == 32'h0000_0005 ? add_81026 : array_index_81020[5];
  assign array_update_81028[6] = add_80936 == 32'h0000_0006 ? add_81026 : array_index_81020[6];
  assign array_update_81028[7] = add_80936 == 32'h0000_0007 ? add_81026 : array_index_81020[7];
  assign array_update_81028[8] = add_80936 == 32'h0000_0008 ? add_81026 : array_index_81020[8];
  assign array_update_81028[9] = add_80936 == 32'h0000_0009 ? add_81026 : array_index_81020[9];
  assign add_81029 = add_81016 + 32'h0000_0001;
  assign array_update_81030[0] = add_80123 == 32'h0000_0000 ? array_update_81028 : array_update_81017[0];
  assign array_update_81030[1] = add_80123 == 32'h0000_0001 ? array_update_81028 : array_update_81017[1];
  assign array_update_81030[2] = add_80123 == 32'h0000_0002 ? array_update_81028 : array_update_81017[2];
  assign array_update_81030[3] = add_80123 == 32'h0000_0003 ? array_update_81028 : array_update_81017[3];
  assign array_update_81030[4] = add_80123 == 32'h0000_0004 ? array_update_81028 : array_update_81017[4];
  assign array_update_81030[5] = add_80123 == 32'h0000_0005 ? array_update_81028 : array_update_81017[5];
  assign array_update_81030[6] = add_80123 == 32'h0000_0006 ? array_update_81028 : array_update_81017[6];
  assign array_update_81030[7] = add_80123 == 32'h0000_0007 ? array_update_81028 : array_update_81017[7];
  assign array_update_81030[8] = add_80123 == 32'h0000_0008 ? array_update_81028 : array_update_81017[8];
  assign array_update_81030[9] = add_80123 == 32'h0000_0009 ? array_update_81028 : array_update_81017[9];
  assign array_index_81032 = array_update_72021[add_81029 > 32'h0000_0009 ? 4'h9 : add_81029[3:0]];
  assign array_index_81033 = array_update_81030[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_81037 = smul32b_32b_x_32b(array_index_80130[add_81029 > 32'h0000_0009 ? 4'h9 : add_81029[3:0]], array_index_81032[add_80936 > 32'h0000_0009 ? 4'h9 : add_80936[3:0]]);
  assign add_81039 = array_index_81033[add_80936 > 32'h0000_0009 ? 4'h9 : add_80936[3:0]] + smul_81037;
  assign array_update_81041[0] = add_80936 == 32'h0000_0000 ? add_81039 : array_index_81033[0];
  assign array_update_81041[1] = add_80936 == 32'h0000_0001 ? add_81039 : array_index_81033[1];
  assign array_update_81041[2] = add_80936 == 32'h0000_0002 ? add_81039 : array_index_81033[2];
  assign array_update_81041[3] = add_80936 == 32'h0000_0003 ? add_81039 : array_index_81033[3];
  assign array_update_81041[4] = add_80936 == 32'h0000_0004 ? add_81039 : array_index_81033[4];
  assign array_update_81041[5] = add_80936 == 32'h0000_0005 ? add_81039 : array_index_81033[5];
  assign array_update_81041[6] = add_80936 == 32'h0000_0006 ? add_81039 : array_index_81033[6];
  assign array_update_81041[7] = add_80936 == 32'h0000_0007 ? add_81039 : array_index_81033[7];
  assign array_update_81041[8] = add_80936 == 32'h0000_0008 ? add_81039 : array_index_81033[8];
  assign array_update_81041[9] = add_80936 == 32'h0000_0009 ? add_81039 : array_index_81033[9];
  assign add_81042 = add_81029 + 32'h0000_0001;
  assign array_update_81043[0] = add_80123 == 32'h0000_0000 ? array_update_81041 : array_update_81030[0];
  assign array_update_81043[1] = add_80123 == 32'h0000_0001 ? array_update_81041 : array_update_81030[1];
  assign array_update_81043[2] = add_80123 == 32'h0000_0002 ? array_update_81041 : array_update_81030[2];
  assign array_update_81043[3] = add_80123 == 32'h0000_0003 ? array_update_81041 : array_update_81030[3];
  assign array_update_81043[4] = add_80123 == 32'h0000_0004 ? array_update_81041 : array_update_81030[4];
  assign array_update_81043[5] = add_80123 == 32'h0000_0005 ? array_update_81041 : array_update_81030[5];
  assign array_update_81043[6] = add_80123 == 32'h0000_0006 ? array_update_81041 : array_update_81030[6];
  assign array_update_81043[7] = add_80123 == 32'h0000_0007 ? array_update_81041 : array_update_81030[7];
  assign array_update_81043[8] = add_80123 == 32'h0000_0008 ? array_update_81041 : array_update_81030[8];
  assign array_update_81043[9] = add_80123 == 32'h0000_0009 ? array_update_81041 : array_update_81030[9];
  assign array_index_81045 = array_update_72021[add_81042 > 32'h0000_0009 ? 4'h9 : add_81042[3:0]];
  assign array_index_81046 = array_update_81043[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_81050 = smul32b_32b_x_32b(array_index_80130[add_81042 > 32'h0000_0009 ? 4'h9 : add_81042[3:0]], array_index_81045[add_80936 > 32'h0000_0009 ? 4'h9 : add_80936[3:0]]);
  assign add_81052 = array_index_81046[add_80936 > 32'h0000_0009 ? 4'h9 : add_80936[3:0]] + smul_81050;
  assign array_update_81054[0] = add_80936 == 32'h0000_0000 ? add_81052 : array_index_81046[0];
  assign array_update_81054[1] = add_80936 == 32'h0000_0001 ? add_81052 : array_index_81046[1];
  assign array_update_81054[2] = add_80936 == 32'h0000_0002 ? add_81052 : array_index_81046[2];
  assign array_update_81054[3] = add_80936 == 32'h0000_0003 ? add_81052 : array_index_81046[3];
  assign array_update_81054[4] = add_80936 == 32'h0000_0004 ? add_81052 : array_index_81046[4];
  assign array_update_81054[5] = add_80936 == 32'h0000_0005 ? add_81052 : array_index_81046[5];
  assign array_update_81054[6] = add_80936 == 32'h0000_0006 ? add_81052 : array_index_81046[6];
  assign array_update_81054[7] = add_80936 == 32'h0000_0007 ? add_81052 : array_index_81046[7];
  assign array_update_81054[8] = add_80936 == 32'h0000_0008 ? add_81052 : array_index_81046[8];
  assign array_update_81054[9] = add_80936 == 32'h0000_0009 ? add_81052 : array_index_81046[9];
  assign add_81055 = add_81042 + 32'h0000_0001;
  assign array_update_81056[0] = add_80123 == 32'h0000_0000 ? array_update_81054 : array_update_81043[0];
  assign array_update_81056[1] = add_80123 == 32'h0000_0001 ? array_update_81054 : array_update_81043[1];
  assign array_update_81056[2] = add_80123 == 32'h0000_0002 ? array_update_81054 : array_update_81043[2];
  assign array_update_81056[3] = add_80123 == 32'h0000_0003 ? array_update_81054 : array_update_81043[3];
  assign array_update_81056[4] = add_80123 == 32'h0000_0004 ? array_update_81054 : array_update_81043[4];
  assign array_update_81056[5] = add_80123 == 32'h0000_0005 ? array_update_81054 : array_update_81043[5];
  assign array_update_81056[6] = add_80123 == 32'h0000_0006 ? array_update_81054 : array_update_81043[6];
  assign array_update_81056[7] = add_80123 == 32'h0000_0007 ? array_update_81054 : array_update_81043[7];
  assign array_update_81056[8] = add_80123 == 32'h0000_0008 ? array_update_81054 : array_update_81043[8];
  assign array_update_81056[9] = add_80123 == 32'h0000_0009 ? array_update_81054 : array_update_81043[9];
  assign array_index_81058 = array_update_72021[add_81055 > 32'h0000_0009 ? 4'h9 : add_81055[3:0]];
  assign array_index_81059 = array_update_81056[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_81063 = smul32b_32b_x_32b(array_index_80130[add_81055 > 32'h0000_0009 ? 4'h9 : add_81055[3:0]], array_index_81058[add_80936 > 32'h0000_0009 ? 4'h9 : add_80936[3:0]]);
  assign add_81065 = array_index_81059[add_80936 > 32'h0000_0009 ? 4'h9 : add_80936[3:0]] + smul_81063;
  assign array_update_81066[0] = add_80936 == 32'h0000_0000 ? add_81065 : array_index_81059[0];
  assign array_update_81066[1] = add_80936 == 32'h0000_0001 ? add_81065 : array_index_81059[1];
  assign array_update_81066[2] = add_80936 == 32'h0000_0002 ? add_81065 : array_index_81059[2];
  assign array_update_81066[3] = add_80936 == 32'h0000_0003 ? add_81065 : array_index_81059[3];
  assign array_update_81066[4] = add_80936 == 32'h0000_0004 ? add_81065 : array_index_81059[4];
  assign array_update_81066[5] = add_80936 == 32'h0000_0005 ? add_81065 : array_index_81059[5];
  assign array_update_81066[6] = add_80936 == 32'h0000_0006 ? add_81065 : array_index_81059[6];
  assign array_update_81066[7] = add_80936 == 32'h0000_0007 ? add_81065 : array_index_81059[7];
  assign array_update_81066[8] = add_80936 == 32'h0000_0008 ? add_81065 : array_index_81059[8];
  assign array_update_81066[9] = add_80936 == 32'h0000_0009 ? add_81065 : array_index_81059[9];
  assign array_update_81067[0] = add_80123 == 32'h0000_0000 ? array_update_81066 : array_update_81056[0];
  assign array_update_81067[1] = add_80123 == 32'h0000_0001 ? array_update_81066 : array_update_81056[1];
  assign array_update_81067[2] = add_80123 == 32'h0000_0002 ? array_update_81066 : array_update_81056[2];
  assign array_update_81067[3] = add_80123 == 32'h0000_0003 ? array_update_81066 : array_update_81056[3];
  assign array_update_81067[4] = add_80123 == 32'h0000_0004 ? array_update_81066 : array_update_81056[4];
  assign array_update_81067[5] = add_80123 == 32'h0000_0005 ? array_update_81066 : array_update_81056[5];
  assign array_update_81067[6] = add_80123 == 32'h0000_0006 ? array_update_81066 : array_update_81056[6];
  assign array_update_81067[7] = add_80123 == 32'h0000_0007 ? array_update_81066 : array_update_81056[7];
  assign array_update_81067[8] = add_80123 == 32'h0000_0008 ? array_update_81066 : array_update_81056[8];
  assign array_update_81067[9] = add_80123 == 32'h0000_0009 ? array_update_81066 : array_update_81056[9];
  assign array_index_81069 = array_update_81067[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign add_81071 = add_80936 + 32'h0000_0001;
  assign array_update_81072[0] = add_81071 == 32'h0000_0000 ? 32'h0000_0000 : array_index_81069[0];
  assign array_update_81072[1] = add_81071 == 32'h0000_0001 ? 32'h0000_0000 : array_index_81069[1];
  assign array_update_81072[2] = add_81071 == 32'h0000_0002 ? 32'h0000_0000 : array_index_81069[2];
  assign array_update_81072[3] = add_81071 == 32'h0000_0003 ? 32'h0000_0000 : array_index_81069[3];
  assign array_update_81072[4] = add_81071 == 32'h0000_0004 ? 32'h0000_0000 : array_index_81069[4];
  assign array_update_81072[5] = add_81071 == 32'h0000_0005 ? 32'h0000_0000 : array_index_81069[5];
  assign array_update_81072[6] = add_81071 == 32'h0000_0006 ? 32'h0000_0000 : array_index_81069[6];
  assign array_update_81072[7] = add_81071 == 32'h0000_0007 ? 32'h0000_0000 : array_index_81069[7];
  assign array_update_81072[8] = add_81071 == 32'h0000_0008 ? 32'h0000_0000 : array_index_81069[8];
  assign array_update_81072[9] = add_81071 == 32'h0000_0009 ? 32'h0000_0000 : array_index_81069[9];
  assign literal_81073 = 32'h0000_0000;
  assign array_update_81074[0] = add_80123 == 32'h0000_0000 ? array_update_81072 : array_update_81067[0];
  assign array_update_81074[1] = add_80123 == 32'h0000_0001 ? array_update_81072 : array_update_81067[1];
  assign array_update_81074[2] = add_80123 == 32'h0000_0002 ? array_update_81072 : array_update_81067[2];
  assign array_update_81074[3] = add_80123 == 32'h0000_0003 ? array_update_81072 : array_update_81067[3];
  assign array_update_81074[4] = add_80123 == 32'h0000_0004 ? array_update_81072 : array_update_81067[4];
  assign array_update_81074[5] = add_80123 == 32'h0000_0005 ? array_update_81072 : array_update_81067[5];
  assign array_update_81074[6] = add_80123 == 32'h0000_0006 ? array_update_81072 : array_update_81067[6];
  assign array_update_81074[7] = add_80123 == 32'h0000_0007 ? array_update_81072 : array_update_81067[7];
  assign array_update_81074[8] = add_80123 == 32'h0000_0008 ? array_update_81072 : array_update_81067[8];
  assign array_update_81074[9] = add_80123 == 32'h0000_0009 ? array_update_81072 : array_update_81067[9];
  assign array_index_81076 = array_update_72021[literal_81073 > 32'h0000_0009 ? 4'h9 : literal_81073[3:0]];
  assign array_index_81077 = array_update_81074[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_81081 = smul32b_32b_x_32b(array_index_80130[literal_81073 > 32'h0000_0009 ? 4'h9 : literal_81073[3:0]], array_index_81076[add_81071 > 32'h0000_0009 ? 4'h9 : add_81071[3:0]]);
  assign add_81083 = array_index_81077[add_81071 > 32'h0000_0009 ? 4'h9 : add_81071[3:0]] + smul_81081;
  assign array_update_81085[0] = add_81071 == 32'h0000_0000 ? add_81083 : array_index_81077[0];
  assign array_update_81085[1] = add_81071 == 32'h0000_0001 ? add_81083 : array_index_81077[1];
  assign array_update_81085[2] = add_81071 == 32'h0000_0002 ? add_81083 : array_index_81077[2];
  assign array_update_81085[3] = add_81071 == 32'h0000_0003 ? add_81083 : array_index_81077[3];
  assign array_update_81085[4] = add_81071 == 32'h0000_0004 ? add_81083 : array_index_81077[4];
  assign array_update_81085[5] = add_81071 == 32'h0000_0005 ? add_81083 : array_index_81077[5];
  assign array_update_81085[6] = add_81071 == 32'h0000_0006 ? add_81083 : array_index_81077[6];
  assign array_update_81085[7] = add_81071 == 32'h0000_0007 ? add_81083 : array_index_81077[7];
  assign array_update_81085[8] = add_81071 == 32'h0000_0008 ? add_81083 : array_index_81077[8];
  assign array_update_81085[9] = add_81071 == 32'h0000_0009 ? add_81083 : array_index_81077[9];
  assign add_81086 = literal_81073 + 32'h0000_0001;
  assign array_update_81087[0] = add_80123 == 32'h0000_0000 ? array_update_81085 : array_update_81074[0];
  assign array_update_81087[1] = add_80123 == 32'h0000_0001 ? array_update_81085 : array_update_81074[1];
  assign array_update_81087[2] = add_80123 == 32'h0000_0002 ? array_update_81085 : array_update_81074[2];
  assign array_update_81087[3] = add_80123 == 32'h0000_0003 ? array_update_81085 : array_update_81074[3];
  assign array_update_81087[4] = add_80123 == 32'h0000_0004 ? array_update_81085 : array_update_81074[4];
  assign array_update_81087[5] = add_80123 == 32'h0000_0005 ? array_update_81085 : array_update_81074[5];
  assign array_update_81087[6] = add_80123 == 32'h0000_0006 ? array_update_81085 : array_update_81074[6];
  assign array_update_81087[7] = add_80123 == 32'h0000_0007 ? array_update_81085 : array_update_81074[7];
  assign array_update_81087[8] = add_80123 == 32'h0000_0008 ? array_update_81085 : array_update_81074[8];
  assign array_update_81087[9] = add_80123 == 32'h0000_0009 ? array_update_81085 : array_update_81074[9];
  assign array_index_81089 = array_update_72021[add_81086 > 32'h0000_0009 ? 4'h9 : add_81086[3:0]];
  assign array_index_81090 = array_update_81087[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_81094 = smul32b_32b_x_32b(array_index_80130[add_81086 > 32'h0000_0009 ? 4'h9 : add_81086[3:0]], array_index_81089[add_81071 > 32'h0000_0009 ? 4'h9 : add_81071[3:0]]);
  assign add_81096 = array_index_81090[add_81071 > 32'h0000_0009 ? 4'h9 : add_81071[3:0]] + smul_81094;
  assign array_update_81098[0] = add_81071 == 32'h0000_0000 ? add_81096 : array_index_81090[0];
  assign array_update_81098[1] = add_81071 == 32'h0000_0001 ? add_81096 : array_index_81090[1];
  assign array_update_81098[2] = add_81071 == 32'h0000_0002 ? add_81096 : array_index_81090[2];
  assign array_update_81098[3] = add_81071 == 32'h0000_0003 ? add_81096 : array_index_81090[3];
  assign array_update_81098[4] = add_81071 == 32'h0000_0004 ? add_81096 : array_index_81090[4];
  assign array_update_81098[5] = add_81071 == 32'h0000_0005 ? add_81096 : array_index_81090[5];
  assign array_update_81098[6] = add_81071 == 32'h0000_0006 ? add_81096 : array_index_81090[6];
  assign array_update_81098[7] = add_81071 == 32'h0000_0007 ? add_81096 : array_index_81090[7];
  assign array_update_81098[8] = add_81071 == 32'h0000_0008 ? add_81096 : array_index_81090[8];
  assign array_update_81098[9] = add_81071 == 32'h0000_0009 ? add_81096 : array_index_81090[9];
  assign add_81099 = add_81086 + 32'h0000_0001;
  assign array_update_81100[0] = add_80123 == 32'h0000_0000 ? array_update_81098 : array_update_81087[0];
  assign array_update_81100[1] = add_80123 == 32'h0000_0001 ? array_update_81098 : array_update_81087[1];
  assign array_update_81100[2] = add_80123 == 32'h0000_0002 ? array_update_81098 : array_update_81087[2];
  assign array_update_81100[3] = add_80123 == 32'h0000_0003 ? array_update_81098 : array_update_81087[3];
  assign array_update_81100[4] = add_80123 == 32'h0000_0004 ? array_update_81098 : array_update_81087[4];
  assign array_update_81100[5] = add_80123 == 32'h0000_0005 ? array_update_81098 : array_update_81087[5];
  assign array_update_81100[6] = add_80123 == 32'h0000_0006 ? array_update_81098 : array_update_81087[6];
  assign array_update_81100[7] = add_80123 == 32'h0000_0007 ? array_update_81098 : array_update_81087[7];
  assign array_update_81100[8] = add_80123 == 32'h0000_0008 ? array_update_81098 : array_update_81087[8];
  assign array_update_81100[9] = add_80123 == 32'h0000_0009 ? array_update_81098 : array_update_81087[9];
  assign array_index_81102 = array_update_72021[add_81099 > 32'h0000_0009 ? 4'h9 : add_81099[3:0]];
  assign array_index_81103 = array_update_81100[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_81107 = smul32b_32b_x_32b(array_index_80130[add_81099 > 32'h0000_0009 ? 4'h9 : add_81099[3:0]], array_index_81102[add_81071 > 32'h0000_0009 ? 4'h9 : add_81071[3:0]]);
  assign add_81109 = array_index_81103[add_81071 > 32'h0000_0009 ? 4'h9 : add_81071[3:0]] + smul_81107;
  assign array_update_81111[0] = add_81071 == 32'h0000_0000 ? add_81109 : array_index_81103[0];
  assign array_update_81111[1] = add_81071 == 32'h0000_0001 ? add_81109 : array_index_81103[1];
  assign array_update_81111[2] = add_81071 == 32'h0000_0002 ? add_81109 : array_index_81103[2];
  assign array_update_81111[3] = add_81071 == 32'h0000_0003 ? add_81109 : array_index_81103[3];
  assign array_update_81111[4] = add_81071 == 32'h0000_0004 ? add_81109 : array_index_81103[4];
  assign array_update_81111[5] = add_81071 == 32'h0000_0005 ? add_81109 : array_index_81103[5];
  assign array_update_81111[6] = add_81071 == 32'h0000_0006 ? add_81109 : array_index_81103[6];
  assign array_update_81111[7] = add_81071 == 32'h0000_0007 ? add_81109 : array_index_81103[7];
  assign array_update_81111[8] = add_81071 == 32'h0000_0008 ? add_81109 : array_index_81103[8];
  assign array_update_81111[9] = add_81071 == 32'h0000_0009 ? add_81109 : array_index_81103[9];
  assign add_81112 = add_81099 + 32'h0000_0001;
  assign array_update_81113[0] = add_80123 == 32'h0000_0000 ? array_update_81111 : array_update_81100[0];
  assign array_update_81113[1] = add_80123 == 32'h0000_0001 ? array_update_81111 : array_update_81100[1];
  assign array_update_81113[2] = add_80123 == 32'h0000_0002 ? array_update_81111 : array_update_81100[2];
  assign array_update_81113[3] = add_80123 == 32'h0000_0003 ? array_update_81111 : array_update_81100[3];
  assign array_update_81113[4] = add_80123 == 32'h0000_0004 ? array_update_81111 : array_update_81100[4];
  assign array_update_81113[5] = add_80123 == 32'h0000_0005 ? array_update_81111 : array_update_81100[5];
  assign array_update_81113[6] = add_80123 == 32'h0000_0006 ? array_update_81111 : array_update_81100[6];
  assign array_update_81113[7] = add_80123 == 32'h0000_0007 ? array_update_81111 : array_update_81100[7];
  assign array_update_81113[8] = add_80123 == 32'h0000_0008 ? array_update_81111 : array_update_81100[8];
  assign array_update_81113[9] = add_80123 == 32'h0000_0009 ? array_update_81111 : array_update_81100[9];
  assign array_index_81115 = array_update_72021[add_81112 > 32'h0000_0009 ? 4'h9 : add_81112[3:0]];
  assign array_index_81116 = array_update_81113[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_81120 = smul32b_32b_x_32b(array_index_80130[add_81112 > 32'h0000_0009 ? 4'h9 : add_81112[3:0]], array_index_81115[add_81071 > 32'h0000_0009 ? 4'h9 : add_81071[3:0]]);
  assign add_81122 = array_index_81116[add_81071 > 32'h0000_0009 ? 4'h9 : add_81071[3:0]] + smul_81120;
  assign array_update_81124[0] = add_81071 == 32'h0000_0000 ? add_81122 : array_index_81116[0];
  assign array_update_81124[1] = add_81071 == 32'h0000_0001 ? add_81122 : array_index_81116[1];
  assign array_update_81124[2] = add_81071 == 32'h0000_0002 ? add_81122 : array_index_81116[2];
  assign array_update_81124[3] = add_81071 == 32'h0000_0003 ? add_81122 : array_index_81116[3];
  assign array_update_81124[4] = add_81071 == 32'h0000_0004 ? add_81122 : array_index_81116[4];
  assign array_update_81124[5] = add_81071 == 32'h0000_0005 ? add_81122 : array_index_81116[5];
  assign array_update_81124[6] = add_81071 == 32'h0000_0006 ? add_81122 : array_index_81116[6];
  assign array_update_81124[7] = add_81071 == 32'h0000_0007 ? add_81122 : array_index_81116[7];
  assign array_update_81124[8] = add_81071 == 32'h0000_0008 ? add_81122 : array_index_81116[8];
  assign array_update_81124[9] = add_81071 == 32'h0000_0009 ? add_81122 : array_index_81116[9];
  assign add_81125 = add_81112 + 32'h0000_0001;
  assign array_update_81126[0] = add_80123 == 32'h0000_0000 ? array_update_81124 : array_update_81113[0];
  assign array_update_81126[1] = add_80123 == 32'h0000_0001 ? array_update_81124 : array_update_81113[1];
  assign array_update_81126[2] = add_80123 == 32'h0000_0002 ? array_update_81124 : array_update_81113[2];
  assign array_update_81126[3] = add_80123 == 32'h0000_0003 ? array_update_81124 : array_update_81113[3];
  assign array_update_81126[4] = add_80123 == 32'h0000_0004 ? array_update_81124 : array_update_81113[4];
  assign array_update_81126[5] = add_80123 == 32'h0000_0005 ? array_update_81124 : array_update_81113[5];
  assign array_update_81126[6] = add_80123 == 32'h0000_0006 ? array_update_81124 : array_update_81113[6];
  assign array_update_81126[7] = add_80123 == 32'h0000_0007 ? array_update_81124 : array_update_81113[7];
  assign array_update_81126[8] = add_80123 == 32'h0000_0008 ? array_update_81124 : array_update_81113[8];
  assign array_update_81126[9] = add_80123 == 32'h0000_0009 ? array_update_81124 : array_update_81113[9];
  assign array_index_81128 = array_update_72021[add_81125 > 32'h0000_0009 ? 4'h9 : add_81125[3:0]];
  assign array_index_81129 = array_update_81126[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_81133 = smul32b_32b_x_32b(array_index_80130[add_81125 > 32'h0000_0009 ? 4'h9 : add_81125[3:0]], array_index_81128[add_81071 > 32'h0000_0009 ? 4'h9 : add_81071[3:0]]);
  assign add_81135 = array_index_81129[add_81071 > 32'h0000_0009 ? 4'h9 : add_81071[3:0]] + smul_81133;
  assign array_update_81137[0] = add_81071 == 32'h0000_0000 ? add_81135 : array_index_81129[0];
  assign array_update_81137[1] = add_81071 == 32'h0000_0001 ? add_81135 : array_index_81129[1];
  assign array_update_81137[2] = add_81071 == 32'h0000_0002 ? add_81135 : array_index_81129[2];
  assign array_update_81137[3] = add_81071 == 32'h0000_0003 ? add_81135 : array_index_81129[3];
  assign array_update_81137[4] = add_81071 == 32'h0000_0004 ? add_81135 : array_index_81129[4];
  assign array_update_81137[5] = add_81071 == 32'h0000_0005 ? add_81135 : array_index_81129[5];
  assign array_update_81137[6] = add_81071 == 32'h0000_0006 ? add_81135 : array_index_81129[6];
  assign array_update_81137[7] = add_81071 == 32'h0000_0007 ? add_81135 : array_index_81129[7];
  assign array_update_81137[8] = add_81071 == 32'h0000_0008 ? add_81135 : array_index_81129[8];
  assign array_update_81137[9] = add_81071 == 32'h0000_0009 ? add_81135 : array_index_81129[9];
  assign add_81138 = add_81125 + 32'h0000_0001;
  assign array_update_81139[0] = add_80123 == 32'h0000_0000 ? array_update_81137 : array_update_81126[0];
  assign array_update_81139[1] = add_80123 == 32'h0000_0001 ? array_update_81137 : array_update_81126[1];
  assign array_update_81139[2] = add_80123 == 32'h0000_0002 ? array_update_81137 : array_update_81126[2];
  assign array_update_81139[3] = add_80123 == 32'h0000_0003 ? array_update_81137 : array_update_81126[3];
  assign array_update_81139[4] = add_80123 == 32'h0000_0004 ? array_update_81137 : array_update_81126[4];
  assign array_update_81139[5] = add_80123 == 32'h0000_0005 ? array_update_81137 : array_update_81126[5];
  assign array_update_81139[6] = add_80123 == 32'h0000_0006 ? array_update_81137 : array_update_81126[6];
  assign array_update_81139[7] = add_80123 == 32'h0000_0007 ? array_update_81137 : array_update_81126[7];
  assign array_update_81139[8] = add_80123 == 32'h0000_0008 ? array_update_81137 : array_update_81126[8];
  assign array_update_81139[9] = add_80123 == 32'h0000_0009 ? array_update_81137 : array_update_81126[9];
  assign array_index_81141 = array_update_72021[add_81138 > 32'h0000_0009 ? 4'h9 : add_81138[3:0]];
  assign array_index_81142 = array_update_81139[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_81146 = smul32b_32b_x_32b(array_index_80130[add_81138 > 32'h0000_0009 ? 4'h9 : add_81138[3:0]], array_index_81141[add_81071 > 32'h0000_0009 ? 4'h9 : add_81071[3:0]]);
  assign add_81148 = array_index_81142[add_81071 > 32'h0000_0009 ? 4'h9 : add_81071[3:0]] + smul_81146;
  assign array_update_81150[0] = add_81071 == 32'h0000_0000 ? add_81148 : array_index_81142[0];
  assign array_update_81150[1] = add_81071 == 32'h0000_0001 ? add_81148 : array_index_81142[1];
  assign array_update_81150[2] = add_81071 == 32'h0000_0002 ? add_81148 : array_index_81142[2];
  assign array_update_81150[3] = add_81071 == 32'h0000_0003 ? add_81148 : array_index_81142[3];
  assign array_update_81150[4] = add_81071 == 32'h0000_0004 ? add_81148 : array_index_81142[4];
  assign array_update_81150[5] = add_81071 == 32'h0000_0005 ? add_81148 : array_index_81142[5];
  assign array_update_81150[6] = add_81071 == 32'h0000_0006 ? add_81148 : array_index_81142[6];
  assign array_update_81150[7] = add_81071 == 32'h0000_0007 ? add_81148 : array_index_81142[7];
  assign array_update_81150[8] = add_81071 == 32'h0000_0008 ? add_81148 : array_index_81142[8];
  assign array_update_81150[9] = add_81071 == 32'h0000_0009 ? add_81148 : array_index_81142[9];
  assign add_81151 = add_81138 + 32'h0000_0001;
  assign array_update_81152[0] = add_80123 == 32'h0000_0000 ? array_update_81150 : array_update_81139[0];
  assign array_update_81152[1] = add_80123 == 32'h0000_0001 ? array_update_81150 : array_update_81139[1];
  assign array_update_81152[2] = add_80123 == 32'h0000_0002 ? array_update_81150 : array_update_81139[2];
  assign array_update_81152[3] = add_80123 == 32'h0000_0003 ? array_update_81150 : array_update_81139[3];
  assign array_update_81152[4] = add_80123 == 32'h0000_0004 ? array_update_81150 : array_update_81139[4];
  assign array_update_81152[5] = add_80123 == 32'h0000_0005 ? array_update_81150 : array_update_81139[5];
  assign array_update_81152[6] = add_80123 == 32'h0000_0006 ? array_update_81150 : array_update_81139[6];
  assign array_update_81152[7] = add_80123 == 32'h0000_0007 ? array_update_81150 : array_update_81139[7];
  assign array_update_81152[8] = add_80123 == 32'h0000_0008 ? array_update_81150 : array_update_81139[8];
  assign array_update_81152[9] = add_80123 == 32'h0000_0009 ? array_update_81150 : array_update_81139[9];
  assign array_index_81154 = array_update_72021[add_81151 > 32'h0000_0009 ? 4'h9 : add_81151[3:0]];
  assign array_index_81155 = array_update_81152[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_81159 = smul32b_32b_x_32b(array_index_80130[add_81151 > 32'h0000_0009 ? 4'h9 : add_81151[3:0]], array_index_81154[add_81071 > 32'h0000_0009 ? 4'h9 : add_81071[3:0]]);
  assign add_81161 = array_index_81155[add_81071 > 32'h0000_0009 ? 4'h9 : add_81071[3:0]] + smul_81159;
  assign array_update_81163[0] = add_81071 == 32'h0000_0000 ? add_81161 : array_index_81155[0];
  assign array_update_81163[1] = add_81071 == 32'h0000_0001 ? add_81161 : array_index_81155[1];
  assign array_update_81163[2] = add_81071 == 32'h0000_0002 ? add_81161 : array_index_81155[2];
  assign array_update_81163[3] = add_81071 == 32'h0000_0003 ? add_81161 : array_index_81155[3];
  assign array_update_81163[4] = add_81071 == 32'h0000_0004 ? add_81161 : array_index_81155[4];
  assign array_update_81163[5] = add_81071 == 32'h0000_0005 ? add_81161 : array_index_81155[5];
  assign array_update_81163[6] = add_81071 == 32'h0000_0006 ? add_81161 : array_index_81155[6];
  assign array_update_81163[7] = add_81071 == 32'h0000_0007 ? add_81161 : array_index_81155[7];
  assign array_update_81163[8] = add_81071 == 32'h0000_0008 ? add_81161 : array_index_81155[8];
  assign array_update_81163[9] = add_81071 == 32'h0000_0009 ? add_81161 : array_index_81155[9];
  assign add_81164 = add_81151 + 32'h0000_0001;
  assign array_update_81165[0] = add_80123 == 32'h0000_0000 ? array_update_81163 : array_update_81152[0];
  assign array_update_81165[1] = add_80123 == 32'h0000_0001 ? array_update_81163 : array_update_81152[1];
  assign array_update_81165[2] = add_80123 == 32'h0000_0002 ? array_update_81163 : array_update_81152[2];
  assign array_update_81165[3] = add_80123 == 32'h0000_0003 ? array_update_81163 : array_update_81152[3];
  assign array_update_81165[4] = add_80123 == 32'h0000_0004 ? array_update_81163 : array_update_81152[4];
  assign array_update_81165[5] = add_80123 == 32'h0000_0005 ? array_update_81163 : array_update_81152[5];
  assign array_update_81165[6] = add_80123 == 32'h0000_0006 ? array_update_81163 : array_update_81152[6];
  assign array_update_81165[7] = add_80123 == 32'h0000_0007 ? array_update_81163 : array_update_81152[7];
  assign array_update_81165[8] = add_80123 == 32'h0000_0008 ? array_update_81163 : array_update_81152[8];
  assign array_update_81165[9] = add_80123 == 32'h0000_0009 ? array_update_81163 : array_update_81152[9];
  assign array_index_81167 = array_update_72021[add_81164 > 32'h0000_0009 ? 4'h9 : add_81164[3:0]];
  assign array_index_81168 = array_update_81165[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_81172 = smul32b_32b_x_32b(array_index_80130[add_81164 > 32'h0000_0009 ? 4'h9 : add_81164[3:0]], array_index_81167[add_81071 > 32'h0000_0009 ? 4'h9 : add_81071[3:0]]);
  assign add_81174 = array_index_81168[add_81071 > 32'h0000_0009 ? 4'h9 : add_81071[3:0]] + smul_81172;
  assign array_update_81176[0] = add_81071 == 32'h0000_0000 ? add_81174 : array_index_81168[0];
  assign array_update_81176[1] = add_81071 == 32'h0000_0001 ? add_81174 : array_index_81168[1];
  assign array_update_81176[2] = add_81071 == 32'h0000_0002 ? add_81174 : array_index_81168[2];
  assign array_update_81176[3] = add_81071 == 32'h0000_0003 ? add_81174 : array_index_81168[3];
  assign array_update_81176[4] = add_81071 == 32'h0000_0004 ? add_81174 : array_index_81168[4];
  assign array_update_81176[5] = add_81071 == 32'h0000_0005 ? add_81174 : array_index_81168[5];
  assign array_update_81176[6] = add_81071 == 32'h0000_0006 ? add_81174 : array_index_81168[6];
  assign array_update_81176[7] = add_81071 == 32'h0000_0007 ? add_81174 : array_index_81168[7];
  assign array_update_81176[8] = add_81071 == 32'h0000_0008 ? add_81174 : array_index_81168[8];
  assign array_update_81176[9] = add_81071 == 32'h0000_0009 ? add_81174 : array_index_81168[9];
  assign add_81177 = add_81164 + 32'h0000_0001;
  assign array_update_81178[0] = add_80123 == 32'h0000_0000 ? array_update_81176 : array_update_81165[0];
  assign array_update_81178[1] = add_80123 == 32'h0000_0001 ? array_update_81176 : array_update_81165[1];
  assign array_update_81178[2] = add_80123 == 32'h0000_0002 ? array_update_81176 : array_update_81165[2];
  assign array_update_81178[3] = add_80123 == 32'h0000_0003 ? array_update_81176 : array_update_81165[3];
  assign array_update_81178[4] = add_80123 == 32'h0000_0004 ? array_update_81176 : array_update_81165[4];
  assign array_update_81178[5] = add_80123 == 32'h0000_0005 ? array_update_81176 : array_update_81165[5];
  assign array_update_81178[6] = add_80123 == 32'h0000_0006 ? array_update_81176 : array_update_81165[6];
  assign array_update_81178[7] = add_80123 == 32'h0000_0007 ? array_update_81176 : array_update_81165[7];
  assign array_update_81178[8] = add_80123 == 32'h0000_0008 ? array_update_81176 : array_update_81165[8];
  assign array_update_81178[9] = add_80123 == 32'h0000_0009 ? array_update_81176 : array_update_81165[9];
  assign array_index_81180 = array_update_72021[add_81177 > 32'h0000_0009 ? 4'h9 : add_81177[3:0]];
  assign array_index_81181 = array_update_81178[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_81185 = smul32b_32b_x_32b(array_index_80130[add_81177 > 32'h0000_0009 ? 4'h9 : add_81177[3:0]], array_index_81180[add_81071 > 32'h0000_0009 ? 4'h9 : add_81071[3:0]]);
  assign add_81187 = array_index_81181[add_81071 > 32'h0000_0009 ? 4'h9 : add_81071[3:0]] + smul_81185;
  assign array_update_81189[0] = add_81071 == 32'h0000_0000 ? add_81187 : array_index_81181[0];
  assign array_update_81189[1] = add_81071 == 32'h0000_0001 ? add_81187 : array_index_81181[1];
  assign array_update_81189[2] = add_81071 == 32'h0000_0002 ? add_81187 : array_index_81181[2];
  assign array_update_81189[3] = add_81071 == 32'h0000_0003 ? add_81187 : array_index_81181[3];
  assign array_update_81189[4] = add_81071 == 32'h0000_0004 ? add_81187 : array_index_81181[4];
  assign array_update_81189[5] = add_81071 == 32'h0000_0005 ? add_81187 : array_index_81181[5];
  assign array_update_81189[6] = add_81071 == 32'h0000_0006 ? add_81187 : array_index_81181[6];
  assign array_update_81189[7] = add_81071 == 32'h0000_0007 ? add_81187 : array_index_81181[7];
  assign array_update_81189[8] = add_81071 == 32'h0000_0008 ? add_81187 : array_index_81181[8];
  assign array_update_81189[9] = add_81071 == 32'h0000_0009 ? add_81187 : array_index_81181[9];
  assign add_81190 = add_81177 + 32'h0000_0001;
  assign array_update_81191[0] = add_80123 == 32'h0000_0000 ? array_update_81189 : array_update_81178[0];
  assign array_update_81191[1] = add_80123 == 32'h0000_0001 ? array_update_81189 : array_update_81178[1];
  assign array_update_81191[2] = add_80123 == 32'h0000_0002 ? array_update_81189 : array_update_81178[2];
  assign array_update_81191[3] = add_80123 == 32'h0000_0003 ? array_update_81189 : array_update_81178[3];
  assign array_update_81191[4] = add_80123 == 32'h0000_0004 ? array_update_81189 : array_update_81178[4];
  assign array_update_81191[5] = add_80123 == 32'h0000_0005 ? array_update_81189 : array_update_81178[5];
  assign array_update_81191[6] = add_80123 == 32'h0000_0006 ? array_update_81189 : array_update_81178[6];
  assign array_update_81191[7] = add_80123 == 32'h0000_0007 ? array_update_81189 : array_update_81178[7];
  assign array_update_81191[8] = add_80123 == 32'h0000_0008 ? array_update_81189 : array_update_81178[8];
  assign array_update_81191[9] = add_80123 == 32'h0000_0009 ? array_update_81189 : array_update_81178[9];
  assign array_index_81193 = array_update_72021[add_81190 > 32'h0000_0009 ? 4'h9 : add_81190[3:0]];
  assign array_index_81194 = array_update_81191[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_81198 = smul32b_32b_x_32b(array_index_80130[add_81190 > 32'h0000_0009 ? 4'h9 : add_81190[3:0]], array_index_81193[add_81071 > 32'h0000_0009 ? 4'h9 : add_81071[3:0]]);
  assign add_81200 = array_index_81194[add_81071 > 32'h0000_0009 ? 4'h9 : add_81071[3:0]] + smul_81198;
  assign array_update_81201[0] = add_81071 == 32'h0000_0000 ? add_81200 : array_index_81194[0];
  assign array_update_81201[1] = add_81071 == 32'h0000_0001 ? add_81200 : array_index_81194[1];
  assign array_update_81201[2] = add_81071 == 32'h0000_0002 ? add_81200 : array_index_81194[2];
  assign array_update_81201[3] = add_81071 == 32'h0000_0003 ? add_81200 : array_index_81194[3];
  assign array_update_81201[4] = add_81071 == 32'h0000_0004 ? add_81200 : array_index_81194[4];
  assign array_update_81201[5] = add_81071 == 32'h0000_0005 ? add_81200 : array_index_81194[5];
  assign array_update_81201[6] = add_81071 == 32'h0000_0006 ? add_81200 : array_index_81194[6];
  assign array_update_81201[7] = add_81071 == 32'h0000_0007 ? add_81200 : array_index_81194[7];
  assign array_update_81201[8] = add_81071 == 32'h0000_0008 ? add_81200 : array_index_81194[8];
  assign array_update_81201[9] = add_81071 == 32'h0000_0009 ? add_81200 : array_index_81194[9];
  assign array_update_81202[0] = add_80123 == 32'h0000_0000 ? array_update_81201 : array_update_81191[0];
  assign array_update_81202[1] = add_80123 == 32'h0000_0001 ? array_update_81201 : array_update_81191[1];
  assign array_update_81202[2] = add_80123 == 32'h0000_0002 ? array_update_81201 : array_update_81191[2];
  assign array_update_81202[3] = add_80123 == 32'h0000_0003 ? array_update_81201 : array_update_81191[3];
  assign array_update_81202[4] = add_80123 == 32'h0000_0004 ? array_update_81201 : array_update_81191[4];
  assign array_update_81202[5] = add_80123 == 32'h0000_0005 ? array_update_81201 : array_update_81191[5];
  assign array_update_81202[6] = add_80123 == 32'h0000_0006 ? array_update_81201 : array_update_81191[6];
  assign array_update_81202[7] = add_80123 == 32'h0000_0007 ? array_update_81201 : array_update_81191[7];
  assign array_update_81202[8] = add_80123 == 32'h0000_0008 ? array_update_81201 : array_update_81191[8];
  assign array_update_81202[9] = add_80123 == 32'h0000_0009 ? array_update_81201 : array_update_81191[9];
  assign array_index_81204 = array_update_81202[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign add_81206 = add_81071 + 32'h0000_0001;
  assign array_update_81207[0] = add_81206 == 32'h0000_0000 ? 32'h0000_0000 : array_index_81204[0];
  assign array_update_81207[1] = add_81206 == 32'h0000_0001 ? 32'h0000_0000 : array_index_81204[1];
  assign array_update_81207[2] = add_81206 == 32'h0000_0002 ? 32'h0000_0000 : array_index_81204[2];
  assign array_update_81207[3] = add_81206 == 32'h0000_0003 ? 32'h0000_0000 : array_index_81204[3];
  assign array_update_81207[4] = add_81206 == 32'h0000_0004 ? 32'h0000_0000 : array_index_81204[4];
  assign array_update_81207[5] = add_81206 == 32'h0000_0005 ? 32'h0000_0000 : array_index_81204[5];
  assign array_update_81207[6] = add_81206 == 32'h0000_0006 ? 32'h0000_0000 : array_index_81204[6];
  assign array_update_81207[7] = add_81206 == 32'h0000_0007 ? 32'h0000_0000 : array_index_81204[7];
  assign array_update_81207[8] = add_81206 == 32'h0000_0008 ? 32'h0000_0000 : array_index_81204[8];
  assign array_update_81207[9] = add_81206 == 32'h0000_0009 ? 32'h0000_0000 : array_index_81204[9];
  assign literal_81208 = 32'h0000_0000;
  assign array_update_81209[0] = add_80123 == 32'h0000_0000 ? array_update_81207 : array_update_81202[0];
  assign array_update_81209[1] = add_80123 == 32'h0000_0001 ? array_update_81207 : array_update_81202[1];
  assign array_update_81209[2] = add_80123 == 32'h0000_0002 ? array_update_81207 : array_update_81202[2];
  assign array_update_81209[3] = add_80123 == 32'h0000_0003 ? array_update_81207 : array_update_81202[3];
  assign array_update_81209[4] = add_80123 == 32'h0000_0004 ? array_update_81207 : array_update_81202[4];
  assign array_update_81209[5] = add_80123 == 32'h0000_0005 ? array_update_81207 : array_update_81202[5];
  assign array_update_81209[6] = add_80123 == 32'h0000_0006 ? array_update_81207 : array_update_81202[6];
  assign array_update_81209[7] = add_80123 == 32'h0000_0007 ? array_update_81207 : array_update_81202[7];
  assign array_update_81209[8] = add_80123 == 32'h0000_0008 ? array_update_81207 : array_update_81202[8];
  assign array_update_81209[9] = add_80123 == 32'h0000_0009 ? array_update_81207 : array_update_81202[9];
  assign array_index_81211 = array_update_72021[literal_81208 > 32'h0000_0009 ? 4'h9 : literal_81208[3:0]];
  assign array_index_81212 = array_update_81209[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_81216 = smul32b_32b_x_32b(array_index_80130[literal_81208 > 32'h0000_0009 ? 4'h9 : literal_81208[3:0]], array_index_81211[add_81206 > 32'h0000_0009 ? 4'h9 : add_81206[3:0]]);
  assign add_81218 = array_index_81212[add_81206 > 32'h0000_0009 ? 4'h9 : add_81206[3:0]] + smul_81216;
  assign array_update_81220[0] = add_81206 == 32'h0000_0000 ? add_81218 : array_index_81212[0];
  assign array_update_81220[1] = add_81206 == 32'h0000_0001 ? add_81218 : array_index_81212[1];
  assign array_update_81220[2] = add_81206 == 32'h0000_0002 ? add_81218 : array_index_81212[2];
  assign array_update_81220[3] = add_81206 == 32'h0000_0003 ? add_81218 : array_index_81212[3];
  assign array_update_81220[4] = add_81206 == 32'h0000_0004 ? add_81218 : array_index_81212[4];
  assign array_update_81220[5] = add_81206 == 32'h0000_0005 ? add_81218 : array_index_81212[5];
  assign array_update_81220[6] = add_81206 == 32'h0000_0006 ? add_81218 : array_index_81212[6];
  assign array_update_81220[7] = add_81206 == 32'h0000_0007 ? add_81218 : array_index_81212[7];
  assign array_update_81220[8] = add_81206 == 32'h0000_0008 ? add_81218 : array_index_81212[8];
  assign array_update_81220[9] = add_81206 == 32'h0000_0009 ? add_81218 : array_index_81212[9];
  assign add_81221 = literal_81208 + 32'h0000_0001;
  assign array_update_81222[0] = add_80123 == 32'h0000_0000 ? array_update_81220 : array_update_81209[0];
  assign array_update_81222[1] = add_80123 == 32'h0000_0001 ? array_update_81220 : array_update_81209[1];
  assign array_update_81222[2] = add_80123 == 32'h0000_0002 ? array_update_81220 : array_update_81209[2];
  assign array_update_81222[3] = add_80123 == 32'h0000_0003 ? array_update_81220 : array_update_81209[3];
  assign array_update_81222[4] = add_80123 == 32'h0000_0004 ? array_update_81220 : array_update_81209[4];
  assign array_update_81222[5] = add_80123 == 32'h0000_0005 ? array_update_81220 : array_update_81209[5];
  assign array_update_81222[6] = add_80123 == 32'h0000_0006 ? array_update_81220 : array_update_81209[6];
  assign array_update_81222[7] = add_80123 == 32'h0000_0007 ? array_update_81220 : array_update_81209[7];
  assign array_update_81222[8] = add_80123 == 32'h0000_0008 ? array_update_81220 : array_update_81209[8];
  assign array_update_81222[9] = add_80123 == 32'h0000_0009 ? array_update_81220 : array_update_81209[9];
  assign array_index_81224 = array_update_72021[add_81221 > 32'h0000_0009 ? 4'h9 : add_81221[3:0]];
  assign array_index_81225 = array_update_81222[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_81229 = smul32b_32b_x_32b(array_index_80130[add_81221 > 32'h0000_0009 ? 4'h9 : add_81221[3:0]], array_index_81224[add_81206 > 32'h0000_0009 ? 4'h9 : add_81206[3:0]]);
  assign add_81231 = array_index_81225[add_81206 > 32'h0000_0009 ? 4'h9 : add_81206[3:0]] + smul_81229;
  assign array_update_81233[0] = add_81206 == 32'h0000_0000 ? add_81231 : array_index_81225[0];
  assign array_update_81233[1] = add_81206 == 32'h0000_0001 ? add_81231 : array_index_81225[1];
  assign array_update_81233[2] = add_81206 == 32'h0000_0002 ? add_81231 : array_index_81225[2];
  assign array_update_81233[3] = add_81206 == 32'h0000_0003 ? add_81231 : array_index_81225[3];
  assign array_update_81233[4] = add_81206 == 32'h0000_0004 ? add_81231 : array_index_81225[4];
  assign array_update_81233[5] = add_81206 == 32'h0000_0005 ? add_81231 : array_index_81225[5];
  assign array_update_81233[6] = add_81206 == 32'h0000_0006 ? add_81231 : array_index_81225[6];
  assign array_update_81233[7] = add_81206 == 32'h0000_0007 ? add_81231 : array_index_81225[7];
  assign array_update_81233[8] = add_81206 == 32'h0000_0008 ? add_81231 : array_index_81225[8];
  assign array_update_81233[9] = add_81206 == 32'h0000_0009 ? add_81231 : array_index_81225[9];
  assign add_81234 = add_81221 + 32'h0000_0001;
  assign array_update_81235[0] = add_80123 == 32'h0000_0000 ? array_update_81233 : array_update_81222[0];
  assign array_update_81235[1] = add_80123 == 32'h0000_0001 ? array_update_81233 : array_update_81222[1];
  assign array_update_81235[2] = add_80123 == 32'h0000_0002 ? array_update_81233 : array_update_81222[2];
  assign array_update_81235[3] = add_80123 == 32'h0000_0003 ? array_update_81233 : array_update_81222[3];
  assign array_update_81235[4] = add_80123 == 32'h0000_0004 ? array_update_81233 : array_update_81222[4];
  assign array_update_81235[5] = add_80123 == 32'h0000_0005 ? array_update_81233 : array_update_81222[5];
  assign array_update_81235[6] = add_80123 == 32'h0000_0006 ? array_update_81233 : array_update_81222[6];
  assign array_update_81235[7] = add_80123 == 32'h0000_0007 ? array_update_81233 : array_update_81222[7];
  assign array_update_81235[8] = add_80123 == 32'h0000_0008 ? array_update_81233 : array_update_81222[8];
  assign array_update_81235[9] = add_80123 == 32'h0000_0009 ? array_update_81233 : array_update_81222[9];
  assign array_index_81237 = array_update_72021[add_81234 > 32'h0000_0009 ? 4'h9 : add_81234[3:0]];
  assign array_index_81238 = array_update_81235[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_81242 = smul32b_32b_x_32b(array_index_80130[add_81234 > 32'h0000_0009 ? 4'h9 : add_81234[3:0]], array_index_81237[add_81206 > 32'h0000_0009 ? 4'h9 : add_81206[3:0]]);
  assign add_81244 = array_index_81238[add_81206 > 32'h0000_0009 ? 4'h9 : add_81206[3:0]] + smul_81242;
  assign array_update_81246[0] = add_81206 == 32'h0000_0000 ? add_81244 : array_index_81238[0];
  assign array_update_81246[1] = add_81206 == 32'h0000_0001 ? add_81244 : array_index_81238[1];
  assign array_update_81246[2] = add_81206 == 32'h0000_0002 ? add_81244 : array_index_81238[2];
  assign array_update_81246[3] = add_81206 == 32'h0000_0003 ? add_81244 : array_index_81238[3];
  assign array_update_81246[4] = add_81206 == 32'h0000_0004 ? add_81244 : array_index_81238[4];
  assign array_update_81246[5] = add_81206 == 32'h0000_0005 ? add_81244 : array_index_81238[5];
  assign array_update_81246[6] = add_81206 == 32'h0000_0006 ? add_81244 : array_index_81238[6];
  assign array_update_81246[7] = add_81206 == 32'h0000_0007 ? add_81244 : array_index_81238[7];
  assign array_update_81246[8] = add_81206 == 32'h0000_0008 ? add_81244 : array_index_81238[8];
  assign array_update_81246[9] = add_81206 == 32'h0000_0009 ? add_81244 : array_index_81238[9];
  assign add_81247 = add_81234 + 32'h0000_0001;
  assign array_update_81248[0] = add_80123 == 32'h0000_0000 ? array_update_81246 : array_update_81235[0];
  assign array_update_81248[1] = add_80123 == 32'h0000_0001 ? array_update_81246 : array_update_81235[1];
  assign array_update_81248[2] = add_80123 == 32'h0000_0002 ? array_update_81246 : array_update_81235[2];
  assign array_update_81248[3] = add_80123 == 32'h0000_0003 ? array_update_81246 : array_update_81235[3];
  assign array_update_81248[4] = add_80123 == 32'h0000_0004 ? array_update_81246 : array_update_81235[4];
  assign array_update_81248[5] = add_80123 == 32'h0000_0005 ? array_update_81246 : array_update_81235[5];
  assign array_update_81248[6] = add_80123 == 32'h0000_0006 ? array_update_81246 : array_update_81235[6];
  assign array_update_81248[7] = add_80123 == 32'h0000_0007 ? array_update_81246 : array_update_81235[7];
  assign array_update_81248[8] = add_80123 == 32'h0000_0008 ? array_update_81246 : array_update_81235[8];
  assign array_update_81248[9] = add_80123 == 32'h0000_0009 ? array_update_81246 : array_update_81235[9];
  assign array_index_81250 = array_update_72021[add_81247 > 32'h0000_0009 ? 4'h9 : add_81247[3:0]];
  assign array_index_81251 = array_update_81248[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_81255 = smul32b_32b_x_32b(array_index_80130[add_81247 > 32'h0000_0009 ? 4'h9 : add_81247[3:0]], array_index_81250[add_81206 > 32'h0000_0009 ? 4'h9 : add_81206[3:0]]);
  assign add_81257 = array_index_81251[add_81206 > 32'h0000_0009 ? 4'h9 : add_81206[3:0]] + smul_81255;
  assign array_update_81259[0] = add_81206 == 32'h0000_0000 ? add_81257 : array_index_81251[0];
  assign array_update_81259[1] = add_81206 == 32'h0000_0001 ? add_81257 : array_index_81251[1];
  assign array_update_81259[2] = add_81206 == 32'h0000_0002 ? add_81257 : array_index_81251[2];
  assign array_update_81259[3] = add_81206 == 32'h0000_0003 ? add_81257 : array_index_81251[3];
  assign array_update_81259[4] = add_81206 == 32'h0000_0004 ? add_81257 : array_index_81251[4];
  assign array_update_81259[5] = add_81206 == 32'h0000_0005 ? add_81257 : array_index_81251[5];
  assign array_update_81259[6] = add_81206 == 32'h0000_0006 ? add_81257 : array_index_81251[6];
  assign array_update_81259[7] = add_81206 == 32'h0000_0007 ? add_81257 : array_index_81251[7];
  assign array_update_81259[8] = add_81206 == 32'h0000_0008 ? add_81257 : array_index_81251[8];
  assign array_update_81259[9] = add_81206 == 32'h0000_0009 ? add_81257 : array_index_81251[9];
  assign add_81260 = add_81247 + 32'h0000_0001;
  assign array_update_81261[0] = add_80123 == 32'h0000_0000 ? array_update_81259 : array_update_81248[0];
  assign array_update_81261[1] = add_80123 == 32'h0000_0001 ? array_update_81259 : array_update_81248[1];
  assign array_update_81261[2] = add_80123 == 32'h0000_0002 ? array_update_81259 : array_update_81248[2];
  assign array_update_81261[3] = add_80123 == 32'h0000_0003 ? array_update_81259 : array_update_81248[3];
  assign array_update_81261[4] = add_80123 == 32'h0000_0004 ? array_update_81259 : array_update_81248[4];
  assign array_update_81261[5] = add_80123 == 32'h0000_0005 ? array_update_81259 : array_update_81248[5];
  assign array_update_81261[6] = add_80123 == 32'h0000_0006 ? array_update_81259 : array_update_81248[6];
  assign array_update_81261[7] = add_80123 == 32'h0000_0007 ? array_update_81259 : array_update_81248[7];
  assign array_update_81261[8] = add_80123 == 32'h0000_0008 ? array_update_81259 : array_update_81248[8];
  assign array_update_81261[9] = add_80123 == 32'h0000_0009 ? array_update_81259 : array_update_81248[9];
  assign array_index_81263 = array_update_72021[add_81260 > 32'h0000_0009 ? 4'h9 : add_81260[3:0]];
  assign array_index_81264 = array_update_81261[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_81268 = smul32b_32b_x_32b(array_index_80130[add_81260 > 32'h0000_0009 ? 4'h9 : add_81260[3:0]], array_index_81263[add_81206 > 32'h0000_0009 ? 4'h9 : add_81206[3:0]]);
  assign add_81270 = array_index_81264[add_81206 > 32'h0000_0009 ? 4'h9 : add_81206[3:0]] + smul_81268;
  assign array_update_81272[0] = add_81206 == 32'h0000_0000 ? add_81270 : array_index_81264[0];
  assign array_update_81272[1] = add_81206 == 32'h0000_0001 ? add_81270 : array_index_81264[1];
  assign array_update_81272[2] = add_81206 == 32'h0000_0002 ? add_81270 : array_index_81264[2];
  assign array_update_81272[3] = add_81206 == 32'h0000_0003 ? add_81270 : array_index_81264[3];
  assign array_update_81272[4] = add_81206 == 32'h0000_0004 ? add_81270 : array_index_81264[4];
  assign array_update_81272[5] = add_81206 == 32'h0000_0005 ? add_81270 : array_index_81264[5];
  assign array_update_81272[6] = add_81206 == 32'h0000_0006 ? add_81270 : array_index_81264[6];
  assign array_update_81272[7] = add_81206 == 32'h0000_0007 ? add_81270 : array_index_81264[7];
  assign array_update_81272[8] = add_81206 == 32'h0000_0008 ? add_81270 : array_index_81264[8];
  assign array_update_81272[9] = add_81206 == 32'h0000_0009 ? add_81270 : array_index_81264[9];
  assign add_81273 = add_81260 + 32'h0000_0001;
  assign array_update_81274[0] = add_80123 == 32'h0000_0000 ? array_update_81272 : array_update_81261[0];
  assign array_update_81274[1] = add_80123 == 32'h0000_0001 ? array_update_81272 : array_update_81261[1];
  assign array_update_81274[2] = add_80123 == 32'h0000_0002 ? array_update_81272 : array_update_81261[2];
  assign array_update_81274[3] = add_80123 == 32'h0000_0003 ? array_update_81272 : array_update_81261[3];
  assign array_update_81274[4] = add_80123 == 32'h0000_0004 ? array_update_81272 : array_update_81261[4];
  assign array_update_81274[5] = add_80123 == 32'h0000_0005 ? array_update_81272 : array_update_81261[5];
  assign array_update_81274[6] = add_80123 == 32'h0000_0006 ? array_update_81272 : array_update_81261[6];
  assign array_update_81274[7] = add_80123 == 32'h0000_0007 ? array_update_81272 : array_update_81261[7];
  assign array_update_81274[8] = add_80123 == 32'h0000_0008 ? array_update_81272 : array_update_81261[8];
  assign array_update_81274[9] = add_80123 == 32'h0000_0009 ? array_update_81272 : array_update_81261[9];
  assign array_index_81276 = array_update_72021[add_81273 > 32'h0000_0009 ? 4'h9 : add_81273[3:0]];
  assign array_index_81277 = array_update_81274[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_81281 = smul32b_32b_x_32b(array_index_80130[add_81273 > 32'h0000_0009 ? 4'h9 : add_81273[3:0]], array_index_81276[add_81206 > 32'h0000_0009 ? 4'h9 : add_81206[3:0]]);
  assign add_81283 = array_index_81277[add_81206 > 32'h0000_0009 ? 4'h9 : add_81206[3:0]] + smul_81281;
  assign array_update_81285[0] = add_81206 == 32'h0000_0000 ? add_81283 : array_index_81277[0];
  assign array_update_81285[1] = add_81206 == 32'h0000_0001 ? add_81283 : array_index_81277[1];
  assign array_update_81285[2] = add_81206 == 32'h0000_0002 ? add_81283 : array_index_81277[2];
  assign array_update_81285[3] = add_81206 == 32'h0000_0003 ? add_81283 : array_index_81277[3];
  assign array_update_81285[4] = add_81206 == 32'h0000_0004 ? add_81283 : array_index_81277[4];
  assign array_update_81285[5] = add_81206 == 32'h0000_0005 ? add_81283 : array_index_81277[5];
  assign array_update_81285[6] = add_81206 == 32'h0000_0006 ? add_81283 : array_index_81277[6];
  assign array_update_81285[7] = add_81206 == 32'h0000_0007 ? add_81283 : array_index_81277[7];
  assign array_update_81285[8] = add_81206 == 32'h0000_0008 ? add_81283 : array_index_81277[8];
  assign array_update_81285[9] = add_81206 == 32'h0000_0009 ? add_81283 : array_index_81277[9];
  assign add_81286 = add_81273 + 32'h0000_0001;
  assign array_update_81287[0] = add_80123 == 32'h0000_0000 ? array_update_81285 : array_update_81274[0];
  assign array_update_81287[1] = add_80123 == 32'h0000_0001 ? array_update_81285 : array_update_81274[1];
  assign array_update_81287[2] = add_80123 == 32'h0000_0002 ? array_update_81285 : array_update_81274[2];
  assign array_update_81287[3] = add_80123 == 32'h0000_0003 ? array_update_81285 : array_update_81274[3];
  assign array_update_81287[4] = add_80123 == 32'h0000_0004 ? array_update_81285 : array_update_81274[4];
  assign array_update_81287[5] = add_80123 == 32'h0000_0005 ? array_update_81285 : array_update_81274[5];
  assign array_update_81287[6] = add_80123 == 32'h0000_0006 ? array_update_81285 : array_update_81274[6];
  assign array_update_81287[7] = add_80123 == 32'h0000_0007 ? array_update_81285 : array_update_81274[7];
  assign array_update_81287[8] = add_80123 == 32'h0000_0008 ? array_update_81285 : array_update_81274[8];
  assign array_update_81287[9] = add_80123 == 32'h0000_0009 ? array_update_81285 : array_update_81274[9];
  assign array_index_81289 = array_update_72021[add_81286 > 32'h0000_0009 ? 4'h9 : add_81286[3:0]];
  assign array_index_81290 = array_update_81287[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_81294 = smul32b_32b_x_32b(array_index_80130[add_81286 > 32'h0000_0009 ? 4'h9 : add_81286[3:0]], array_index_81289[add_81206 > 32'h0000_0009 ? 4'h9 : add_81206[3:0]]);
  assign add_81296 = array_index_81290[add_81206 > 32'h0000_0009 ? 4'h9 : add_81206[3:0]] + smul_81294;
  assign array_update_81298[0] = add_81206 == 32'h0000_0000 ? add_81296 : array_index_81290[0];
  assign array_update_81298[1] = add_81206 == 32'h0000_0001 ? add_81296 : array_index_81290[1];
  assign array_update_81298[2] = add_81206 == 32'h0000_0002 ? add_81296 : array_index_81290[2];
  assign array_update_81298[3] = add_81206 == 32'h0000_0003 ? add_81296 : array_index_81290[3];
  assign array_update_81298[4] = add_81206 == 32'h0000_0004 ? add_81296 : array_index_81290[4];
  assign array_update_81298[5] = add_81206 == 32'h0000_0005 ? add_81296 : array_index_81290[5];
  assign array_update_81298[6] = add_81206 == 32'h0000_0006 ? add_81296 : array_index_81290[6];
  assign array_update_81298[7] = add_81206 == 32'h0000_0007 ? add_81296 : array_index_81290[7];
  assign array_update_81298[8] = add_81206 == 32'h0000_0008 ? add_81296 : array_index_81290[8];
  assign array_update_81298[9] = add_81206 == 32'h0000_0009 ? add_81296 : array_index_81290[9];
  assign add_81299 = add_81286 + 32'h0000_0001;
  assign array_update_81300[0] = add_80123 == 32'h0000_0000 ? array_update_81298 : array_update_81287[0];
  assign array_update_81300[1] = add_80123 == 32'h0000_0001 ? array_update_81298 : array_update_81287[1];
  assign array_update_81300[2] = add_80123 == 32'h0000_0002 ? array_update_81298 : array_update_81287[2];
  assign array_update_81300[3] = add_80123 == 32'h0000_0003 ? array_update_81298 : array_update_81287[3];
  assign array_update_81300[4] = add_80123 == 32'h0000_0004 ? array_update_81298 : array_update_81287[4];
  assign array_update_81300[5] = add_80123 == 32'h0000_0005 ? array_update_81298 : array_update_81287[5];
  assign array_update_81300[6] = add_80123 == 32'h0000_0006 ? array_update_81298 : array_update_81287[6];
  assign array_update_81300[7] = add_80123 == 32'h0000_0007 ? array_update_81298 : array_update_81287[7];
  assign array_update_81300[8] = add_80123 == 32'h0000_0008 ? array_update_81298 : array_update_81287[8];
  assign array_update_81300[9] = add_80123 == 32'h0000_0009 ? array_update_81298 : array_update_81287[9];
  assign array_index_81302 = array_update_72021[add_81299 > 32'h0000_0009 ? 4'h9 : add_81299[3:0]];
  assign array_index_81303 = array_update_81300[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_81307 = smul32b_32b_x_32b(array_index_80130[add_81299 > 32'h0000_0009 ? 4'h9 : add_81299[3:0]], array_index_81302[add_81206 > 32'h0000_0009 ? 4'h9 : add_81206[3:0]]);
  assign add_81309 = array_index_81303[add_81206 > 32'h0000_0009 ? 4'h9 : add_81206[3:0]] + smul_81307;
  assign array_update_81311[0] = add_81206 == 32'h0000_0000 ? add_81309 : array_index_81303[0];
  assign array_update_81311[1] = add_81206 == 32'h0000_0001 ? add_81309 : array_index_81303[1];
  assign array_update_81311[2] = add_81206 == 32'h0000_0002 ? add_81309 : array_index_81303[2];
  assign array_update_81311[3] = add_81206 == 32'h0000_0003 ? add_81309 : array_index_81303[3];
  assign array_update_81311[4] = add_81206 == 32'h0000_0004 ? add_81309 : array_index_81303[4];
  assign array_update_81311[5] = add_81206 == 32'h0000_0005 ? add_81309 : array_index_81303[5];
  assign array_update_81311[6] = add_81206 == 32'h0000_0006 ? add_81309 : array_index_81303[6];
  assign array_update_81311[7] = add_81206 == 32'h0000_0007 ? add_81309 : array_index_81303[7];
  assign array_update_81311[8] = add_81206 == 32'h0000_0008 ? add_81309 : array_index_81303[8];
  assign array_update_81311[9] = add_81206 == 32'h0000_0009 ? add_81309 : array_index_81303[9];
  assign add_81312 = add_81299 + 32'h0000_0001;
  assign array_update_81313[0] = add_80123 == 32'h0000_0000 ? array_update_81311 : array_update_81300[0];
  assign array_update_81313[1] = add_80123 == 32'h0000_0001 ? array_update_81311 : array_update_81300[1];
  assign array_update_81313[2] = add_80123 == 32'h0000_0002 ? array_update_81311 : array_update_81300[2];
  assign array_update_81313[3] = add_80123 == 32'h0000_0003 ? array_update_81311 : array_update_81300[3];
  assign array_update_81313[4] = add_80123 == 32'h0000_0004 ? array_update_81311 : array_update_81300[4];
  assign array_update_81313[5] = add_80123 == 32'h0000_0005 ? array_update_81311 : array_update_81300[5];
  assign array_update_81313[6] = add_80123 == 32'h0000_0006 ? array_update_81311 : array_update_81300[6];
  assign array_update_81313[7] = add_80123 == 32'h0000_0007 ? array_update_81311 : array_update_81300[7];
  assign array_update_81313[8] = add_80123 == 32'h0000_0008 ? array_update_81311 : array_update_81300[8];
  assign array_update_81313[9] = add_80123 == 32'h0000_0009 ? array_update_81311 : array_update_81300[9];
  assign array_index_81315 = array_update_72021[add_81312 > 32'h0000_0009 ? 4'h9 : add_81312[3:0]];
  assign array_index_81316 = array_update_81313[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_81320 = smul32b_32b_x_32b(array_index_80130[add_81312 > 32'h0000_0009 ? 4'h9 : add_81312[3:0]], array_index_81315[add_81206 > 32'h0000_0009 ? 4'h9 : add_81206[3:0]]);
  assign add_81322 = array_index_81316[add_81206 > 32'h0000_0009 ? 4'h9 : add_81206[3:0]] + smul_81320;
  assign array_update_81324[0] = add_81206 == 32'h0000_0000 ? add_81322 : array_index_81316[0];
  assign array_update_81324[1] = add_81206 == 32'h0000_0001 ? add_81322 : array_index_81316[1];
  assign array_update_81324[2] = add_81206 == 32'h0000_0002 ? add_81322 : array_index_81316[2];
  assign array_update_81324[3] = add_81206 == 32'h0000_0003 ? add_81322 : array_index_81316[3];
  assign array_update_81324[4] = add_81206 == 32'h0000_0004 ? add_81322 : array_index_81316[4];
  assign array_update_81324[5] = add_81206 == 32'h0000_0005 ? add_81322 : array_index_81316[5];
  assign array_update_81324[6] = add_81206 == 32'h0000_0006 ? add_81322 : array_index_81316[6];
  assign array_update_81324[7] = add_81206 == 32'h0000_0007 ? add_81322 : array_index_81316[7];
  assign array_update_81324[8] = add_81206 == 32'h0000_0008 ? add_81322 : array_index_81316[8];
  assign array_update_81324[9] = add_81206 == 32'h0000_0009 ? add_81322 : array_index_81316[9];
  assign add_81325 = add_81312 + 32'h0000_0001;
  assign array_update_81326[0] = add_80123 == 32'h0000_0000 ? array_update_81324 : array_update_81313[0];
  assign array_update_81326[1] = add_80123 == 32'h0000_0001 ? array_update_81324 : array_update_81313[1];
  assign array_update_81326[2] = add_80123 == 32'h0000_0002 ? array_update_81324 : array_update_81313[2];
  assign array_update_81326[3] = add_80123 == 32'h0000_0003 ? array_update_81324 : array_update_81313[3];
  assign array_update_81326[4] = add_80123 == 32'h0000_0004 ? array_update_81324 : array_update_81313[4];
  assign array_update_81326[5] = add_80123 == 32'h0000_0005 ? array_update_81324 : array_update_81313[5];
  assign array_update_81326[6] = add_80123 == 32'h0000_0006 ? array_update_81324 : array_update_81313[6];
  assign array_update_81326[7] = add_80123 == 32'h0000_0007 ? array_update_81324 : array_update_81313[7];
  assign array_update_81326[8] = add_80123 == 32'h0000_0008 ? array_update_81324 : array_update_81313[8];
  assign array_update_81326[9] = add_80123 == 32'h0000_0009 ? array_update_81324 : array_update_81313[9];
  assign array_index_81328 = array_update_72021[add_81325 > 32'h0000_0009 ? 4'h9 : add_81325[3:0]];
  assign array_index_81329 = array_update_81326[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_81333 = smul32b_32b_x_32b(array_index_80130[add_81325 > 32'h0000_0009 ? 4'h9 : add_81325[3:0]], array_index_81328[add_81206 > 32'h0000_0009 ? 4'h9 : add_81206[3:0]]);
  assign add_81335 = array_index_81329[add_81206 > 32'h0000_0009 ? 4'h9 : add_81206[3:0]] + smul_81333;
  assign array_update_81336[0] = add_81206 == 32'h0000_0000 ? add_81335 : array_index_81329[0];
  assign array_update_81336[1] = add_81206 == 32'h0000_0001 ? add_81335 : array_index_81329[1];
  assign array_update_81336[2] = add_81206 == 32'h0000_0002 ? add_81335 : array_index_81329[2];
  assign array_update_81336[3] = add_81206 == 32'h0000_0003 ? add_81335 : array_index_81329[3];
  assign array_update_81336[4] = add_81206 == 32'h0000_0004 ? add_81335 : array_index_81329[4];
  assign array_update_81336[5] = add_81206 == 32'h0000_0005 ? add_81335 : array_index_81329[5];
  assign array_update_81336[6] = add_81206 == 32'h0000_0006 ? add_81335 : array_index_81329[6];
  assign array_update_81336[7] = add_81206 == 32'h0000_0007 ? add_81335 : array_index_81329[7];
  assign array_update_81336[8] = add_81206 == 32'h0000_0008 ? add_81335 : array_index_81329[8];
  assign array_update_81336[9] = add_81206 == 32'h0000_0009 ? add_81335 : array_index_81329[9];
  assign array_update_81337[0] = add_80123 == 32'h0000_0000 ? array_update_81336 : array_update_81326[0];
  assign array_update_81337[1] = add_80123 == 32'h0000_0001 ? array_update_81336 : array_update_81326[1];
  assign array_update_81337[2] = add_80123 == 32'h0000_0002 ? array_update_81336 : array_update_81326[2];
  assign array_update_81337[3] = add_80123 == 32'h0000_0003 ? array_update_81336 : array_update_81326[3];
  assign array_update_81337[4] = add_80123 == 32'h0000_0004 ? array_update_81336 : array_update_81326[4];
  assign array_update_81337[5] = add_80123 == 32'h0000_0005 ? array_update_81336 : array_update_81326[5];
  assign array_update_81337[6] = add_80123 == 32'h0000_0006 ? array_update_81336 : array_update_81326[6];
  assign array_update_81337[7] = add_80123 == 32'h0000_0007 ? array_update_81336 : array_update_81326[7];
  assign array_update_81337[8] = add_80123 == 32'h0000_0008 ? array_update_81336 : array_update_81326[8];
  assign array_update_81337[9] = add_80123 == 32'h0000_0009 ? array_update_81336 : array_update_81326[9];
  assign array_index_81339 = array_update_81337[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign add_81341 = add_81206 + 32'h0000_0001;
  assign array_update_81342[0] = add_81341 == 32'h0000_0000 ? 32'h0000_0000 : array_index_81339[0];
  assign array_update_81342[1] = add_81341 == 32'h0000_0001 ? 32'h0000_0000 : array_index_81339[1];
  assign array_update_81342[2] = add_81341 == 32'h0000_0002 ? 32'h0000_0000 : array_index_81339[2];
  assign array_update_81342[3] = add_81341 == 32'h0000_0003 ? 32'h0000_0000 : array_index_81339[3];
  assign array_update_81342[4] = add_81341 == 32'h0000_0004 ? 32'h0000_0000 : array_index_81339[4];
  assign array_update_81342[5] = add_81341 == 32'h0000_0005 ? 32'h0000_0000 : array_index_81339[5];
  assign array_update_81342[6] = add_81341 == 32'h0000_0006 ? 32'h0000_0000 : array_index_81339[6];
  assign array_update_81342[7] = add_81341 == 32'h0000_0007 ? 32'h0000_0000 : array_index_81339[7];
  assign array_update_81342[8] = add_81341 == 32'h0000_0008 ? 32'h0000_0000 : array_index_81339[8];
  assign array_update_81342[9] = add_81341 == 32'h0000_0009 ? 32'h0000_0000 : array_index_81339[9];
  assign literal_81343 = 32'h0000_0000;
  assign array_update_81344[0] = add_80123 == 32'h0000_0000 ? array_update_81342 : array_update_81337[0];
  assign array_update_81344[1] = add_80123 == 32'h0000_0001 ? array_update_81342 : array_update_81337[1];
  assign array_update_81344[2] = add_80123 == 32'h0000_0002 ? array_update_81342 : array_update_81337[2];
  assign array_update_81344[3] = add_80123 == 32'h0000_0003 ? array_update_81342 : array_update_81337[3];
  assign array_update_81344[4] = add_80123 == 32'h0000_0004 ? array_update_81342 : array_update_81337[4];
  assign array_update_81344[5] = add_80123 == 32'h0000_0005 ? array_update_81342 : array_update_81337[5];
  assign array_update_81344[6] = add_80123 == 32'h0000_0006 ? array_update_81342 : array_update_81337[6];
  assign array_update_81344[7] = add_80123 == 32'h0000_0007 ? array_update_81342 : array_update_81337[7];
  assign array_update_81344[8] = add_80123 == 32'h0000_0008 ? array_update_81342 : array_update_81337[8];
  assign array_update_81344[9] = add_80123 == 32'h0000_0009 ? array_update_81342 : array_update_81337[9];
  assign array_index_81346 = array_update_72021[literal_81343 > 32'h0000_0009 ? 4'h9 : literal_81343[3:0]];
  assign array_index_81347 = array_update_81344[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_81351 = smul32b_32b_x_32b(array_index_80130[literal_81343 > 32'h0000_0009 ? 4'h9 : literal_81343[3:0]], array_index_81346[add_81341 > 32'h0000_0009 ? 4'h9 : add_81341[3:0]]);
  assign add_81353 = array_index_81347[add_81341 > 32'h0000_0009 ? 4'h9 : add_81341[3:0]] + smul_81351;
  assign array_update_81355[0] = add_81341 == 32'h0000_0000 ? add_81353 : array_index_81347[0];
  assign array_update_81355[1] = add_81341 == 32'h0000_0001 ? add_81353 : array_index_81347[1];
  assign array_update_81355[2] = add_81341 == 32'h0000_0002 ? add_81353 : array_index_81347[2];
  assign array_update_81355[3] = add_81341 == 32'h0000_0003 ? add_81353 : array_index_81347[3];
  assign array_update_81355[4] = add_81341 == 32'h0000_0004 ? add_81353 : array_index_81347[4];
  assign array_update_81355[5] = add_81341 == 32'h0000_0005 ? add_81353 : array_index_81347[5];
  assign array_update_81355[6] = add_81341 == 32'h0000_0006 ? add_81353 : array_index_81347[6];
  assign array_update_81355[7] = add_81341 == 32'h0000_0007 ? add_81353 : array_index_81347[7];
  assign array_update_81355[8] = add_81341 == 32'h0000_0008 ? add_81353 : array_index_81347[8];
  assign array_update_81355[9] = add_81341 == 32'h0000_0009 ? add_81353 : array_index_81347[9];
  assign add_81356 = literal_81343 + 32'h0000_0001;
  assign array_update_81357[0] = add_80123 == 32'h0000_0000 ? array_update_81355 : array_update_81344[0];
  assign array_update_81357[1] = add_80123 == 32'h0000_0001 ? array_update_81355 : array_update_81344[1];
  assign array_update_81357[2] = add_80123 == 32'h0000_0002 ? array_update_81355 : array_update_81344[2];
  assign array_update_81357[3] = add_80123 == 32'h0000_0003 ? array_update_81355 : array_update_81344[3];
  assign array_update_81357[4] = add_80123 == 32'h0000_0004 ? array_update_81355 : array_update_81344[4];
  assign array_update_81357[5] = add_80123 == 32'h0000_0005 ? array_update_81355 : array_update_81344[5];
  assign array_update_81357[6] = add_80123 == 32'h0000_0006 ? array_update_81355 : array_update_81344[6];
  assign array_update_81357[7] = add_80123 == 32'h0000_0007 ? array_update_81355 : array_update_81344[7];
  assign array_update_81357[8] = add_80123 == 32'h0000_0008 ? array_update_81355 : array_update_81344[8];
  assign array_update_81357[9] = add_80123 == 32'h0000_0009 ? array_update_81355 : array_update_81344[9];
  assign array_index_81359 = array_update_72021[add_81356 > 32'h0000_0009 ? 4'h9 : add_81356[3:0]];
  assign array_index_81360 = array_update_81357[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_81364 = smul32b_32b_x_32b(array_index_80130[add_81356 > 32'h0000_0009 ? 4'h9 : add_81356[3:0]], array_index_81359[add_81341 > 32'h0000_0009 ? 4'h9 : add_81341[3:0]]);
  assign add_81366 = array_index_81360[add_81341 > 32'h0000_0009 ? 4'h9 : add_81341[3:0]] + smul_81364;
  assign array_update_81368[0] = add_81341 == 32'h0000_0000 ? add_81366 : array_index_81360[0];
  assign array_update_81368[1] = add_81341 == 32'h0000_0001 ? add_81366 : array_index_81360[1];
  assign array_update_81368[2] = add_81341 == 32'h0000_0002 ? add_81366 : array_index_81360[2];
  assign array_update_81368[3] = add_81341 == 32'h0000_0003 ? add_81366 : array_index_81360[3];
  assign array_update_81368[4] = add_81341 == 32'h0000_0004 ? add_81366 : array_index_81360[4];
  assign array_update_81368[5] = add_81341 == 32'h0000_0005 ? add_81366 : array_index_81360[5];
  assign array_update_81368[6] = add_81341 == 32'h0000_0006 ? add_81366 : array_index_81360[6];
  assign array_update_81368[7] = add_81341 == 32'h0000_0007 ? add_81366 : array_index_81360[7];
  assign array_update_81368[8] = add_81341 == 32'h0000_0008 ? add_81366 : array_index_81360[8];
  assign array_update_81368[9] = add_81341 == 32'h0000_0009 ? add_81366 : array_index_81360[9];
  assign add_81369 = add_81356 + 32'h0000_0001;
  assign array_update_81370[0] = add_80123 == 32'h0000_0000 ? array_update_81368 : array_update_81357[0];
  assign array_update_81370[1] = add_80123 == 32'h0000_0001 ? array_update_81368 : array_update_81357[1];
  assign array_update_81370[2] = add_80123 == 32'h0000_0002 ? array_update_81368 : array_update_81357[2];
  assign array_update_81370[3] = add_80123 == 32'h0000_0003 ? array_update_81368 : array_update_81357[3];
  assign array_update_81370[4] = add_80123 == 32'h0000_0004 ? array_update_81368 : array_update_81357[4];
  assign array_update_81370[5] = add_80123 == 32'h0000_0005 ? array_update_81368 : array_update_81357[5];
  assign array_update_81370[6] = add_80123 == 32'h0000_0006 ? array_update_81368 : array_update_81357[6];
  assign array_update_81370[7] = add_80123 == 32'h0000_0007 ? array_update_81368 : array_update_81357[7];
  assign array_update_81370[8] = add_80123 == 32'h0000_0008 ? array_update_81368 : array_update_81357[8];
  assign array_update_81370[9] = add_80123 == 32'h0000_0009 ? array_update_81368 : array_update_81357[9];
  assign array_index_81372 = array_update_72021[add_81369 > 32'h0000_0009 ? 4'h9 : add_81369[3:0]];
  assign array_index_81373 = array_update_81370[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_81377 = smul32b_32b_x_32b(array_index_80130[add_81369 > 32'h0000_0009 ? 4'h9 : add_81369[3:0]], array_index_81372[add_81341 > 32'h0000_0009 ? 4'h9 : add_81341[3:0]]);
  assign add_81379 = array_index_81373[add_81341 > 32'h0000_0009 ? 4'h9 : add_81341[3:0]] + smul_81377;
  assign array_update_81381[0] = add_81341 == 32'h0000_0000 ? add_81379 : array_index_81373[0];
  assign array_update_81381[1] = add_81341 == 32'h0000_0001 ? add_81379 : array_index_81373[1];
  assign array_update_81381[2] = add_81341 == 32'h0000_0002 ? add_81379 : array_index_81373[2];
  assign array_update_81381[3] = add_81341 == 32'h0000_0003 ? add_81379 : array_index_81373[3];
  assign array_update_81381[4] = add_81341 == 32'h0000_0004 ? add_81379 : array_index_81373[4];
  assign array_update_81381[5] = add_81341 == 32'h0000_0005 ? add_81379 : array_index_81373[5];
  assign array_update_81381[6] = add_81341 == 32'h0000_0006 ? add_81379 : array_index_81373[6];
  assign array_update_81381[7] = add_81341 == 32'h0000_0007 ? add_81379 : array_index_81373[7];
  assign array_update_81381[8] = add_81341 == 32'h0000_0008 ? add_81379 : array_index_81373[8];
  assign array_update_81381[9] = add_81341 == 32'h0000_0009 ? add_81379 : array_index_81373[9];
  assign add_81382 = add_81369 + 32'h0000_0001;
  assign array_update_81383[0] = add_80123 == 32'h0000_0000 ? array_update_81381 : array_update_81370[0];
  assign array_update_81383[1] = add_80123 == 32'h0000_0001 ? array_update_81381 : array_update_81370[1];
  assign array_update_81383[2] = add_80123 == 32'h0000_0002 ? array_update_81381 : array_update_81370[2];
  assign array_update_81383[3] = add_80123 == 32'h0000_0003 ? array_update_81381 : array_update_81370[3];
  assign array_update_81383[4] = add_80123 == 32'h0000_0004 ? array_update_81381 : array_update_81370[4];
  assign array_update_81383[5] = add_80123 == 32'h0000_0005 ? array_update_81381 : array_update_81370[5];
  assign array_update_81383[6] = add_80123 == 32'h0000_0006 ? array_update_81381 : array_update_81370[6];
  assign array_update_81383[7] = add_80123 == 32'h0000_0007 ? array_update_81381 : array_update_81370[7];
  assign array_update_81383[8] = add_80123 == 32'h0000_0008 ? array_update_81381 : array_update_81370[8];
  assign array_update_81383[9] = add_80123 == 32'h0000_0009 ? array_update_81381 : array_update_81370[9];
  assign array_index_81385 = array_update_72021[add_81382 > 32'h0000_0009 ? 4'h9 : add_81382[3:0]];
  assign array_index_81386 = array_update_81383[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_81390 = smul32b_32b_x_32b(array_index_80130[add_81382 > 32'h0000_0009 ? 4'h9 : add_81382[3:0]], array_index_81385[add_81341 > 32'h0000_0009 ? 4'h9 : add_81341[3:0]]);
  assign add_81392 = array_index_81386[add_81341 > 32'h0000_0009 ? 4'h9 : add_81341[3:0]] + smul_81390;
  assign array_update_81394[0] = add_81341 == 32'h0000_0000 ? add_81392 : array_index_81386[0];
  assign array_update_81394[1] = add_81341 == 32'h0000_0001 ? add_81392 : array_index_81386[1];
  assign array_update_81394[2] = add_81341 == 32'h0000_0002 ? add_81392 : array_index_81386[2];
  assign array_update_81394[3] = add_81341 == 32'h0000_0003 ? add_81392 : array_index_81386[3];
  assign array_update_81394[4] = add_81341 == 32'h0000_0004 ? add_81392 : array_index_81386[4];
  assign array_update_81394[5] = add_81341 == 32'h0000_0005 ? add_81392 : array_index_81386[5];
  assign array_update_81394[6] = add_81341 == 32'h0000_0006 ? add_81392 : array_index_81386[6];
  assign array_update_81394[7] = add_81341 == 32'h0000_0007 ? add_81392 : array_index_81386[7];
  assign array_update_81394[8] = add_81341 == 32'h0000_0008 ? add_81392 : array_index_81386[8];
  assign array_update_81394[9] = add_81341 == 32'h0000_0009 ? add_81392 : array_index_81386[9];
  assign add_81395 = add_81382 + 32'h0000_0001;
  assign array_update_81396[0] = add_80123 == 32'h0000_0000 ? array_update_81394 : array_update_81383[0];
  assign array_update_81396[1] = add_80123 == 32'h0000_0001 ? array_update_81394 : array_update_81383[1];
  assign array_update_81396[2] = add_80123 == 32'h0000_0002 ? array_update_81394 : array_update_81383[2];
  assign array_update_81396[3] = add_80123 == 32'h0000_0003 ? array_update_81394 : array_update_81383[3];
  assign array_update_81396[4] = add_80123 == 32'h0000_0004 ? array_update_81394 : array_update_81383[4];
  assign array_update_81396[5] = add_80123 == 32'h0000_0005 ? array_update_81394 : array_update_81383[5];
  assign array_update_81396[6] = add_80123 == 32'h0000_0006 ? array_update_81394 : array_update_81383[6];
  assign array_update_81396[7] = add_80123 == 32'h0000_0007 ? array_update_81394 : array_update_81383[7];
  assign array_update_81396[8] = add_80123 == 32'h0000_0008 ? array_update_81394 : array_update_81383[8];
  assign array_update_81396[9] = add_80123 == 32'h0000_0009 ? array_update_81394 : array_update_81383[9];
  assign array_index_81398 = array_update_72021[add_81395 > 32'h0000_0009 ? 4'h9 : add_81395[3:0]];
  assign array_index_81399 = array_update_81396[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_81403 = smul32b_32b_x_32b(array_index_80130[add_81395 > 32'h0000_0009 ? 4'h9 : add_81395[3:0]], array_index_81398[add_81341 > 32'h0000_0009 ? 4'h9 : add_81341[3:0]]);
  assign add_81405 = array_index_81399[add_81341 > 32'h0000_0009 ? 4'h9 : add_81341[3:0]] + smul_81403;
  assign array_update_81407[0] = add_81341 == 32'h0000_0000 ? add_81405 : array_index_81399[0];
  assign array_update_81407[1] = add_81341 == 32'h0000_0001 ? add_81405 : array_index_81399[1];
  assign array_update_81407[2] = add_81341 == 32'h0000_0002 ? add_81405 : array_index_81399[2];
  assign array_update_81407[3] = add_81341 == 32'h0000_0003 ? add_81405 : array_index_81399[3];
  assign array_update_81407[4] = add_81341 == 32'h0000_0004 ? add_81405 : array_index_81399[4];
  assign array_update_81407[5] = add_81341 == 32'h0000_0005 ? add_81405 : array_index_81399[5];
  assign array_update_81407[6] = add_81341 == 32'h0000_0006 ? add_81405 : array_index_81399[6];
  assign array_update_81407[7] = add_81341 == 32'h0000_0007 ? add_81405 : array_index_81399[7];
  assign array_update_81407[8] = add_81341 == 32'h0000_0008 ? add_81405 : array_index_81399[8];
  assign array_update_81407[9] = add_81341 == 32'h0000_0009 ? add_81405 : array_index_81399[9];
  assign add_81408 = add_81395 + 32'h0000_0001;
  assign array_update_81409[0] = add_80123 == 32'h0000_0000 ? array_update_81407 : array_update_81396[0];
  assign array_update_81409[1] = add_80123 == 32'h0000_0001 ? array_update_81407 : array_update_81396[1];
  assign array_update_81409[2] = add_80123 == 32'h0000_0002 ? array_update_81407 : array_update_81396[2];
  assign array_update_81409[3] = add_80123 == 32'h0000_0003 ? array_update_81407 : array_update_81396[3];
  assign array_update_81409[4] = add_80123 == 32'h0000_0004 ? array_update_81407 : array_update_81396[4];
  assign array_update_81409[5] = add_80123 == 32'h0000_0005 ? array_update_81407 : array_update_81396[5];
  assign array_update_81409[6] = add_80123 == 32'h0000_0006 ? array_update_81407 : array_update_81396[6];
  assign array_update_81409[7] = add_80123 == 32'h0000_0007 ? array_update_81407 : array_update_81396[7];
  assign array_update_81409[8] = add_80123 == 32'h0000_0008 ? array_update_81407 : array_update_81396[8];
  assign array_update_81409[9] = add_80123 == 32'h0000_0009 ? array_update_81407 : array_update_81396[9];
  assign array_index_81411 = array_update_72021[add_81408 > 32'h0000_0009 ? 4'h9 : add_81408[3:0]];
  assign array_index_81412 = array_update_81409[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_81416 = smul32b_32b_x_32b(array_index_80130[add_81408 > 32'h0000_0009 ? 4'h9 : add_81408[3:0]], array_index_81411[add_81341 > 32'h0000_0009 ? 4'h9 : add_81341[3:0]]);
  assign add_81418 = array_index_81412[add_81341 > 32'h0000_0009 ? 4'h9 : add_81341[3:0]] + smul_81416;
  assign array_update_81420[0] = add_81341 == 32'h0000_0000 ? add_81418 : array_index_81412[0];
  assign array_update_81420[1] = add_81341 == 32'h0000_0001 ? add_81418 : array_index_81412[1];
  assign array_update_81420[2] = add_81341 == 32'h0000_0002 ? add_81418 : array_index_81412[2];
  assign array_update_81420[3] = add_81341 == 32'h0000_0003 ? add_81418 : array_index_81412[3];
  assign array_update_81420[4] = add_81341 == 32'h0000_0004 ? add_81418 : array_index_81412[4];
  assign array_update_81420[5] = add_81341 == 32'h0000_0005 ? add_81418 : array_index_81412[5];
  assign array_update_81420[6] = add_81341 == 32'h0000_0006 ? add_81418 : array_index_81412[6];
  assign array_update_81420[7] = add_81341 == 32'h0000_0007 ? add_81418 : array_index_81412[7];
  assign array_update_81420[8] = add_81341 == 32'h0000_0008 ? add_81418 : array_index_81412[8];
  assign array_update_81420[9] = add_81341 == 32'h0000_0009 ? add_81418 : array_index_81412[9];
  assign add_81421 = add_81408 + 32'h0000_0001;
  assign array_update_81422[0] = add_80123 == 32'h0000_0000 ? array_update_81420 : array_update_81409[0];
  assign array_update_81422[1] = add_80123 == 32'h0000_0001 ? array_update_81420 : array_update_81409[1];
  assign array_update_81422[2] = add_80123 == 32'h0000_0002 ? array_update_81420 : array_update_81409[2];
  assign array_update_81422[3] = add_80123 == 32'h0000_0003 ? array_update_81420 : array_update_81409[3];
  assign array_update_81422[4] = add_80123 == 32'h0000_0004 ? array_update_81420 : array_update_81409[4];
  assign array_update_81422[5] = add_80123 == 32'h0000_0005 ? array_update_81420 : array_update_81409[5];
  assign array_update_81422[6] = add_80123 == 32'h0000_0006 ? array_update_81420 : array_update_81409[6];
  assign array_update_81422[7] = add_80123 == 32'h0000_0007 ? array_update_81420 : array_update_81409[7];
  assign array_update_81422[8] = add_80123 == 32'h0000_0008 ? array_update_81420 : array_update_81409[8];
  assign array_update_81422[9] = add_80123 == 32'h0000_0009 ? array_update_81420 : array_update_81409[9];
  assign array_index_81424 = array_update_72021[add_81421 > 32'h0000_0009 ? 4'h9 : add_81421[3:0]];
  assign array_index_81425 = array_update_81422[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_81429 = smul32b_32b_x_32b(array_index_80130[add_81421 > 32'h0000_0009 ? 4'h9 : add_81421[3:0]], array_index_81424[add_81341 > 32'h0000_0009 ? 4'h9 : add_81341[3:0]]);
  assign add_81431 = array_index_81425[add_81341 > 32'h0000_0009 ? 4'h9 : add_81341[3:0]] + smul_81429;
  assign array_update_81433[0] = add_81341 == 32'h0000_0000 ? add_81431 : array_index_81425[0];
  assign array_update_81433[1] = add_81341 == 32'h0000_0001 ? add_81431 : array_index_81425[1];
  assign array_update_81433[2] = add_81341 == 32'h0000_0002 ? add_81431 : array_index_81425[2];
  assign array_update_81433[3] = add_81341 == 32'h0000_0003 ? add_81431 : array_index_81425[3];
  assign array_update_81433[4] = add_81341 == 32'h0000_0004 ? add_81431 : array_index_81425[4];
  assign array_update_81433[5] = add_81341 == 32'h0000_0005 ? add_81431 : array_index_81425[5];
  assign array_update_81433[6] = add_81341 == 32'h0000_0006 ? add_81431 : array_index_81425[6];
  assign array_update_81433[7] = add_81341 == 32'h0000_0007 ? add_81431 : array_index_81425[7];
  assign array_update_81433[8] = add_81341 == 32'h0000_0008 ? add_81431 : array_index_81425[8];
  assign array_update_81433[9] = add_81341 == 32'h0000_0009 ? add_81431 : array_index_81425[9];
  assign add_81434 = add_81421 + 32'h0000_0001;
  assign array_update_81435[0] = add_80123 == 32'h0000_0000 ? array_update_81433 : array_update_81422[0];
  assign array_update_81435[1] = add_80123 == 32'h0000_0001 ? array_update_81433 : array_update_81422[1];
  assign array_update_81435[2] = add_80123 == 32'h0000_0002 ? array_update_81433 : array_update_81422[2];
  assign array_update_81435[3] = add_80123 == 32'h0000_0003 ? array_update_81433 : array_update_81422[3];
  assign array_update_81435[4] = add_80123 == 32'h0000_0004 ? array_update_81433 : array_update_81422[4];
  assign array_update_81435[5] = add_80123 == 32'h0000_0005 ? array_update_81433 : array_update_81422[5];
  assign array_update_81435[6] = add_80123 == 32'h0000_0006 ? array_update_81433 : array_update_81422[6];
  assign array_update_81435[7] = add_80123 == 32'h0000_0007 ? array_update_81433 : array_update_81422[7];
  assign array_update_81435[8] = add_80123 == 32'h0000_0008 ? array_update_81433 : array_update_81422[8];
  assign array_update_81435[9] = add_80123 == 32'h0000_0009 ? array_update_81433 : array_update_81422[9];
  assign array_index_81437 = array_update_72021[add_81434 > 32'h0000_0009 ? 4'h9 : add_81434[3:0]];
  assign array_index_81438 = array_update_81435[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_81442 = smul32b_32b_x_32b(array_index_80130[add_81434 > 32'h0000_0009 ? 4'h9 : add_81434[3:0]], array_index_81437[add_81341 > 32'h0000_0009 ? 4'h9 : add_81341[3:0]]);
  assign add_81444 = array_index_81438[add_81341 > 32'h0000_0009 ? 4'h9 : add_81341[3:0]] + smul_81442;
  assign array_update_81446[0] = add_81341 == 32'h0000_0000 ? add_81444 : array_index_81438[0];
  assign array_update_81446[1] = add_81341 == 32'h0000_0001 ? add_81444 : array_index_81438[1];
  assign array_update_81446[2] = add_81341 == 32'h0000_0002 ? add_81444 : array_index_81438[2];
  assign array_update_81446[3] = add_81341 == 32'h0000_0003 ? add_81444 : array_index_81438[3];
  assign array_update_81446[4] = add_81341 == 32'h0000_0004 ? add_81444 : array_index_81438[4];
  assign array_update_81446[5] = add_81341 == 32'h0000_0005 ? add_81444 : array_index_81438[5];
  assign array_update_81446[6] = add_81341 == 32'h0000_0006 ? add_81444 : array_index_81438[6];
  assign array_update_81446[7] = add_81341 == 32'h0000_0007 ? add_81444 : array_index_81438[7];
  assign array_update_81446[8] = add_81341 == 32'h0000_0008 ? add_81444 : array_index_81438[8];
  assign array_update_81446[9] = add_81341 == 32'h0000_0009 ? add_81444 : array_index_81438[9];
  assign add_81447 = add_81434 + 32'h0000_0001;
  assign array_update_81448[0] = add_80123 == 32'h0000_0000 ? array_update_81446 : array_update_81435[0];
  assign array_update_81448[1] = add_80123 == 32'h0000_0001 ? array_update_81446 : array_update_81435[1];
  assign array_update_81448[2] = add_80123 == 32'h0000_0002 ? array_update_81446 : array_update_81435[2];
  assign array_update_81448[3] = add_80123 == 32'h0000_0003 ? array_update_81446 : array_update_81435[3];
  assign array_update_81448[4] = add_80123 == 32'h0000_0004 ? array_update_81446 : array_update_81435[4];
  assign array_update_81448[5] = add_80123 == 32'h0000_0005 ? array_update_81446 : array_update_81435[5];
  assign array_update_81448[6] = add_80123 == 32'h0000_0006 ? array_update_81446 : array_update_81435[6];
  assign array_update_81448[7] = add_80123 == 32'h0000_0007 ? array_update_81446 : array_update_81435[7];
  assign array_update_81448[8] = add_80123 == 32'h0000_0008 ? array_update_81446 : array_update_81435[8];
  assign array_update_81448[9] = add_80123 == 32'h0000_0009 ? array_update_81446 : array_update_81435[9];
  assign array_index_81450 = array_update_72021[add_81447 > 32'h0000_0009 ? 4'h9 : add_81447[3:0]];
  assign array_index_81451 = array_update_81448[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_81455 = smul32b_32b_x_32b(array_index_80130[add_81447 > 32'h0000_0009 ? 4'h9 : add_81447[3:0]], array_index_81450[add_81341 > 32'h0000_0009 ? 4'h9 : add_81341[3:0]]);
  assign add_81457 = array_index_81451[add_81341 > 32'h0000_0009 ? 4'h9 : add_81341[3:0]] + smul_81455;
  assign array_update_81459[0] = add_81341 == 32'h0000_0000 ? add_81457 : array_index_81451[0];
  assign array_update_81459[1] = add_81341 == 32'h0000_0001 ? add_81457 : array_index_81451[1];
  assign array_update_81459[2] = add_81341 == 32'h0000_0002 ? add_81457 : array_index_81451[2];
  assign array_update_81459[3] = add_81341 == 32'h0000_0003 ? add_81457 : array_index_81451[3];
  assign array_update_81459[4] = add_81341 == 32'h0000_0004 ? add_81457 : array_index_81451[4];
  assign array_update_81459[5] = add_81341 == 32'h0000_0005 ? add_81457 : array_index_81451[5];
  assign array_update_81459[6] = add_81341 == 32'h0000_0006 ? add_81457 : array_index_81451[6];
  assign array_update_81459[7] = add_81341 == 32'h0000_0007 ? add_81457 : array_index_81451[7];
  assign array_update_81459[8] = add_81341 == 32'h0000_0008 ? add_81457 : array_index_81451[8];
  assign array_update_81459[9] = add_81341 == 32'h0000_0009 ? add_81457 : array_index_81451[9];
  assign add_81460 = add_81447 + 32'h0000_0001;
  assign array_update_81461[0] = add_80123 == 32'h0000_0000 ? array_update_81459 : array_update_81448[0];
  assign array_update_81461[1] = add_80123 == 32'h0000_0001 ? array_update_81459 : array_update_81448[1];
  assign array_update_81461[2] = add_80123 == 32'h0000_0002 ? array_update_81459 : array_update_81448[2];
  assign array_update_81461[3] = add_80123 == 32'h0000_0003 ? array_update_81459 : array_update_81448[3];
  assign array_update_81461[4] = add_80123 == 32'h0000_0004 ? array_update_81459 : array_update_81448[4];
  assign array_update_81461[5] = add_80123 == 32'h0000_0005 ? array_update_81459 : array_update_81448[5];
  assign array_update_81461[6] = add_80123 == 32'h0000_0006 ? array_update_81459 : array_update_81448[6];
  assign array_update_81461[7] = add_80123 == 32'h0000_0007 ? array_update_81459 : array_update_81448[7];
  assign array_update_81461[8] = add_80123 == 32'h0000_0008 ? array_update_81459 : array_update_81448[8];
  assign array_update_81461[9] = add_80123 == 32'h0000_0009 ? array_update_81459 : array_update_81448[9];
  assign array_index_81463 = array_update_72021[add_81460 > 32'h0000_0009 ? 4'h9 : add_81460[3:0]];
  assign array_index_81464 = array_update_81461[add_80123 > 32'h0000_0009 ? 4'h9 : add_80123[3:0]];
  assign smul_81468 = smul32b_32b_x_32b(array_index_80130[add_81460 > 32'h0000_0009 ? 4'h9 : add_81460[3:0]], array_index_81463[add_81341 > 32'h0000_0009 ? 4'h9 : add_81341[3:0]]);
  assign add_81470 = array_index_81464[add_81341 > 32'h0000_0009 ? 4'h9 : add_81341[3:0]] + smul_81468;
  assign array_update_81471[0] = add_81341 == 32'h0000_0000 ? add_81470 : array_index_81464[0];
  assign array_update_81471[1] = add_81341 == 32'h0000_0001 ? add_81470 : array_index_81464[1];
  assign array_update_81471[2] = add_81341 == 32'h0000_0002 ? add_81470 : array_index_81464[2];
  assign array_update_81471[3] = add_81341 == 32'h0000_0003 ? add_81470 : array_index_81464[3];
  assign array_update_81471[4] = add_81341 == 32'h0000_0004 ? add_81470 : array_index_81464[4];
  assign array_update_81471[5] = add_81341 == 32'h0000_0005 ? add_81470 : array_index_81464[5];
  assign array_update_81471[6] = add_81341 == 32'h0000_0006 ? add_81470 : array_index_81464[6];
  assign array_update_81471[7] = add_81341 == 32'h0000_0007 ? add_81470 : array_index_81464[7];
  assign array_update_81471[8] = add_81341 == 32'h0000_0008 ? add_81470 : array_index_81464[8];
  assign array_update_81471[9] = add_81341 == 32'h0000_0009 ? add_81470 : array_index_81464[9];
  assign array_update_81473[0] = add_80123 == 32'h0000_0000 ? array_update_81471 : array_update_81461[0];
  assign array_update_81473[1] = add_80123 == 32'h0000_0001 ? array_update_81471 : array_update_81461[1];
  assign array_update_81473[2] = add_80123 == 32'h0000_0002 ? array_update_81471 : array_update_81461[2];
  assign array_update_81473[3] = add_80123 == 32'h0000_0003 ? array_update_81471 : array_update_81461[3];
  assign array_update_81473[4] = add_80123 == 32'h0000_0004 ? array_update_81471 : array_update_81461[4];
  assign array_update_81473[5] = add_80123 == 32'h0000_0005 ? array_update_81471 : array_update_81461[5];
  assign array_update_81473[6] = add_80123 == 32'h0000_0006 ? array_update_81471 : array_update_81461[6];
  assign array_update_81473[7] = add_80123 == 32'h0000_0007 ? array_update_81471 : array_update_81461[7];
  assign array_update_81473[8] = add_80123 == 32'h0000_0008 ? array_update_81471 : array_update_81461[8];
  assign array_update_81473[9] = add_80123 == 32'h0000_0009 ? array_update_81471 : array_update_81461[9];
  assign add_81474 = add_80123 + 32'h0000_0001;
  assign array_index_81475 = array_update_81473[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign literal_81477 = 32'h0000_0000;
  assign array_update_81478[0] = literal_81477 == 32'h0000_0000 ? 32'h0000_0000 : array_index_81475[0];
  assign array_update_81478[1] = literal_81477 == 32'h0000_0001 ? 32'h0000_0000 : array_index_81475[1];
  assign array_update_81478[2] = literal_81477 == 32'h0000_0002 ? 32'h0000_0000 : array_index_81475[2];
  assign array_update_81478[3] = literal_81477 == 32'h0000_0003 ? 32'h0000_0000 : array_index_81475[3];
  assign array_update_81478[4] = literal_81477 == 32'h0000_0004 ? 32'h0000_0000 : array_index_81475[4];
  assign array_update_81478[5] = literal_81477 == 32'h0000_0005 ? 32'h0000_0000 : array_index_81475[5];
  assign array_update_81478[6] = literal_81477 == 32'h0000_0006 ? 32'h0000_0000 : array_index_81475[6];
  assign array_update_81478[7] = literal_81477 == 32'h0000_0007 ? 32'h0000_0000 : array_index_81475[7];
  assign array_update_81478[8] = literal_81477 == 32'h0000_0008 ? 32'h0000_0000 : array_index_81475[8];
  assign array_update_81478[9] = literal_81477 == 32'h0000_0009 ? 32'h0000_0000 : array_index_81475[9];
  assign literal_81479 = 32'h0000_0000;
  assign array_update_81480[0] = add_81474 == 32'h0000_0000 ? array_update_81478 : array_update_81473[0];
  assign array_update_81480[1] = add_81474 == 32'h0000_0001 ? array_update_81478 : array_update_81473[1];
  assign array_update_81480[2] = add_81474 == 32'h0000_0002 ? array_update_81478 : array_update_81473[2];
  assign array_update_81480[3] = add_81474 == 32'h0000_0003 ? array_update_81478 : array_update_81473[3];
  assign array_update_81480[4] = add_81474 == 32'h0000_0004 ? array_update_81478 : array_update_81473[4];
  assign array_update_81480[5] = add_81474 == 32'h0000_0005 ? array_update_81478 : array_update_81473[5];
  assign array_update_81480[6] = add_81474 == 32'h0000_0006 ? array_update_81478 : array_update_81473[6];
  assign array_update_81480[7] = add_81474 == 32'h0000_0007 ? array_update_81478 : array_update_81473[7];
  assign array_update_81480[8] = add_81474 == 32'h0000_0008 ? array_update_81478 : array_update_81473[8];
  assign array_update_81480[9] = add_81474 == 32'h0000_0009 ? array_update_81478 : array_update_81473[9];
  assign array_index_81481 = array_update_72020[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign array_index_81482 = array_update_72021[literal_81479 > 32'h0000_0009 ? 4'h9 : literal_81479[3:0]];
  assign array_index_81483 = array_update_81480[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_81487 = smul32b_32b_x_32b(array_index_81481[literal_81479 > 32'h0000_0009 ? 4'h9 : literal_81479[3:0]], array_index_81482[literal_81477 > 32'h0000_0009 ? 4'h9 : literal_81477[3:0]]);
  assign add_81489 = array_index_81483[literal_81477 > 32'h0000_0009 ? 4'h9 : literal_81477[3:0]] + smul_81487;
  assign array_update_81491[0] = literal_81477 == 32'h0000_0000 ? add_81489 : array_index_81483[0];
  assign array_update_81491[1] = literal_81477 == 32'h0000_0001 ? add_81489 : array_index_81483[1];
  assign array_update_81491[2] = literal_81477 == 32'h0000_0002 ? add_81489 : array_index_81483[2];
  assign array_update_81491[3] = literal_81477 == 32'h0000_0003 ? add_81489 : array_index_81483[3];
  assign array_update_81491[4] = literal_81477 == 32'h0000_0004 ? add_81489 : array_index_81483[4];
  assign array_update_81491[5] = literal_81477 == 32'h0000_0005 ? add_81489 : array_index_81483[5];
  assign array_update_81491[6] = literal_81477 == 32'h0000_0006 ? add_81489 : array_index_81483[6];
  assign array_update_81491[7] = literal_81477 == 32'h0000_0007 ? add_81489 : array_index_81483[7];
  assign array_update_81491[8] = literal_81477 == 32'h0000_0008 ? add_81489 : array_index_81483[8];
  assign array_update_81491[9] = literal_81477 == 32'h0000_0009 ? add_81489 : array_index_81483[9];
  assign add_81492 = literal_81479 + 32'h0000_0001;
  assign array_update_81493[0] = add_81474 == 32'h0000_0000 ? array_update_81491 : array_update_81480[0];
  assign array_update_81493[1] = add_81474 == 32'h0000_0001 ? array_update_81491 : array_update_81480[1];
  assign array_update_81493[2] = add_81474 == 32'h0000_0002 ? array_update_81491 : array_update_81480[2];
  assign array_update_81493[3] = add_81474 == 32'h0000_0003 ? array_update_81491 : array_update_81480[3];
  assign array_update_81493[4] = add_81474 == 32'h0000_0004 ? array_update_81491 : array_update_81480[4];
  assign array_update_81493[5] = add_81474 == 32'h0000_0005 ? array_update_81491 : array_update_81480[5];
  assign array_update_81493[6] = add_81474 == 32'h0000_0006 ? array_update_81491 : array_update_81480[6];
  assign array_update_81493[7] = add_81474 == 32'h0000_0007 ? array_update_81491 : array_update_81480[7];
  assign array_update_81493[8] = add_81474 == 32'h0000_0008 ? array_update_81491 : array_update_81480[8];
  assign array_update_81493[9] = add_81474 == 32'h0000_0009 ? array_update_81491 : array_update_81480[9];
  assign array_index_81495 = array_update_72021[add_81492 > 32'h0000_0009 ? 4'h9 : add_81492[3:0]];
  assign array_index_81496 = array_update_81493[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_81500 = smul32b_32b_x_32b(array_index_81481[add_81492 > 32'h0000_0009 ? 4'h9 : add_81492[3:0]], array_index_81495[literal_81477 > 32'h0000_0009 ? 4'h9 : literal_81477[3:0]]);
  assign add_81502 = array_index_81496[literal_81477 > 32'h0000_0009 ? 4'h9 : literal_81477[3:0]] + smul_81500;
  assign array_update_81504[0] = literal_81477 == 32'h0000_0000 ? add_81502 : array_index_81496[0];
  assign array_update_81504[1] = literal_81477 == 32'h0000_0001 ? add_81502 : array_index_81496[1];
  assign array_update_81504[2] = literal_81477 == 32'h0000_0002 ? add_81502 : array_index_81496[2];
  assign array_update_81504[3] = literal_81477 == 32'h0000_0003 ? add_81502 : array_index_81496[3];
  assign array_update_81504[4] = literal_81477 == 32'h0000_0004 ? add_81502 : array_index_81496[4];
  assign array_update_81504[5] = literal_81477 == 32'h0000_0005 ? add_81502 : array_index_81496[5];
  assign array_update_81504[6] = literal_81477 == 32'h0000_0006 ? add_81502 : array_index_81496[6];
  assign array_update_81504[7] = literal_81477 == 32'h0000_0007 ? add_81502 : array_index_81496[7];
  assign array_update_81504[8] = literal_81477 == 32'h0000_0008 ? add_81502 : array_index_81496[8];
  assign array_update_81504[9] = literal_81477 == 32'h0000_0009 ? add_81502 : array_index_81496[9];
  assign add_81505 = add_81492 + 32'h0000_0001;
  assign array_update_81506[0] = add_81474 == 32'h0000_0000 ? array_update_81504 : array_update_81493[0];
  assign array_update_81506[1] = add_81474 == 32'h0000_0001 ? array_update_81504 : array_update_81493[1];
  assign array_update_81506[2] = add_81474 == 32'h0000_0002 ? array_update_81504 : array_update_81493[2];
  assign array_update_81506[3] = add_81474 == 32'h0000_0003 ? array_update_81504 : array_update_81493[3];
  assign array_update_81506[4] = add_81474 == 32'h0000_0004 ? array_update_81504 : array_update_81493[4];
  assign array_update_81506[5] = add_81474 == 32'h0000_0005 ? array_update_81504 : array_update_81493[5];
  assign array_update_81506[6] = add_81474 == 32'h0000_0006 ? array_update_81504 : array_update_81493[6];
  assign array_update_81506[7] = add_81474 == 32'h0000_0007 ? array_update_81504 : array_update_81493[7];
  assign array_update_81506[8] = add_81474 == 32'h0000_0008 ? array_update_81504 : array_update_81493[8];
  assign array_update_81506[9] = add_81474 == 32'h0000_0009 ? array_update_81504 : array_update_81493[9];
  assign array_index_81508 = array_update_72021[add_81505 > 32'h0000_0009 ? 4'h9 : add_81505[3:0]];
  assign array_index_81509 = array_update_81506[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_81513 = smul32b_32b_x_32b(array_index_81481[add_81505 > 32'h0000_0009 ? 4'h9 : add_81505[3:0]], array_index_81508[literal_81477 > 32'h0000_0009 ? 4'h9 : literal_81477[3:0]]);
  assign add_81515 = array_index_81509[literal_81477 > 32'h0000_0009 ? 4'h9 : literal_81477[3:0]] + smul_81513;
  assign array_update_81517[0] = literal_81477 == 32'h0000_0000 ? add_81515 : array_index_81509[0];
  assign array_update_81517[1] = literal_81477 == 32'h0000_0001 ? add_81515 : array_index_81509[1];
  assign array_update_81517[2] = literal_81477 == 32'h0000_0002 ? add_81515 : array_index_81509[2];
  assign array_update_81517[3] = literal_81477 == 32'h0000_0003 ? add_81515 : array_index_81509[3];
  assign array_update_81517[4] = literal_81477 == 32'h0000_0004 ? add_81515 : array_index_81509[4];
  assign array_update_81517[5] = literal_81477 == 32'h0000_0005 ? add_81515 : array_index_81509[5];
  assign array_update_81517[6] = literal_81477 == 32'h0000_0006 ? add_81515 : array_index_81509[6];
  assign array_update_81517[7] = literal_81477 == 32'h0000_0007 ? add_81515 : array_index_81509[7];
  assign array_update_81517[8] = literal_81477 == 32'h0000_0008 ? add_81515 : array_index_81509[8];
  assign array_update_81517[9] = literal_81477 == 32'h0000_0009 ? add_81515 : array_index_81509[9];
  assign add_81518 = add_81505 + 32'h0000_0001;
  assign array_update_81519[0] = add_81474 == 32'h0000_0000 ? array_update_81517 : array_update_81506[0];
  assign array_update_81519[1] = add_81474 == 32'h0000_0001 ? array_update_81517 : array_update_81506[1];
  assign array_update_81519[2] = add_81474 == 32'h0000_0002 ? array_update_81517 : array_update_81506[2];
  assign array_update_81519[3] = add_81474 == 32'h0000_0003 ? array_update_81517 : array_update_81506[3];
  assign array_update_81519[4] = add_81474 == 32'h0000_0004 ? array_update_81517 : array_update_81506[4];
  assign array_update_81519[5] = add_81474 == 32'h0000_0005 ? array_update_81517 : array_update_81506[5];
  assign array_update_81519[6] = add_81474 == 32'h0000_0006 ? array_update_81517 : array_update_81506[6];
  assign array_update_81519[7] = add_81474 == 32'h0000_0007 ? array_update_81517 : array_update_81506[7];
  assign array_update_81519[8] = add_81474 == 32'h0000_0008 ? array_update_81517 : array_update_81506[8];
  assign array_update_81519[9] = add_81474 == 32'h0000_0009 ? array_update_81517 : array_update_81506[9];
  assign array_index_81521 = array_update_72021[add_81518 > 32'h0000_0009 ? 4'h9 : add_81518[3:0]];
  assign array_index_81522 = array_update_81519[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_81526 = smul32b_32b_x_32b(array_index_81481[add_81518 > 32'h0000_0009 ? 4'h9 : add_81518[3:0]], array_index_81521[literal_81477 > 32'h0000_0009 ? 4'h9 : literal_81477[3:0]]);
  assign add_81528 = array_index_81522[literal_81477 > 32'h0000_0009 ? 4'h9 : literal_81477[3:0]] + smul_81526;
  assign array_update_81530[0] = literal_81477 == 32'h0000_0000 ? add_81528 : array_index_81522[0];
  assign array_update_81530[1] = literal_81477 == 32'h0000_0001 ? add_81528 : array_index_81522[1];
  assign array_update_81530[2] = literal_81477 == 32'h0000_0002 ? add_81528 : array_index_81522[2];
  assign array_update_81530[3] = literal_81477 == 32'h0000_0003 ? add_81528 : array_index_81522[3];
  assign array_update_81530[4] = literal_81477 == 32'h0000_0004 ? add_81528 : array_index_81522[4];
  assign array_update_81530[5] = literal_81477 == 32'h0000_0005 ? add_81528 : array_index_81522[5];
  assign array_update_81530[6] = literal_81477 == 32'h0000_0006 ? add_81528 : array_index_81522[6];
  assign array_update_81530[7] = literal_81477 == 32'h0000_0007 ? add_81528 : array_index_81522[7];
  assign array_update_81530[8] = literal_81477 == 32'h0000_0008 ? add_81528 : array_index_81522[8];
  assign array_update_81530[9] = literal_81477 == 32'h0000_0009 ? add_81528 : array_index_81522[9];
  assign add_81531 = add_81518 + 32'h0000_0001;
  assign array_update_81532[0] = add_81474 == 32'h0000_0000 ? array_update_81530 : array_update_81519[0];
  assign array_update_81532[1] = add_81474 == 32'h0000_0001 ? array_update_81530 : array_update_81519[1];
  assign array_update_81532[2] = add_81474 == 32'h0000_0002 ? array_update_81530 : array_update_81519[2];
  assign array_update_81532[3] = add_81474 == 32'h0000_0003 ? array_update_81530 : array_update_81519[3];
  assign array_update_81532[4] = add_81474 == 32'h0000_0004 ? array_update_81530 : array_update_81519[4];
  assign array_update_81532[5] = add_81474 == 32'h0000_0005 ? array_update_81530 : array_update_81519[5];
  assign array_update_81532[6] = add_81474 == 32'h0000_0006 ? array_update_81530 : array_update_81519[6];
  assign array_update_81532[7] = add_81474 == 32'h0000_0007 ? array_update_81530 : array_update_81519[7];
  assign array_update_81532[8] = add_81474 == 32'h0000_0008 ? array_update_81530 : array_update_81519[8];
  assign array_update_81532[9] = add_81474 == 32'h0000_0009 ? array_update_81530 : array_update_81519[9];
  assign array_index_81534 = array_update_72021[add_81531 > 32'h0000_0009 ? 4'h9 : add_81531[3:0]];
  assign array_index_81535 = array_update_81532[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_81539 = smul32b_32b_x_32b(array_index_81481[add_81531 > 32'h0000_0009 ? 4'h9 : add_81531[3:0]], array_index_81534[literal_81477 > 32'h0000_0009 ? 4'h9 : literal_81477[3:0]]);
  assign add_81541 = array_index_81535[literal_81477 > 32'h0000_0009 ? 4'h9 : literal_81477[3:0]] + smul_81539;
  assign array_update_81543[0] = literal_81477 == 32'h0000_0000 ? add_81541 : array_index_81535[0];
  assign array_update_81543[1] = literal_81477 == 32'h0000_0001 ? add_81541 : array_index_81535[1];
  assign array_update_81543[2] = literal_81477 == 32'h0000_0002 ? add_81541 : array_index_81535[2];
  assign array_update_81543[3] = literal_81477 == 32'h0000_0003 ? add_81541 : array_index_81535[3];
  assign array_update_81543[4] = literal_81477 == 32'h0000_0004 ? add_81541 : array_index_81535[4];
  assign array_update_81543[5] = literal_81477 == 32'h0000_0005 ? add_81541 : array_index_81535[5];
  assign array_update_81543[6] = literal_81477 == 32'h0000_0006 ? add_81541 : array_index_81535[6];
  assign array_update_81543[7] = literal_81477 == 32'h0000_0007 ? add_81541 : array_index_81535[7];
  assign array_update_81543[8] = literal_81477 == 32'h0000_0008 ? add_81541 : array_index_81535[8];
  assign array_update_81543[9] = literal_81477 == 32'h0000_0009 ? add_81541 : array_index_81535[9];
  assign add_81544 = add_81531 + 32'h0000_0001;
  assign array_update_81545[0] = add_81474 == 32'h0000_0000 ? array_update_81543 : array_update_81532[0];
  assign array_update_81545[1] = add_81474 == 32'h0000_0001 ? array_update_81543 : array_update_81532[1];
  assign array_update_81545[2] = add_81474 == 32'h0000_0002 ? array_update_81543 : array_update_81532[2];
  assign array_update_81545[3] = add_81474 == 32'h0000_0003 ? array_update_81543 : array_update_81532[3];
  assign array_update_81545[4] = add_81474 == 32'h0000_0004 ? array_update_81543 : array_update_81532[4];
  assign array_update_81545[5] = add_81474 == 32'h0000_0005 ? array_update_81543 : array_update_81532[5];
  assign array_update_81545[6] = add_81474 == 32'h0000_0006 ? array_update_81543 : array_update_81532[6];
  assign array_update_81545[7] = add_81474 == 32'h0000_0007 ? array_update_81543 : array_update_81532[7];
  assign array_update_81545[8] = add_81474 == 32'h0000_0008 ? array_update_81543 : array_update_81532[8];
  assign array_update_81545[9] = add_81474 == 32'h0000_0009 ? array_update_81543 : array_update_81532[9];
  assign array_index_81547 = array_update_72021[add_81544 > 32'h0000_0009 ? 4'h9 : add_81544[3:0]];
  assign array_index_81548 = array_update_81545[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_81552 = smul32b_32b_x_32b(array_index_81481[add_81544 > 32'h0000_0009 ? 4'h9 : add_81544[3:0]], array_index_81547[literal_81477 > 32'h0000_0009 ? 4'h9 : literal_81477[3:0]]);
  assign add_81554 = array_index_81548[literal_81477 > 32'h0000_0009 ? 4'h9 : literal_81477[3:0]] + smul_81552;
  assign array_update_81556[0] = literal_81477 == 32'h0000_0000 ? add_81554 : array_index_81548[0];
  assign array_update_81556[1] = literal_81477 == 32'h0000_0001 ? add_81554 : array_index_81548[1];
  assign array_update_81556[2] = literal_81477 == 32'h0000_0002 ? add_81554 : array_index_81548[2];
  assign array_update_81556[3] = literal_81477 == 32'h0000_0003 ? add_81554 : array_index_81548[3];
  assign array_update_81556[4] = literal_81477 == 32'h0000_0004 ? add_81554 : array_index_81548[4];
  assign array_update_81556[5] = literal_81477 == 32'h0000_0005 ? add_81554 : array_index_81548[5];
  assign array_update_81556[6] = literal_81477 == 32'h0000_0006 ? add_81554 : array_index_81548[6];
  assign array_update_81556[7] = literal_81477 == 32'h0000_0007 ? add_81554 : array_index_81548[7];
  assign array_update_81556[8] = literal_81477 == 32'h0000_0008 ? add_81554 : array_index_81548[8];
  assign array_update_81556[9] = literal_81477 == 32'h0000_0009 ? add_81554 : array_index_81548[9];
  assign add_81557 = add_81544 + 32'h0000_0001;
  assign array_update_81558[0] = add_81474 == 32'h0000_0000 ? array_update_81556 : array_update_81545[0];
  assign array_update_81558[1] = add_81474 == 32'h0000_0001 ? array_update_81556 : array_update_81545[1];
  assign array_update_81558[2] = add_81474 == 32'h0000_0002 ? array_update_81556 : array_update_81545[2];
  assign array_update_81558[3] = add_81474 == 32'h0000_0003 ? array_update_81556 : array_update_81545[3];
  assign array_update_81558[4] = add_81474 == 32'h0000_0004 ? array_update_81556 : array_update_81545[4];
  assign array_update_81558[5] = add_81474 == 32'h0000_0005 ? array_update_81556 : array_update_81545[5];
  assign array_update_81558[6] = add_81474 == 32'h0000_0006 ? array_update_81556 : array_update_81545[6];
  assign array_update_81558[7] = add_81474 == 32'h0000_0007 ? array_update_81556 : array_update_81545[7];
  assign array_update_81558[8] = add_81474 == 32'h0000_0008 ? array_update_81556 : array_update_81545[8];
  assign array_update_81558[9] = add_81474 == 32'h0000_0009 ? array_update_81556 : array_update_81545[9];
  assign array_index_81560 = array_update_72021[add_81557 > 32'h0000_0009 ? 4'h9 : add_81557[3:0]];
  assign array_index_81561 = array_update_81558[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_81565 = smul32b_32b_x_32b(array_index_81481[add_81557 > 32'h0000_0009 ? 4'h9 : add_81557[3:0]], array_index_81560[literal_81477 > 32'h0000_0009 ? 4'h9 : literal_81477[3:0]]);
  assign add_81567 = array_index_81561[literal_81477 > 32'h0000_0009 ? 4'h9 : literal_81477[3:0]] + smul_81565;
  assign array_update_81569[0] = literal_81477 == 32'h0000_0000 ? add_81567 : array_index_81561[0];
  assign array_update_81569[1] = literal_81477 == 32'h0000_0001 ? add_81567 : array_index_81561[1];
  assign array_update_81569[2] = literal_81477 == 32'h0000_0002 ? add_81567 : array_index_81561[2];
  assign array_update_81569[3] = literal_81477 == 32'h0000_0003 ? add_81567 : array_index_81561[3];
  assign array_update_81569[4] = literal_81477 == 32'h0000_0004 ? add_81567 : array_index_81561[4];
  assign array_update_81569[5] = literal_81477 == 32'h0000_0005 ? add_81567 : array_index_81561[5];
  assign array_update_81569[6] = literal_81477 == 32'h0000_0006 ? add_81567 : array_index_81561[6];
  assign array_update_81569[7] = literal_81477 == 32'h0000_0007 ? add_81567 : array_index_81561[7];
  assign array_update_81569[8] = literal_81477 == 32'h0000_0008 ? add_81567 : array_index_81561[8];
  assign array_update_81569[9] = literal_81477 == 32'h0000_0009 ? add_81567 : array_index_81561[9];
  assign add_81570 = add_81557 + 32'h0000_0001;
  assign array_update_81571[0] = add_81474 == 32'h0000_0000 ? array_update_81569 : array_update_81558[0];
  assign array_update_81571[1] = add_81474 == 32'h0000_0001 ? array_update_81569 : array_update_81558[1];
  assign array_update_81571[2] = add_81474 == 32'h0000_0002 ? array_update_81569 : array_update_81558[2];
  assign array_update_81571[3] = add_81474 == 32'h0000_0003 ? array_update_81569 : array_update_81558[3];
  assign array_update_81571[4] = add_81474 == 32'h0000_0004 ? array_update_81569 : array_update_81558[4];
  assign array_update_81571[5] = add_81474 == 32'h0000_0005 ? array_update_81569 : array_update_81558[5];
  assign array_update_81571[6] = add_81474 == 32'h0000_0006 ? array_update_81569 : array_update_81558[6];
  assign array_update_81571[7] = add_81474 == 32'h0000_0007 ? array_update_81569 : array_update_81558[7];
  assign array_update_81571[8] = add_81474 == 32'h0000_0008 ? array_update_81569 : array_update_81558[8];
  assign array_update_81571[9] = add_81474 == 32'h0000_0009 ? array_update_81569 : array_update_81558[9];
  assign array_index_81573 = array_update_72021[add_81570 > 32'h0000_0009 ? 4'h9 : add_81570[3:0]];
  assign array_index_81574 = array_update_81571[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_81578 = smul32b_32b_x_32b(array_index_81481[add_81570 > 32'h0000_0009 ? 4'h9 : add_81570[3:0]], array_index_81573[literal_81477 > 32'h0000_0009 ? 4'h9 : literal_81477[3:0]]);
  assign add_81580 = array_index_81574[literal_81477 > 32'h0000_0009 ? 4'h9 : literal_81477[3:0]] + smul_81578;
  assign array_update_81582[0] = literal_81477 == 32'h0000_0000 ? add_81580 : array_index_81574[0];
  assign array_update_81582[1] = literal_81477 == 32'h0000_0001 ? add_81580 : array_index_81574[1];
  assign array_update_81582[2] = literal_81477 == 32'h0000_0002 ? add_81580 : array_index_81574[2];
  assign array_update_81582[3] = literal_81477 == 32'h0000_0003 ? add_81580 : array_index_81574[3];
  assign array_update_81582[4] = literal_81477 == 32'h0000_0004 ? add_81580 : array_index_81574[4];
  assign array_update_81582[5] = literal_81477 == 32'h0000_0005 ? add_81580 : array_index_81574[5];
  assign array_update_81582[6] = literal_81477 == 32'h0000_0006 ? add_81580 : array_index_81574[6];
  assign array_update_81582[7] = literal_81477 == 32'h0000_0007 ? add_81580 : array_index_81574[7];
  assign array_update_81582[8] = literal_81477 == 32'h0000_0008 ? add_81580 : array_index_81574[8];
  assign array_update_81582[9] = literal_81477 == 32'h0000_0009 ? add_81580 : array_index_81574[9];
  assign add_81583 = add_81570 + 32'h0000_0001;
  assign array_update_81584[0] = add_81474 == 32'h0000_0000 ? array_update_81582 : array_update_81571[0];
  assign array_update_81584[1] = add_81474 == 32'h0000_0001 ? array_update_81582 : array_update_81571[1];
  assign array_update_81584[2] = add_81474 == 32'h0000_0002 ? array_update_81582 : array_update_81571[2];
  assign array_update_81584[3] = add_81474 == 32'h0000_0003 ? array_update_81582 : array_update_81571[3];
  assign array_update_81584[4] = add_81474 == 32'h0000_0004 ? array_update_81582 : array_update_81571[4];
  assign array_update_81584[5] = add_81474 == 32'h0000_0005 ? array_update_81582 : array_update_81571[5];
  assign array_update_81584[6] = add_81474 == 32'h0000_0006 ? array_update_81582 : array_update_81571[6];
  assign array_update_81584[7] = add_81474 == 32'h0000_0007 ? array_update_81582 : array_update_81571[7];
  assign array_update_81584[8] = add_81474 == 32'h0000_0008 ? array_update_81582 : array_update_81571[8];
  assign array_update_81584[9] = add_81474 == 32'h0000_0009 ? array_update_81582 : array_update_81571[9];
  assign array_index_81586 = array_update_72021[add_81583 > 32'h0000_0009 ? 4'h9 : add_81583[3:0]];
  assign array_index_81587 = array_update_81584[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_81591 = smul32b_32b_x_32b(array_index_81481[add_81583 > 32'h0000_0009 ? 4'h9 : add_81583[3:0]], array_index_81586[literal_81477 > 32'h0000_0009 ? 4'h9 : literal_81477[3:0]]);
  assign add_81593 = array_index_81587[literal_81477 > 32'h0000_0009 ? 4'h9 : literal_81477[3:0]] + smul_81591;
  assign array_update_81595[0] = literal_81477 == 32'h0000_0000 ? add_81593 : array_index_81587[0];
  assign array_update_81595[1] = literal_81477 == 32'h0000_0001 ? add_81593 : array_index_81587[1];
  assign array_update_81595[2] = literal_81477 == 32'h0000_0002 ? add_81593 : array_index_81587[2];
  assign array_update_81595[3] = literal_81477 == 32'h0000_0003 ? add_81593 : array_index_81587[3];
  assign array_update_81595[4] = literal_81477 == 32'h0000_0004 ? add_81593 : array_index_81587[4];
  assign array_update_81595[5] = literal_81477 == 32'h0000_0005 ? add_81593 : array_index_81587[5];
  assign array_update_81595[6] = literal_81477 == 32'h0000_0006 ? add_81593 : array_index_81587[6];
  assign array_update_81595[7] = literal_81477 == 32'h0000_0007 ? add_81593 : array_index_81587[7];
  assign array_update_81595[8] = literal_81477 == 32'h0000_0008 ? add_81593 : array_index_81587[8];
  assign array_update_81595[9] = literal_81477 == 32'h0000_0009 ? add_81593 : array_index_81587[9];
  assign add_81596 = add_81583 + 32'h0000_0001;
  assign array_update_81597[0] = add_81474 == 32'h0000_0000 ? array_update_81595 : array_update_81584[0];
  assign array_update_81597[1] = add_81474 == 32'h0000_0001 ? array_update_81595 : array_update_81584[1];
  assign array_update_81597[2] = add_81474 == 32'h0000_0002 ? array_update_81595 : array_update_81584[2];
  assign array_update_81597[3] = add_81474 == 32'h0000_0003 ? array_update_81595 : array_update_81584[3];
  assign array_update_81597[4] = add_81474 == 32'h0000_0004 ? array_update_81595 : array_update_81584[4];
  assign array_update_81597[5] = add_81474 == 32'h0000_0005 ? array_update_81595 : array_update_81584[5];
  assign array_update_81597[6] = add_81474 == 32'h0000_0006 ? array_update_81595 : array_update_81584[6];
  assign array_update_81597[7] = add_81474 == 32'h0000_0007 ? array_update_81595 : array_update_81584[7];
  assign array_update_81597[8] = add_81474 == 32'h0000_0008 ? array_update_81595 : array_update_81584[8];
  assign array_update_81597[9] = add_81474 == 32'h0000_0009 ? array_update_81595 : array_update_81584[9];
  assign array_index_81599 = array_update_72021[add_81596 > 32'h0000_0009 ? 4'h9 : add_81596[3:0]];
  assign array_index_81600 = array_update_81597[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_81604 = smul32b_32b_x_32b(array_index_81481[add_81596 > 32'h0000_0009 ? 4'h9 : add_81596[3:0]], array_index_81599[literal_81477 > 32'h0000_0009 ? 4'h9 : literal_81477[3:0]]);
  assign add_81606 = array_index_81600[literal_81477 > 32'h0000_0009 ? 4'h9 : literal_81477[3:0]] + smul_81604;
  assign array_update_81607[0] = literal_81477 == 32'h0000_0000 ? add_81606 : array_index_81600[0];
  assign array_update_81607[1] = literal_81477 == 32'h0000_0001 ? add_81606 : array_index_81600[1];
  assign array_update_81607[2] = literal_81477 == 32'h0000_0002 ? add_81606 : array_index_81600[2];
  assign array_update_81607[3] = literal_81477 == 32'h0000_0003 ? add_81606 : array_index_81600[3];
  assign array_update_81607[4] = literal_81477 == 32'h0000_0004 ? add_81606 : array_index_81600[4];
  assign array_update_81607[5] = literal_81477 == 32'h0000_0005 ? add_81606 : array_index_81600[5];
  assign array_update_81607[6] = literal_81477 == 32'h0000_0006 ? add_81606 : array_index_81600[6];
  assign array_update_81607[7] = literal_81477 == 32'h0000_0007 ? add_81606 : array_index_81600[7];
  assign array_update_81607[8] = literal_81477 == 32'h0000_0008 ? add_81606 : array_index_81600[8];
  assign array_update_81607[9] = literal_81477 == 32'h0000_0009 ? add_81606 : array_index_81600[9];
  assign array_update_81608[0] = add_81474 == 32'h0000_0000 ? array_update_81607 : array_update_81597[0];
  assign array_update_81608[1] = add_81474 == 32'h0000_0001 ? array_update_81607 : array_update_81597[1];
  assign array_update_81608[2] = add_81474 == 32'h0000_0002 ? array_update_81607 : array_update_81597[2];
  assign array_update_81608[3] = add_81474 == 32'h0000_0003 ? array_update_81607 : array_update_81597[3];
  assign array_update_81608[4] = add_81474 == 32'h0000_0004 ? array_update_81607 : array_update_81597[4];
  assign array_update_81608[5] = add_81474 == 32'h0000_0005 ? array_update_81607 : array_update_81597[5];
  assign array_update_81608[6] = add_81474 == 32'h0000_0006 ? array_update_81607 : array_update_81597[6];
  assign array_update_81608[7] = add_81474 == 32'h0000_0007 ? array_update_81607 : array_update_81597[7];
  assign array_update_81608[8] = add_81474 == 32'h0000_0008 ? array_update_81607 : array_update_81597[8];
  assign array_update_81608[9] = add_81474 == 32'h0000_0009 ? array_update_81607 : array_update_81597[9];
  assign array_index_81610 = array_update_81608[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign add_81612 = literal_81477 + 32'h0000_0001;
  assign array_update_81613[0] = add_81612 == 32'h0000_0000 ? 32'h0000_0000 : array_index_81610[0];
  assign array_update_81613[1] = add_81612 == 32'h0000_0001 ? 32'h0000_0000 : array_index_81610[1];
  assign array_update_81613[2] = add_81612 == 32'h0000_0002 ? 32'h0000_0000 : array_index_81610[2];
  assign array_update_81613[3] = add_81612 == 32'h0000_0003 ? 32'h0000_0000 : array_index_81610[3];
  assign array_update_81613[4] = add_81612 == 32'h0000_0004 ? 32'h0000_0000 : array_index_81610[4];
  assign array_update_81613[5] = add_81612 == 32'h0000_0005 ? 32'h0000_0000 : array_index_81610[5];
  assign array_update_81613[6] = add_81612 == 32'h0000_0006 ? 32'h0000_0000 : array_index_81610[6];
  assign array_update_81613[7] = add_81612 == 32'h0000_0007 ? 32'h0000_0000 : array_index_81610[7];
  assign array_update_81613[8] = add_81612 == 32'h0000_0008 ? 32'h0000_0000 : array_index_81610[8];
  assign array_update_81613[9] = add_81612 == 32'h0000_0009 ? 32'h0000_0000 : array_index_81610[9];
  assign literal_81614 = 32'h0000_0000;
  assign array_update_81615[0] = add_81474 == 32'h0000_0000 ? array_update_81613 : array_update_81608[0];
  assign array_update_81615[1] = add_81474 == 32'h0000_0001 ? array_update_81613 : array_update_81608[1];
  assign array_update_81615[2] = add_81474 == 32'h0000_0002 ? array_update_81613 : array_update_81608[2];
  assign array_update_81615[3] = add_81474 == 32'h0000_0003 ? array_update_81613 : array_update_81608[3];
  assign array_update_81615[4] = add_81474 == 32'h0000_0004 ? array_update_81613 : array_update_81608[4];
  assign array_update_81615[5] = add_81474 == 32'h0000_0005 ? array_update_81613 : array_update_81608[5];
  assign array_update_81615[6] = add_81474 == 32'h0000_0006 ? array_update_81613 : array_update_81608[6];
  assign array_update_81615[7] = add_81474 == 32'h0000_0007 ? array_update_81613 : array_update_81608[7];
  assign array_update_81615[8] = add_81474 == 32'h0000_0008 ? array_update_81613 : array_update_81608[8];
  assign array_update_81615[9] = add_81474 == 32'h0000_0009 ? array_update_81613 : array_update_81608[9];
  assign array_index_81617 = array_update_72021[literal_81614 > 32'h0000_0009 ? 4'h9 : literal_81614[3:0]];
  assign array_index_81618 = array_update_81615[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_81622 = smul32b_32b_x_32b(array_index_81481[literal_81614 > 32'h0000_0009 ? 4'h9 : literal_81614[3:0]], array_index_81617[add_81612 > 32'h0000_0009 ? 4'h9 : add_81612[3:0]]);
  assign add_81624 = array_index_81618[add_81612 > 32'h0000_0009 ? 4'h9 : add_81612[3:0]] + smul_81622;
  assign array_update_81626[0] = add_81612 == 32'h0000_0000 ? add_81624 : array_index_81618[0];
  assign array_update_81626[1] = add_81612 == 32'h0000_0001 ? add_81624 : array_index_81618[1];
  assign array_update_81626[2] = add_81612 == 32'h0000_0002 ? add_81624 : array_index_81618[2];
  assign array_update_81626[3] = add_81612 == 32'h0000_0003 ? add_81624 : array_index_81618[3];
  assign array_update_81626[4] = add_81612 == 32'h0000_0004 ? add_81624 : array_index_81618[4];
  assign array_update_81626[5] = add_81612 == 32'h0000_0005 ? add_81624 : array_index_81618[5];
  assign array_update_81626[6] = add_81612 == 32'h0000_0006 ? add_81624 : array_index_81618[6];
  assign array_update_81626[7] = add_81612 == 32'h0000_0007 ? add_81624 : array_index_81618[7];
  assign array_update_81626[8] = add_81612 == 32'h0000_0008 ? add_81624 : array_index_81618[8];
  assign array_update_81626[9] = add_81612 == 32'h0000_0009 ? add_81624 : array_index_81618[9];
  assign add_81627 = literal_81614 + 32'h0000_0001;
  assign array_update_81628[0] = add_81474 == 32'h0000_0000 ? array_update_81626 : array_update_81615[0];
  assign array_update_81628[1] = add_81474 == 32'h0000_0001 ? array_update_81626 : array_update_81615[1];
  assign array_update_81628[2] = add_81474 == 32'h0000_0002 ? array_update_81626 : array_update_81615[2];
  assign array_update_81628[3] = add_81474 == 32'h0000_0003 ? array_update_81626 : array_update_81615[3];
  assign array_update_81628[4] = add_81474 == 32'h0000_0004 ? array_update_81626 : array_update_81615[4];
  assign array_update_81628[5] = add_81474 == 32'h0000_0005 ? array_update_81626 : array_update_81615[5];
  assign array_update_81628[6] = add_81474 == 32'h0000_0006 ? array_update_81626 : array_update_81615[6];
  assign array_update_81628[7] = add_81474 == 32'h0000_0007 ? array_update_81626 : array_update_81615[7];
  assign array_update_81628[8] = add_81474 == 32'h0000_0008 ? array_update_81626 : array_update_81615[8];
  assign array_update_81628[9] = add_81474 == 32'h0000_0009 ? array_update_81626 : array_update_81615[9];
  assign array_index_81630 = array_update_72021[add_81627 > 32'h0000_0009 ? 4'h9 : add_81627[3:0]];
  assign array_index_81631 = array_update_81628[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_81635 = smul32b_32b_x_32b(array_index_81481[add_81627 > 32'h0000_0009 ? 4'h9 : add_81627[3:0]], array_index_81630[add_81612 > 32'h0000_0009 ? 4'h9 : add_81612[3:0]]);
  assign add_81637 = array_index_81631[add_81612 > 32'h0000_0009 ? 4'h9 : add_81612[3:0]] + smul_81635;
  assign array_update_81639[0] = add_81612 == 32'h0000_0000 ? add_81637 : array_index_81631[0];
  assign array_update_81639[1] = add_81612 == 32'h0000_0001 ? add_81637 : array_index_81631[1];
  assign array_update_81639[2] = add_81612 == 32'h0000_0002 ? add_81637 : array_index_81631[2];
  assign array_update_81639[3] = add_81612 == 32'h0000_0003 ? add_81637 : array_index_81631[3];
  assign array_update_81639[4] = add_81612 == 32'h0000_0004 ? add_81637 : array_index_81631[4];
  assign array_update_81639[5] = add_81612 == 32'h0000_0005 ? add_81637 : array_index_81631[5];
  assign array_update_81639[6] = add_81612 == 32'h0000_0006 ? add_81637 : array_index_81631[6];
  assign array_update_81639[7] = add_81612 == 32'h0000_0007 ? add_81637 : array_index_81631[7];
  assign array_update_81639[8] = add_81612 == 32'h0000_0008 ? add_81637 : array_index_81631[8];
  assign array_update_81639[9] = add_81612 == 32'h0000_0009 ? add_81637 : array_index_81631[9];
  assign add_81640 = add_81627 + 32'h0000_0001;
  assign array_update_81641[0] = add_81474 == 32'h0000_0000 ? array_update_81639 : array_update_81628[0];
  assign array_update_81641[1] = add_81474 == 32'h0000_0001 ? array_update_81639 : array_update_81628[1];
  assign array_update_81641[2] = add_81474 == 32'h0000_0002 ? array_update_81639 : array_update_81628[2];
  assign array_update_81641[3] = add_81474 == 32'h0000_0003 ? array_update_81639 : array_update_81628[3];
  assign array_update_81641[4] = add_81474 == 32'h0000_0004 ? array_update_81639 : array_update_81628[4];
  assign array_update_81641[5] = add_81474 == 32'h0000_0005 ? array_update_81639 : array_update_81628[5];
  assign array_update_81641[6] = add_81474 == 32'h0000_0006 ? array_update_81639 : array_update_81628[6];
  assign array_update_81641[7] = add_81474 == 32'h0000_0007 ? array_update_81639 : array_update_81628[7];
  assign array_update_81641[8] = add_81474 == 32'h0000_0008 ? array_update_81639 : array_update_81628[8];
  assign array_update_81641[9] = add_81474 == 32'h0000_0009 ? array_update_81639 : array_update_81628[9];
  assign array_index_81643 = array_update_72021[add_81640 > 32'h0000_0009 ? 4'h9 : add_81640[3:0]];
  assign array_index_81644 = array_update_81641[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_81648 = smul32b_32b_x_32b(array_index_81481[add_81640 > 32'h0000_0009 ? 4'h9 : add_81640[3:0]], array_index_81643[add_81612 > 32'h0000_0009 ? 4'h9 : add_81612[3:0]]);
  assign add_81650 = array_index_81644[add_81612 > 32'h0000_0009 ? 4'h9 : add_81612[3:0]] + smul_81648;
  assign array_update_81652[0] = add_81612 == 32'h0000_0000 ? add_81650 : array_index_81644[0];
  assign array_update_81652[1] = add_81612 == 32'h0000_0001 ? add_81650 : array_index_81644[1];
  assign array_update_81652[2] = add_81612 == 32'h0000_0002 ? add_81650 : array_index_81644[2];
  assign array_update_81652[3] = add_81612 == 32'h0000_0003 ? add_81650 : array_index_81644[3];
  assign array_update_81652[4] = add_81612 == 32'h0000_0004 ? add_81650 : array_index_81644[4];
  assign array_update_81652[5] = add_81612 == 32'h0000_0005 ? add_81650 : array_index_81644[5];
  assign array_update_81652[6] = add_81612 == 32'h0000_0006 ? add_81650 : array_index_81644[6];
  assign array_update_81652[7] = add_81612 == 32'h0000_0007 ? add_81650 : array_index_81644[7];
  assign array_update_81652[8] = add_81612 == 32'h0000_0008 ? add_81650 : array_index_81644[8];
  assign array_update_81652[9] = add_81612 == 32'h0000_0009 ? add_81650 : array_index_81644[9];
  assign add_81653 = add_81640 + 32'h0000_0001;
  assign array_update_81654[0] = add_81474 == 32'h0000_0000 ? array_update_81652 : array_update_81641[0];
  assign array_update_81654[1] = add_81474 == 32'h0000_0001 ? array_update_81652 : array_update_81641[1];
  assign array_update_81654[2] = add_81474 == 32'h0000_0002 ? array_update_81652 : array_update_81641[2];
  assign array_update_81654[3] = add_81474 == 32'h0000_0003 ? array_update_81652 : array_update_81641[3];
  assign array_update_81654[4] = add_81474 == 32'h0000_0004 ? array_update_81652 : array_update_81641[4];
  assign array_update_81654[5] = add_81474 == 32'h0000_0005 ? array_update_81652 : array_update_81641[5];
  assign array_update_81654[6] = add_81474 == 32'h0000_0006 ? array_update_81652 : array_update_81641[6];
  assign array_update_81654[7] = add_81474 == 32'h0000_0007 ? array_update_81652 : array_update_81641[7];
  assign array_update_81654[8] = add_81474 == 32'h0000_0008 ? array_update_81652 : array_update_81641[8];
  assign array_update_81654[9] = add_81474 == 32'h0000_0009 ? array_update_81652 : array_update_81641[9];
  assign array_index_81656 = array_update_72021[add_81653 > 32'h0000_0009 ? 4'h9 : add_81653[3:0]];
  assign array_index_81657 = array_update_81654[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_81661 = smul32b_32b_x_32b(array_index_81481[add_81653 > 32'h0000_0009 ? 4'h9 : add_81653[3:0]], array_index_81656[add_81612 > 32'h0000_0009 ? 4'h9 : add_81612[3:0]]);
  assign add_81663 = array_index_81657[add_81612 > 32'h0000_0009 ? 4'h9 : add_81612[3:0]] + smul_81661;
  assign array_update_81665[0] = add_81612 == 32'h0000_0000 ? add_81663 : array_index_81657[0];
  assign array_update_81665[1] = add_81612 == 32'h0000_0001 ? add_81663 : array_index_81657[1];
  assign array_update_81665[2] = add_81612 == 32'h0000_0002 ? add_81663 : array_index_81657[2];
  assign array_update_81665[3] = add_81612 == 32'h0000_0003 ? add_81663 : array_index_81657[3];
  assign array_update_81665[4] = add_81612 == 32'h0000_0004 ? add_81663 : array_index_81657[4];
  assign array_update_81665[5] = add_81612 == 32'h0000_0005 ? add_81663 : array_index_81657[5];
  assign array_update_81665[6] = add_81612 == 32'h0000_0006 ? add_81663 : array_index_81657[6];
  assign array_update_81665[7] = add_81612 == 32'h0000_0007 ? add_81663 : array_index_81657[7];
  assign array_update_81665[8] = add_81612 == 32'h0000_0008 ? add_81663 : array_index_81657[8];
  assign array_update_81665[9] = add_81612 == 32'h0000_0009 ? add_81663 : array_index_81657[9];
  assign add_81666 = add_81653 + 32'h0000_0001;
  assign array_update_81667[0] = add_81474 == 32'h0000_0000 ? array_update_81665 : array_update_81654[0];
  assign array_update_81667[1] = add_81474 == 32'h0000_0001 ? array_update_81665 : array_update_81654[1];
  assign array_update_81667[2] = add_81474 == 32'h0000_0002 ? array_update_81665 : array_update_81654[2];
  assign array_update_81667[3] = add_81474 == 32'h0000_0003 ? array_update_81665 : array_update_81654[3];
  assign array_update_81667[4] = add_81474 == 32'h0000_0004 ? array_update_81665 : array_update_81654[4];
  assign array_update_81667[5] = add_81474 == 32'h0000_0005 ? array_update_81665 : array_update_81654[5];
  assign array_update_81667[6] = add_81474 == 32'h0000_0006 ? array_update_81665 : array_update_81654[6];
  assign array_update_81667[7] = add_81474 == 32'h0000_0007 ? array_update_81665 : array_update_81654[7];
  assign array_update_81667[8] = add_81474 == 32'h0000_0008 ? array_update_81665 : array_update_81654[8];
  assign array_update_81667[9] = add_81474 == 32'h0000_0009 ? array_update_81665 : array_update_81654[9];
  assign array_index_81669 = array_update_72021[add_81666 > 32'h0000_0009 ? 4'h9 : add_81666[3:0]];
  assign array_index_81670 = array_update_81667[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_81674 = smul32b_32b_x_32b(array_index_81481[add_81666 > 32'h0000_0009 ? 4'h9 : add_81666[3:0]], array_index_81669[add_81612 > 32'h0000_0009 ? 4'h9 : add_81612[3:0]]);
  assign add_81676 = array_index_81670[add_81612 > 32'h0000_0009 ? 4'h9 : add_81612[3:0]] + smul_81674;
  assign array_update_81678[0] = add_81612 == 32'h0000_0000 ? add_81676 : array_index_81670[0];
  assign array_update_81678[1] = add_81612 == 32'h0000_0001 ? add_81676 : array_index_81670[1];
  assign array_update_81678[2] = add_81612 == 32'h0000_0002 ? add_81676 : array_index_81670[2];
  assign array_update_81678[3] = add_81612 == 32'h0000_0003 ? add_81676 : array_index_81670[3];
  assign array_update_81678[4] = add_81612 == 32'h0000_0004 ? add_81676 : array_index_81670[4];
  assign array_update_81678[5] = add_81612 == 32'h0000_0005 ? add_81676 : array_index_81670[5];
  assign array_update_81678[6] = add_81612 == 32'h0000_0006 ? add_81676 : array_index_81670[6];
  assign array_update_81678[7] = add_81612 == 32'h0000_0007 ? add_81676 : array_index_81670[7];
  assign array_update_81678[8] = add_81612 == 32'h0000_0008 ? add_81676 : array_index_81670[8];
  assign array_update_81678[9] = add_81612 == 32'h0000_0009 ? add_81676 : array_index_81670[9];
  assign add_81679 = add_81666 + 32'h0000_0001;
  assign array_update_81680[0] = add_81474 == 32'h0000_0000 ? array_update_81678 : array_update_81667[0];
  assign array_update_81680[1] = add_81474 == 32'h0000_0001 ? array_update_81678 : array_update_81667[1];
  assign array_update_81680[2] = add_81474 == 32'h0000_0002 ? array_update_81678 : array_update_81667[2];
  assign array_update_81680[3] = add_81474 == 32'h0000_0003 ? array_update_81678 : array_update_81667[3];
  assign array_update_81680[4] = add_81474 == 32'h0000_0004 ? array_update_81678 : array_update_81667[4];
  assign array_update_81680[5] = add_81474 == 32'h0000_0005 ? array_update_81678 : array_update_81667[5];
  assign array_update_81680[6] = add_81474 == 32'h0000_0006 ? array_update_81678 : array_update_81667[6];
  assign array_update_81680[7] = add_81474 == 32'h0000_0007 ? array_update_81678 : array_update_81667[7];
  assign array_update_81680[8] = add_81474 == 32'h0000_0008 ? array_update_81678 : array_update_81667[8];
  assign array_update_81680[9] = add_81474 == 32'h0000_0009 ? array_update_81678 : array_update_81667[9];
  assign array_index_81682 = array_update_72021[add_81679 > 32'h0000_0009 ? 4'h9 : add_81679[3:0]];
  assign array_index_81683 = array_update_81680[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_81687 = smul32b_32b_x_32b(array_index_81481[add_81679 > 32'h0000_0009 ? 4'h9 : add_81679[3:0]], array_index_81682[add_81612 > 32'h0000_0009 ? 4'h9 : add_81612[3:0]]);
  assign add_81689 = array_index_81683[add_81612 > 32'h0000_0009 ? 4'h9 : add_81612[3:0]] + smul_81687;
  assign array_update_81691[0] = add_81612 == 32'h0000_0000 ? add_81689 : array_index_81683[0];
  assign array_update_81691[1] = add_81612 == 32'h0000_0001 ? add_81689 : array_index_81683[1];
  assign array_update_81691[2] = add_81612 == 32'h0000_0002 ? add_81689 : array_index_81683[2];
  assign array_update_81691[3] = add_81612 == 32'h0000_0003 ? add_81689 : array_index_81683[3];
  assign array_update_81691[4] = add_81612 == 32'h0000_0004 ? add_81689 : array_index_81683[4];
  assign array_update_81691[5] = add_81612 == 32'h0000_0005 ? add_81689 : array_index_81683[5];
  assign array_update_81691[6] = add_81612 == 32'h0000_0006 ? add_81689 : array_index_81683[6];
  assign array_update_81691[7] = add_81612 == 32'h0000_0007 ? add_81689 : array_index_81683[7];
  assign array_update_81691[8] = add_81612 == 32'h0000_0008 ? add_81689 : array_index_81683[8];
  assign array_update_81691[9] = add_81612 == 32'h0000_0009 ? add_81689 : array_index_81683[9];
  assign add_81692 = add_81679 + 32'h0000_0001;
  assign array_update_81693[0] = add_81474 == 32'h0000_0000 ? array_update_81691 : array_update_81680[0];
  assign array_update_81693[1] = add_81474 == 32'h0000_0001 ? array_update_81691 : array_update_81680[1];
  assign array_update_81693[2] = add_81474 == 32'h0000_0002 ? array_update_81691 : array_update_81680[2];
  assign array_update_81693[3] = add_81474 == 32'h0000_0003 ? array_update_81691 : array_update_81680[3];
  assign array_update_81693[4] = add_81474 == 32'h0000_0004 ? array_update_81691 : array_update_81680[4];
  assign array_update_81693[5] = add_81474 == 32'h0000_0005 ? array_update_81691 : array_update_81680[5];
  assign array_update_81693[6] = add_81474 == 32'h0000_0006 ? array_update_81691 : array_update_81680[6];
  assign array_update_81693[7] = add_81474 == 32'h0000_0007 ? array_update_81691 : array_update_81680[7];
  assign array_update_81693[8] = add_81474 == 32'h0000_0008 ? array_update_81691 : array_update_81680[8];
  assign array_update_81693[9] = add_81474 == 32'h0000_0009 ? array_update_81691 : array_update_81680[9];
  assign array_index_81695 = array_update_72021[add_81692 > 32'h0000_0009 ? 4'h9 : add_81692[3:0]];
  assign array_index_81696 = array_update_81693[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_81700 = smul32b_32b_x_32b(array_index_81481[add_81692 > 32'h0000_0009 ? 4'h9 : add_81692[3:0]], array_index_81695[add_81612 > 32'h0000_0009 ? 4'h9 : add_81612[3:0]]);
  assign add_81702 = array_index_81696[add_81612 > 32'h0000_0009 ? 4'h9 : add_81612[3:0]] + smul_81700;
  assign array_update_81704[0] = add_81612 == 32'h0000_0000 ? add_81702 : array_index_81696[0];
  assign array_update_81704[1] = add_81612 == 32'h0000_0001 ? add_81702 : array_index_81696[1];
  assign array_update_81704[2] = add_81612 == 32'h0000_0002 ? add_81702 : array_index_81696[2];
  assign array_update_81704[3] = add_81612 == 32'h0000_0003 ? add_81702 : array_index_81696[3];
  assign array_update_81704[4] = add_81612 == 32'h0000_0004 ? add_81702 : array_index_81696[4];
  assign array_update_81704[5] = add_81612 == 32'h0000_0005 ? add_81702 : array_index_81696[5];
  assign array_update_81704[6] = add_81612 == 32'h0000_0006 ? add_81702 : array_index_81696[6];
  assign array_update_81704[7] = add_81612 == 32'h0000_0007 ? add_81702 : array_index_81696[7];
  assign array_update_81704[8] = add_81612 == 32'h0000_0008 ? add_81702 : array_index_81696[8];
  assign array_update_81704[9] = add_81612 == 32'h0000_0009 ? add_81702 : array_index_81696[9];
  assign add_81705 = add_81692 + 32'h0000_0001;
  assign array_update_81706[0] = add_81474 == 32'h0000_0000 ? array_update_81704 : array_update_81693[0];
  assign array_update_81706[1] = add_81474 == 32'h0000_0001 ? array_update_81704 : array_update_81693[1];
  assign array_update_81706[2] = add_81474 == 32'h0000_0002 ? array_update_81704 : array_update_81693[2];
  assign array_update_81706[3] = add_81474 == 32'h0000_0003 ? array_update_81704 : array_update_81693[3];
  assign array_update_81706[4] = add_81474 == 32'h0000_0004 ? array_update_81704 : array_update_81693[4];
  assign array_update_81706[5] = add_81474 == 32'h0000_0005 ? array_update_81704 : array_update_81693[5];
  assign array_update_81706[6] = add_81474 == 32'h0000_0006 ? array_update_81704 : array_update_81693[6];
  assign array_update_81706[7] = add_81474 == 32'h0000_0007 ? array_update_81704 : array_update_81693[7];
  assign array_update_81706[8] = add_81474 == 32'h0000_0008 ? array_update_81704 : array_update_81693[8];
  assign array_update_81706[9] = add_81474 == 32'h0000_0009 ? array_update_81704 : array_update_81693[9];
  assign array_index_81708 = array_update_72021[add_81705 > 32'h0000_0009 ? 4'h9 : add_81705[3:0]];
  assign array_index_81709 = array_update_81706[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_81713 = smul32b_32b_x_32b(array_index_81481[add_81705 > 32'h0000_0009 ? 4'h9 : add_81705[3:0]], array_index_81708[add_81612 > 32'h0000_0009 ? 4'h9 : add_81612[3:0]]);
  assign add_81715 = array_index_81709[add_81612 > 32'h0000_0009 ? 4'h9 : add_81612[3:0]] + smul_81713;
  assign array_update_81717[0] = add_81612 == 32'h0000_0000 ? add_81715 : array_index_81709[0];
  assign array_update_81717[1] = add_81612 == 32'h0000_0001 ? add_81715 : array_index_81709[1];
  assign array_update_81717[2] = add_81612 == 32'h0000_0002 ? add_81715 : array_index_81709[2];
  assign array_update_81717[3] = add_81612 == 32'h0000_0003 ? add_81715 : array_index_81709[3];
  assign array_update_81717[4] = add_81612 == 32'h0000_0004 ? add_81715 : array_index_81709[4];
  assign array_update_81717[5] = add_81612 == 32'h0000_0005 ? add_81715 : array_index_81709[5];
  assign array_update_81717[6] = add_81612 == 32'h0000_0006 ? add_81715 : array_index_81709[6];
  assign array_update_81717[7] = add_81612 == 32'h0000_0007 ? add_81715 : array_index_81709[7];
  assign array_update_81717[8] = add_81612 == 32'h0000_0008 ? add_81715 : array_index_81709[8];
  assign array_update_81717[9] = add_81612 == 32'h0000_0009 ? add_81715 : array_index_81709[9];
  assign add_81718 = add_81705 + 32'h0000_0001;
  assign array_update_81719[0] = add_81474 == 32'h0000_0000 ? array_update_81717 : array_update_81706[0];
  assign array_update_81719[1] = add_81474 == 32'h0000_0001 ? array_update_81717 : array_update_81706[1];
  assign array_update_81719[2] = add_81474 == 32'h0000_0002 ? array_update_81717 : array_update_81706[2];
  assign array_update_81719[3] = add_81474 == 32'h0000_0003 ? array_update_81717 : array_update_81706[3];
  assign array_update_81719[4] = add_81474 == 32'h0000_0004 ? array_update_81717 : array_update_81706[4];
  assign array_update_81719[5] = add_81474 == 32'h0000_0005 ? array_update_81717 : array_update_81706[5];
  assign array_update_81719[6] = add_81474 == 32'h0000_0006 ? array_update_81717 : array_update_81706[6];
  assign array_update_81719[7] = add_81474 == 32'h0000_0007 ? array_update_81717 : array_update_81706[7];
  assign array_update_81719[8] = add_81474 == 32'h0000_0008 ? array_update_81717 : array_update_81706[8];
  assign array_update_81719[9] = add_81474 == 32'h0000_0009 ? array_update_81717 : array_update_81706[9];
  assign array_index_81721 = array_update_72021[add_81718 > 32'h0000_0009 ? 4'h9 : add_81718[3:0]];
  assign array_index_81722 = array_update_81719[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_81726 = smul32b_32b_x_32b(array_index_81481[add_81718 > 32'h0000_0009 ? 4'h9 : add_81718[3:0]], array_index_81721[add_81612 > 32'h0000_0009 ? 4'h9 : add_81612[3:0]]);
  assign add_81728 = array_index_81722[add_81612 > 32'h0000_0009 ? 4'h9 : add_81612[3:0]] + smul_81726;
  assign array_update_81730[0] = add_81612 == 32'h0000_0000 ? add_81728 : array_index_81722[0];
  assign array_update_81730[1] = add_81612 == 32'h0000_0001 ? add_81728 : array_index_81722[1];
  assign array_update_81730[2] = add_81612 == 32'h0000_0002 ? add_81728 : array_index_81722[2];
  assign array_update_81730[3] = add_81612 == 32'h0000_0003 ? add_81728 : array_index_81722[3];
  assign array_update_81730[4] = add_81612 == 32'h0000_0004 ? add_81728 : array_index_81722[4];
  assign array_update_81730[5] = add_81612 == 32'h0000_0005 ? add_81728 : array_index_81722[5];
  assign array_update_81730[6] = add_81612 == 32'h0000_0006 ? add_81728 : array_index_81722[6];
  assign array_update_81730[7] = add_81612 == 32'h0000_0007 ? add_81728 : array_index_81722[7];
  assign array_update_81730[8] = add_81612 == 32'h0000_0008 ? add_81728 : array_index_81722[8];
  assign array_update_81730[9] = add_81612 == 32'h0000_0009 ? add_81728 : array_index_81722[9];
  assign add_81731 = add_81718 + 32'h0000_0001;
  assign array_update_81732[0] = add_81474 == 32'h0000_0000 ? array_update_81730 : array_update_81719[0];
  assign array_update_81732[1] = add_81474 == 32'h0000_0001 ? array_update_81730 : array_update_81719[1];
  assign array_update_81732[2] = add_81474 == 32'h0000_0002 ? array_update_81730 : array_update_81719[2];
  assign array_update_81732[3] = add_81474 == 32'h0000_0003 ? array_update_81730 : array_update_81719[3];
  assign array_update_81732[4] = add_81474 == 32'h0000_0004 ? array_update_81730 : array_update_81719[4];
  assign array_update_81732[5] = add_81474 == 32'h0000_0005 ? array_update_81730 : array_update_81719[5];
  assign array_update_81732[6] = add_81474 == 32'h0000_0006 ? array_update_81730 : array_update_81719[6];
  assign array_update_81732[7] = add_81474 == 32'h0000_0007 ? array_update_81730 : array_update_81719[7];
  assign array_update_81732[8] = add_81474 == 32'h0000_0008 ? array_update_81730 : array_update_81719[8];
  assign array_update_81732[9] = add_81474 == 32'h0000_0009 ? array_update_81730 : array_update_81719[9];
  assign array_index_81734 = array_update_72021[add_81731 > 32'h0000_0009 ? 4'h9 : add_81731[3:0]];
  assign array_index_81735 = array_update_81732[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_81739 = smul32b_32b_x_32b(array_index_81481[add_81731 > 32'h0000_0009 ? 4'h9 : add_81731[3:0]], array_index_81734[add_81612 > 32'h0000_0009 ? 4'h9 : add_81612[3:0]]);
  assign add_81741 = array_index_81735[add_81612 > 32'h0000_0009 ? 4'h9 : add_81612[3:0]] + smul_81739;
  assign array_update_81742[0] = add_81612 == 32'h0000_0000 ? add_81741 : array_index_81735[0];
  assign array_update_81742[1] = add_81612 == 32'h0000_0001 ? add_81741 : array_index_81735[1];
  assign array_update_81742[2] = add_81612 == 32'h0000_0002 ? add_81741 : array_index_81735[2];
  assign array_update_81742[3] = add_81612 == 32'h0000_0003 ? add_81741 : array_index_81735[3];
  assign array_update_81742[4] = add_81612 == 32'h0000_0004 ? add_81741 : array_index_81735[4];
  assign array_update_81742[5] = add_81612 == 32'h0000_0005 ? add_81741 : array_index_81735[5];
  assign array_update_81742[6] = add_81612 == 32'h0000_0006 ? add_81741 : array_index_81735[6];
  assign array_update_81742[7] = add_81612 == 32'h0000_0007 ? add_81741 : array_index_81735[7];
  assign array_update_81742[8] = add_81612 == 32'h0000_0008 ? add_81741 : array_index_81735[8];
  assign array_update_81742[9] = add_81612 == 32'h0000_0009 ? add_81741 : array_index_81735[9];
  assign array_update_81743[0] = add_81474 == 32'h0000_0000 ? array_update_81742 : array_update_81732[0];
  assign array_update_81743[1] = add_81474 == 32'h0000_0001 ? array_update_81742 : array_update_81732[1];
  assign array_update_81743[2] = add_81474 == 32'h0000_0002 ? array_update_81742 : array_update_81732[2];
  assign array_update_81743[3] = add_81474 == 32'h0000_0003 ? array_update_81742 : array_update_81732[3];
  assign array_update_81743[4] = add_81474 == 32'h0000_0004 ? array_update_81742 : array_update_81732[4];
  assign array_update_81743[5] = add_81474 == 32'h0000_0005 ? array_update_81742 : array_update_81732[5];
  assign array_update_81743[6] = add_81474 == 32'h0000_0006 ? array_update_81742 : array_update_81732[6];
  assign array_update_81743[7] = add_81474 == 32'h0000_0007 ? array_update_81742 : array_update_81732[7];
  assign array_update_81743[8] = add_81474 == 32'h0000_0008 ? array_update_81742 : array_update_81732[8];
  assign array_update_81743[9] = add_81474 == 32'h0000_0009 ? array_update_81742 : array_update_81732[9];
  assign array_index_81745 = array_update_81743[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign add_81747 = add_81612 + 32'h0000_0001;
  assign array_update_81748[0] = add_81747 == 32'h0000_0000 ? 32'h0000_0000 : array_index_81745[0];
  assign array_update_81748[1] = add_81747 == 32'h0000_0001 ? 32'h0000_0000 : array_index_81745[1];
  assign array_update_81748[2] = add_81747 == 32'h0000_0002 ? 32'h0000_0000 : array_index_81745[2];
  assign array_update_81748[3] = add_81747 == 32'h0000_0003 ? 32'h0000_0000 : array_index_81745[3];
  assign array_update_81748[4] = add_81747 == 32'h0000_0004 ? 32'h0000_0000 : array_index_81745[4];
  assign array_update_81748[5] = add_81747 == 32'h0000_0005 ? 32'h0000_0000 : array_index_81745[5];
  assign array_update_81748[6] = add_81747 == 32'h0000_0006 ? 32'h0000_0000 : array_index_81745[6];
  assign array_update_81748[7] = add_81747 == 32'h0000_0007 ? 32'h0000_0000 : array_index_81745[7];
  assign array_update_81748[8] = add_81747 == 32'h0000_0008 ? 32'h0000_0000 : array_index_81745[8];
  assign array_update_81748[9] = add_81747 == 32'h0000_0009 ? 32'h0000_0000 : array_index_81745[9];
  assign literal_81749 = 32'h0000_0000;
  assign array_update_81750[0] = add_81474 == 32'h0000_0000 ? array_update_81748 : array_update_81743[0];
  assign array_update_81750[1] = add_81474 == 32'h0000_0001 ? array_update_81748 : array_update_81743[1];
  assign array_update_81750[2] = add_81474 == 32'h0000_0002 ? array_update_81748 : array_update_81743[2];
  assign array_update_81750[3] = add_81474 == 32'h0000_0003 ? array_update_81748 : array_update_81743[3];
  assign array_update_81750[4] = add_81474 == 32'h0000_0004 ? array_update_81748 : array_update_81743[4];
  assign array_update_81750[5] = add_81474 == 32'h0000_0005 ? array_update_81748 : array_update_81743[5];
  assign array_update_81750[6] = add_81474 == 32'h0000_0006 ? array_update_81748 : array_update_81743[6];
  assign array_update_81750[7] = add_81474 == 32'h0000_0007 ? array_update_81748 : array_update_81743[7];
  assign array_update_81750[8] = add_81474 == 32'h0000_0008 ? array_update_81748 : array_update_81743[8];
  assign array_update_81750[9] = add_81474 == 32'h0000_0009 ? array_update_81748 : array_update_81743[9];
  assign array_index_81752 = array_update_72021[literal_81749 > 32'h0000_0009 ? 4'h9 : literal_81749[3:0]];
  assign array_index_81753 = array_update_81750[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_81757 = smul32b_32b_x_32b(array_index_81481[literal_81749 > 32'h0000_0009 ? 4'h9 : literal_81749[3:0]], array_index_81752[add_81747 > 32'h0000_0009 ? 4'h9 : add_81747[3:0]]);
  assign add_81759 = array_index_81753[add_81747 > 32'h0000_0009 ? 4'h9 : add_81747[3:0]] + smul_81757;
  assign array_update_81761[0] = add_81747 == 32'h0000_0000 ? add_81759 : array_index_81753[0];
  assign array_update_81761[1] = add_81747 == 32'h0000_0001 ? add_81759 : array_index_81753[1];
  assign array_update_81761[2] = add_81747 == 32'h0000_0002 ? add_81759 : array_index_81753[2];
  assign array_update_81761[3] = add_81747 == 32'h0000_0003 ? add_81759 : array_index_81753[3];
  assign array_update_81761[4] = add_81747 == 32'h0000_0004 ? add_81759 : array_index_81753[4];
  assign array_update_81761[5] = add_81747 == 32'h0000_0005 ? add_81759 : array_index_81753[5];
  assign array_update_81761[6] = add_81747 == 32'h0000_0006 ? add_81759 : array_index_81753[6];
  assign array_update_81761[7] = add_81747 == 32'h0000_0007 ? add_81759 : array_index_81753[7];
  assign array_update_81761[8] = add_81747 == 32'h0000_0008 ? add_81759 : array_index_81753[8];
  assign array_update_81761[9] = add_81747 == 32'h0000_0009 ? add_81759 : array_index_81753[9];
  assign add_81762 = literal_81749 + 32'h0000_0001;
  assign array_update_81763[0] = add_81474 == 32'h0000_0000 ? array_update_81761 : array_update_81750[0];
  assign array_update_81763[1] = add_81474 == 32'h0000_0001 ? array_update_81761 : array_update_81750[1];
  assign array_update_81763[2] = add_81474 == 32'h0000_0002 ? array_update_81761 : array_update_81750[2];
  assign array_update_81763[3] = add_81474 == 32'h0000_0003 ? array_update_81761 : array_update_81750[3];
  assign array_update_81763[4] = add_81474 == 32'h0000_0004 ? array_update_81761 : array_update_81750[4];
  assign array_update_81763[5] = add_81474 == 32'h0000_0005 ? array_update_81761 : array_update_81750[5];
  assign array_update_81763[6] = add_81474 == 32'h0000_0006 ? array_update_81761 : array_update_81750[6];
  assign array_update_81763[7] = add_81474 == 32'h0000_0007 ? array_update_81761 : array_update_81750[7];
  assign array_update_81763[8] = add_81474 == 32'h0000_0008 ? array_update_81761 : array_update_81750[8];
  assign array_update_81763[9] = add_81474 == 32'h0000_0009 ? array_update_81761 : array_update_81750[9];
  assign array_index_81765 = array_update_72021[add_81762 > 32'h0000_0009 ? 4'h9 : add_81762[3:0]];
  assign array_index_81766 = array_update_81763[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_81770 = smul32b_32b_x_32b(array_index_81481[add_81762 > 32'h0000_0009 ? 4'h9 : add_81762[3:0]], array_index_81765[add_81747 > 32'h0000_0009 ? 4'h9 : add_81747[3:0]]);
  assign add_81772 = array_index_81766[add_81747 > 32'h0000_0009 ? 4'h9 : add_81747[3:0]] + smul_81770;
  assign array_update_81774[0] = add_81747 == 32'h0000_0000 ? add_81772 : array_index_81766[0];
  assign array_update_81774[1] = add_81747 == 32'h0000_0001 ? add_81772 : array_index_81766[1];
  assign array_update_81774[2] = add_81747 == 32'h0000_0002 ? add_81772 : array_index_81766[2];
  assign array_update_81774[3] = add_81747 == 32'h0000_0003 ? add_81772 : array_index_81766[3];
  assign array_update_81774[4] = add_81747 == 32'h0000_0004 ? add_81772 : array_index_81766[4];
  assign array_update_81774[5] = add_81747 == 32'h0000_0005 ? add_81772 : array_index_81766[5];
  assign array_update_81774[6] = add_81747 == 32'h0000_0006 ? add_81772 : array_index_81766[6];
  assign array_update_81774[7] = add_81747 == 32'h0000_0007 ? add_81772 : array_index_81766[7];
  assign array_update_81774[8] = add_81747 == 32'h0000_0008 ? add_81772 : array_index_81766[8];
  assign array_update_81774[9] = add_81747 == 32'h0000_0009 ? add_81772 : array_index_81766[9];
  assign add_81775 = add_81762 + 32'h0000_0001;
  assign array_update_81776[0] = add_81474 == 32'h0000_0000 ? array_update_81774 : array_update_81763[0];
  assign array_update_81776[1] = add_81474 == 32'h0000_0001 ? array_update_81774 : array_update_81763[1];
  assign array_update_81776[2] = add_81474 == 32'h0000_0002 ? array_update_81774 : array_update_81763[2];
  assign array_update_81776[3] = add_81474 == 32'h0000_0003 ? array_update_81774 : array_update_81763[3];
  assign array_update_81776[4] = add_81474 == 32'h0000_0004 ? array_update_81774 : array_update_81763[4];
  assign array_update_81776[5] = add_81474 == 32'h0000_0005 ? array_update_81774 : array_update_81763[5];
  assign array_update_81776[6] = add_81474 == 32'h0000_0006 ? array_update_81774 : array_update_81763[6];
  assign array_update_81776[7] = add_81474 == 32'h0000_0007 ? array_update_81774 : array_update_81763[7];
  assign array_update_81776[8] = add_81474 == 32'h0000_0008 ? array_update_81774 : array_update_81763[8];
  assign array_update_81776[9] = add_81474 == 32'h0000_0009 ? array_update_81774 : array_update_81763[9];
  assign array_index_81778 = array_update_72021[add_81775 > 32'h0000_0009 ? 4'h9 : add_81775[3:0]];
  assign array_index_81779 = array_update_81776[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_81783 = smul32b_32b_x_32b(array_index_81481[add_81775 > 32'h0000_0009 ? 4'h9 : add_81775[3:0]], array_index_81778[add_81747 > 32'h0000_0009 ? 4'h9 : add_81747[3:0]]);
  assign add_81785 = array_index_81779[add_81747 > 32'h0000_0009 ? 4'h9 : add_81747[3:0]] + smul_81783;
  assign array_update_81787[0] = add_81747 == 32'h0000_0000 ? add_81785 : array_index_81779[0];
  assign array_update_81787[1] = add_81747 == 32'h0000_0001 ? add_81785 : array_index_81779[1];
  assign array_update_81787[2] = add_81747 == 32'h0000_0002 ? add_81785 : array_index_81779[2];
  assign array_update_81787[3] = add_81747 == 32'h0000_0003 ? add_81785 : array_index_81779[3];
  assign array_update_81787[4] = add_81747 == 32'h0000_0004 ? add_81785 : array_index_81779[4];
  assign array_update_81787[5] = add_81747 == 32'h0000_0005 ? add_81785 : array_index_81779[5];
  assign array_update_81787[6] = add_81747 == 32'h0000_0006 ? add_81785 : array_index_81779[6];
  assign array_update_81787[7] = add_81747 == 32'h0000_0007 ? add_81785 : array_index_81779[7];
  assign array_update_81787[8] = add_81747 == 32'h0000_0008 ? add_81785 : array_index_81779[8];
  assign array_update_81787[9] = add_81747 == 32'h0000_0009 ? add_81785 : array_index_81779[9];
  assign add_81788 = add_81775 + 32'h0000_0001;
  assign array_update_81789[0] = add_81474 == 32'h0000_0000 ? array_update_81787 : array_update_81776[0];
  assign array_update_81789[1] = add_81474 == 32'h0000_0001 ? array_update_81787 : array_update_81776[1];
  assign array_update_81789[2] = add_81474 == 32'h0000_0002 ? array_update_81787 : array_update_81776[2];
  assign array_update_81789[3] = add_81474 == 32'h0000_0003 ? array_update_81787 : array_update_81776[3];
  assign array_update_81789[4] = add_81474 == 32'h0000_0004 ? array_update_81787 : array_update_81776[4];
  assign array_update_81789[5] = add_81474 == 32'h0000_0005 ? array_update_81787 : array_update_81776[5];
  assign array_update_81789[6] = add_81474 == 32'h0000_0006 ? array_update_81787 : array_update_81776[6];
  assign array_update_81789[7] = add_81474 == 32'h0000_0007 ? array_update_81787 : array_update_81776[7];
  assign array_update_81789[8] = add_81474 == 32'h0000_0008 ? array_update_81787 : array_update_81776[8];
  assign array_update_81789[9] = add_81474 == 32'h0000_0009 ? array_update_81787 : array_update_81776[9];
  assign array_index_81791 = array_update_72021[add_81788 > 32'h0000_0009 ? 4'h9 : add_81788[3:0]];
  assign array_index_81792 = array_update_81789[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_81796 = smul32b_32b_x_32b(array_index_81481[add_81788 > 32'h0000_0009 ? 4'h9 : add_81788[3:0]], array_index_81791[add_81747 > 32'h0000_0009 ? 4'h9 : add_81747[3:0]]);
  assign add_81798 = array_index_81792[add_81747 > 32'h0000_0009 ? 4'h9 : add_81747[3:0]] + smul_81796;
  assign array_update_81800[0] = add_81747 == 32'h0000_0000 ? add_81798 : array_index_81792[0];
  assign array_update_81800[1] = add_81747 == 32'h0000_0001 ? add_81798 : array_index_81792[1];
  assign array_update_81800[2] = add_81747 == 32'h0000_0002 ? add_81798 : array_index_81792[2];
  assign array_update_81800[3] = add_81747 == 32'h0000_0003 ? add_81798 : array_index_81792[3];
  assign array_update_81800[4] = add_81747 == 32'h0000_0004 ? add_81798 : array_index_81792[4];
  assign array_update_81800[5] = add_81747 == 32'h0000_0005 ? add_81798 : array_index_81792[5];
  assign array_update_81800[6] = add_81747 == 32'h0000_0006 ? add_81798 : array_index_81792[6];
  assign array_update_81800[7] = add_81747 == 32'h0000_0007 ? add_81798 : array_index_81792[7];
  assign array_update_81800[8] = add_81747 == 32'h0000_0008 ? add_81798 : array_index_81792[8];
  assign array_update_81800[9] = add_81747 == 32'h0000_0009 ? add_81798 : array_index_81792[9];
  assign add_81801 = add_81788 + 32'h0000_0001;
  assign array_update_81802[0] = add_81474 == 32'h0000_0000 ? array_update_81800 : array_update_81789[0];
  assign array_update_81802[1] = add_81474 == 32'h0000_0001 ? array_update_81800 : array_update_81789[1];
  assign array_update_81802[2] = add_81474 == 32'h0000_0002 ? array_update_81800 : array_update_81789[2];
  assign array_update_81802[3] = add_81474 == 32'h0000_0003 ? array_update_81800 : array_update_81789[3];
  assign array_update_81802[4] = add_81474 == 32'h0000_0004 ? array_update_81800 : array_update_81789[4];
  assign array_update_81802[5] = add_81474 == 32'h0000_0005 ? array_update_81800 : array_update_81789[5];
  assign array_update_81802[6] = add_81474 == 32'h0000_0006 ? array_update_81800 : array_update_81789[6];
  assign array_update_81802[7] = add_81474 == 32'h0000_0007 ? array_update_81800 : array_update_81789[7];
  assign array_update_81802[8] = add_81474 == 32'h0000_0008 ? array_update_81800 : array_update_81789[8];
  assign array_update_81802[9] = add_81474 == 32'h0000_0009 ? array_update_81800 : array_update_81789[9];
  assign array_index_81804 = array_update_72021[add_81801 > 32'h0000_0009 ? 4'h9 : add_81801[3:0]];
  assign array_index_81805 = array_update_81802[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_81809 = smul32b_32b_x_32b(array_index_81481[add_81801 > 32'h0000_0009 ? 4'h9 : add_81801[3:0]], array_index_81804[add_81747 > 32'h0000_0009 ? 4'h9 : add_81747[3:0]]);
  assign add_81811 = array_index_81805[add_81747 > 32'h0000_0009 ? 4'h9 : add_81747[3:0]] + smul_81809;
  assign array_update_81813[0] = add_81747 == 32'h0000_0000 ? add_81811 : array_index_81805[0];
  assign array_update_81813[1] = add_81747 == 32'h0000_0001 ? add_81811 : array_index_81805[1];
  assign array_update_81813[2] = add_81747 == 32'h0000_0002 ? add_81811 : array_index_81805[2];
  assign array_update_81813[3] = add_81747 == 32'h0000_0003 ? add_81811 : array_index_81805[3];
  assign array_update_81813[4] = add_81747 == 32'h0000_0004 ? add_81811 : array_index_81805[4];
  assign array_update_81813[5] = add_81747 == 32'h0000_0005 ? add_81811 : array_index_81805[5];
  assign array_update_81813[6] = add_81747 == 32'h0000_0006 ? add_81811 : array_index_81805[6];
  assign array_update_81813[7] = add_81747 == 32'h0000_0007 ? add_81811 : array_index_81805[7];
  assign array_update_81813[8] = add_81747 == 32'h0000_0008 ? add_81811 : array_index_81805[8];
  assign array_update_81813[9] = add_81747 == 32'h0000_0009 ? add_81811 : array_index_81805[9];
  assign add_81814 = add_81801 + 32'h0000_0001;
  assign array_update_81815[0] = add_81474 == 32'h0000_0000 ? array_update_81813 : array_update_81802[0];
  assign array_update_81815[1] = add_81474 == 32'h0000_0001 ? array_update_81813 : array_update_81802[1];
  assign array_update_81815[2] = add_81474 == 32'h0000_0002 ? array_update_81813 : array_update_81802[2];
  assign array_update_81815[3] = add_81474 == 32'h0000_0003 ? array_update_81813 : array_update_81802[3];
  assign array_update_81815[4] = add_81474 == 32'h0000_0004 ? array_update_81813 : array_update_81802[4];
  assign array_update_81815[5] = add_81474 == 32'h0000_0005 ? array_update_81813 : array_update_81802[5];
  assign array_update_81815[6] = add_81474 == 32'h0000_0006 ? array_update_81813 : array_update_81802[6];
  assign array_update_81815[7] = add_81474 == 32'h0000_0007 ? array_update_81813 : array_update_81802[7];
  assign array_update_81815[8] = add_81474 == 32'h0000_0008 ? array_update_81813 : array_update_81802[8];
  assign array_update_81815[9] = add_81474 == 32'h0000_0009 ? array_update_81813 : array_update_81802[9];
  assign array_index_81817 = array_update_72021[add_81814 > 32'h0000_0009 ? 4'h9 : add_81814[3:0]];
  assign array_index_81818 = array_update_81815[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_81822 = smul32b_32b_x_32b(array_index_81481[add_81814 > 32'h0000_0009 ? 4'h9 : add_81814[3:0]], array_index_81817[add_81747 > 32'h0000_0009 ? 4'h9 : add_81747[3:0]]);
  assign add_81824 = array_index_81818[add_81747 > 32'h0000_0009 ? 4'h9 : add_81747[3:0]] + smul_81822;
  assign array_update_81826[0] = add_81747 == 32'h0000_0000 ? add_81824 : array_index_81818[0];
  assign array_update_81826[1] = add_81747 == 32'h0000_0001 ? add_81824 : array_index_81818[1];
  assign array_update_81826[2] = add_81747 == 32'h0000_0002 ? add_81824 : array_index_81818[2];
  assign array_update_81826[3] = add_81747 == 32'h0000_0003 ? add_81824 : array_index_81818[3];
  assign array_update_81826[4] = add_81747 == 32'h0000_0004 ? add_81824 : array_index_81818[4];
  assign array_update_81826[5] = add_81747 == 32'h0000_0005 ? add_81824 : array_index_81818[5];
  assign array_update_81826[6] = add_81747 == 32'h0000_0006 ? add_81824 : array_index_81818[6];
  assign array_update_81826[7] = add_81747 == 32'h0000_0007 ? add_81824 : array_index_81818[7];
  assign array_update_81826[8] = add_81747 == 32'h0000_0008 ? add_81824 : array_index_81818[8];
  assign array_update_81826[9] = add_81747 == 32'h0000_0009 ? add_81824 : array_index_81818[9];
  assign add_81827 = add_81814 + 32'h0000_0001;
  assign array_update_81828[0] = add_81474 == 32'h0000_0000 ? array_update_81826 : array_update_81815[0];
  assign array_update_81828[1] = add_81474 == 32'h0000_0001 ? array_update_81826 : array_update_81815[1];
  assign array_update_81828[2] = add_81474 == 32'h0000_0002 ? array_update_81826 : array_update_81815[2];
  assign array_update_81828[3] = add_81474 == 32'h0000_0003 ? array_update_81826 : array_update_81815[3];
  assign array_update_81828[4] = add_81474 == 32'h0000_0004 ? array_update_81826 : array_update_81815[4];
  assign array_update_81828[5] = add_81474 == 32'h0000_0005 ? array_update_81826 : array_update_81815[5];
  assign array_update_81828[6] = add_81474 == 32'h0000_0006 ? array_update_81826 : array_update_81815[6];
  assign array_update_81828[7] = add_81474 == 32'h0000_0007 ? array_update_81826 : array_update_81815[7];
  assign array_update_81828[8] = add_81474 == 32'h0000_0008 ? array_update_81826 : array_update_81815[8];
  assign array_update_81828[9] = add_81474 == 32'h0000_0009 ? array_update_81826 : array_update_81815[9];
  assign array_index_81830 = array_update_72021[add_81827 > 32'h0000_0009 ? 4'h9 : add_81827[3:0]];
  assign array_index_81831 = array_update_81828[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_81835 = smul32b_32b_x_32b(array_index_81481[add_81827 > 32'h0000_0009 ? 4'h9 : add_81827[3:0]], array_index_81830[add_81747 > 32'h0000_0009 ? 4'h9 : add_81747[3:0]]);
  assign add_81837 = array_index_81831[add_81747 > 32'h0000_0009 ? 4'h9 : add_81747[3:0]] + smul_81835;
  assign array_update_81839[0] = add_81747 == 32'h0000_0000 ? add_81837 : array_index_81831[0];
  assign array_update_81839[1] = add_81747 == 32'h0000_0001 ? add_81837 : array_index_81831[1];
  assign array_update_81839[2] = add_81747 == 32'h0000_0002 ? add_81837 : array_index_81831[2];
  assign array_update_81839[3] = add_81747 == 32'h0000_0003 ? add_81837 : array_index_81831[3];
  assign array_update_81839[4] = add_81747 == 32'h0000_0004 ? add_81837 : array_index_81831[4];
  assign array_update_81839[5] = add_81747 == 32'h0000_0005 ? add_81837 : array_index_81831[5];
  assign array_update_81839[6] = add_81747 == 32'h0000_0006 ? add_81837 : array_index_81831[6];
  assign array_update_81839[7] = add_81747 == 32'h0000_0007 ? add_81837 : array_index_81831[7];
  assign array_update_81839[8] = add_81747 == 32'h0000_0008 ? add_81837 : array_index_81831[8];
  assign array_update_81839[9] = add_81747 == 32'h0000_0009 ? add_81837 : array_index_81831[9];
  assign add_81840 = add_81827 + 32'h0000_0001;
  assign array_update_81841[0] = add_81474 == 32'h0000_0000 ? array_update_81839 : array_update_81828[0];
  assign array_update_81841[1] = add_81474 == 32'h0000_0001 ? array_update_81839 : array_update_81828[1];
  assign array_update_81841[2] = add_81474 == 32'h0000_0002 ? array_update_81839 : array_update_81828[2];
  assign array_update_81841[3] = add_81474 == 32'h0000_0003 ? array_update_81839 : array_update_81828[3];
  assign array_update_81841[4] = add_81474 == 32'h0000_0004 ? array_update_81839 : array_update_81828[4];
  assign array_update_81841[5] = add_81474 == 32'h0000_0005 ? array_update_81839 : array_update_81828[5];
  assign array_update_81841[6] = add_81474 == 32'h0000_0006 ? array_update_81839 : array_update_81828[6];
  assign array_update_81841[7] = add_81474 == 32'h0000_0007 ? array_update_81839 : array_update_81828[7];
  assign array_update_81841[8] = add_81474 == 32'h0000_0008 ? array_update_81839 : array_update_81828[8];
  assign array_update_81841[9] = add_81474 == 32'h0000_0009 ? array_update_81839 : array_update_81828[9];
  assign array_index_81843 = array_update_72021[add_81840 > 32'h0000_0009 ? 4'h9 : add_81840[3:0]];
  assign array_index_81844 = array_update_81841[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_81848 = smul32b_32b_x_32b(array_index_81481[add_81840 > 32'h0000_0009 ? 4'h9 : add_81840[3:0]], array_index_81843[add_81747 > 32'h0000_0009 ? 4'h9 : add_81747[3:0]]);
  assign add_81850 = array_index_81844[add_81747 > 32'h0000_0009 ? 4'h9 : add_81747[3:0]] + smul_81848;
  assign array_update_81852[0] = add_81747 == 32'h0000_0000 ? add_81850 : array_index_81844[0];
  assign array_update_81852[1] = add_81747 == 32'h0000_0001 ? add_81850 : array_index_81844[1];
  assign array_update_81852[2] = add_81747 == 32'h0000_0002 ? add_81850 : array_index_81844[2];
  assign array_update_81852[3] = add_81747 == 32'h0000_0003 ? add_81850 : array_index_81844[3];
  assign array_update_81852[4] = add_81747 == 32'h0000_0004 ? add_81850 : array_index_81844[4];
  assign array_update_81852[5] = add_81747 == 32'h0000_0005 ? add_81850 : array_index_81844[5];
  assign array_update_81852[6] = add_81747 == 32'h0000_0006 ? add_81850 : array_index_81844[6];
  assign array_update_81852[7] = add_81747 == 32'h0000_0007 ? add_81850 : array_index_81844[7];
  assign array_update_81852[8] = add_81747 == 32'h0000_0008 ? add_81850 : array_index_81844[8];
  assign array_update_81852[9] = add_81747 == 32'h0000_0009 ? add_81850 : array_index_81844[9];
  assign add_81853 = add_81840 + 32'h0000_0001;
  assign array_update_81854[0] = add_81474 == 32'h0000_0000 ? array_update_81852 : array_update_81841[0];
  assign array_update_81854[1] = add_81474 == 32'h0000_0001 ? array_update_81852 : array_update_81841[1];
  assign array_update_81854[2] = add_81474 == 32'h0000_0002 ? array_update_81852 : array_update_81841[2];
  assign array_update_81854[3] = add_81474 == 32'h0000_0003 ? array_update_81852 : array_update_81841[3];
  assign array_update_81854[4] = add_81474 == 32'h0000_0004 ? array_update_81852 : array_update_81841[4];
  assign array_update_81854[5] = add_81474 == 32'h0000_0005 ? array_update_81852 : array_update_81841[5];
  assign array_update_81854[6] = add_81474 == 32'h0000_0006 ? array_update_81852 : array_update_81841[6];
  assign array_update_81854[7] = add_81474 == 32'h0000_0007 ? array_update_81852 : array_update_81841[7];
  assign array_update_81854[8] = add_81474 == 32'h0000_0008 ? array_update_81852 : array_update_81841[8];
  assign array_update_81854[9] = add_81474 == 32'h0000_0009 ? array_update_81852 : array_update_81841[9];
  assign array_index_81856 = array_update_72021[add_81853 > 32'h0000_0009 ? 4'h9 : add_81853[3:0]];
  assign array_index_81857 = array_update_81854[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_81861 = smul32b_32b_x_32b(array_index_81481[add_81853 > 32'h0000_0009 ? 4'h9 : add_81853[3:0]], array_index_81856[add_81747 > 32'h0000_0009 ? 4'h9 : add_81747[3:0]]);
  assign add_81863 = array_index_81857[add_81747 > 32'h0000_0009 ? 4'h9 : add_81747[3:0]] + smul_81861;
  assign array_update_81865[0] = add_81747 == 32'h0000_0000 ? add_81863 : array_index_81857[0];
  assign array_update_81865[1] = add_81747 == 32'h0000_0001 ? add_81863 : array_index_81857[1];
  assign array_update_81865[2] = add_81747 == 32'h0000_0002 ? add_81863 : array_index_81857[2];
  assign array_update_81865[3] = add_81747 == 32'h0000_0003 ? add_81863 : array_index_81857[3];
  assign array_update_81865[4] = add_81747 == 32'h0000_0004 ? add_81863 : array_index_81857[4];
  assign array_update_81865[5] = add_81747 == 32'h0000_0005 ? add_81863 : array_index_81857[5];
  assign array_update_81865[6] = add_81747 == 32'h0000_0006 ? add_81863 : array_index_81857[6];
  assign array_update_81865[7] = add_81747 == 32'h0000_0007 ? add_81863 : array_index_81857[7];
  assign array_update_81865[8] = add_81747 == 32'h0000_0008 ? add_81863 : array_index_81857[8];
  assign array_update_81865[9] = add_81747 == 32'h0000_0009 ? add_81863 : array_index_81857[9];
  assign add_81866 = add_81853 + 32'h0000_0001;
  assign array_update_81867[0] = add_81474 == 32'h0000_0000 ? array_update_81865 : array_update_81854[0];
  assign array_update_81867[1] = add_81474 == 32'h0000_0001 ? array_update_81865 : array_update_81854[1];
  assign array_update_81867[2] = add_81474 == 32'h0000_0002 ? array_update_81865 : array_update_81854[2];
  assign array_update_81867[3] = add_81474 == 32'h0000_0003 ? array_update_81865 : array_update_81854[3];
  assign array_update_81867[4] = add_81474 == 32'h0000_0004 ? array_update_81865 : array_update_81854[4];
  assign array_update_81867[5] = add_81474 == 32'h0000_0005 ? array_update_81865 : array_update_81854[5];
  assign array_update_81867[6] = add_81474 == 32'h0000_0006 ? array_update_81865 : array_update_81854[6];
  assign array_update_81867[7] = add_81474 == 32'h0000_0007 ? array_update_81865 : array_update_81854[7];
  assign array_update_81867[8] = add_81474 == 32'h0000_0008 ? array_update_81865 : array_update_81854[8];
  assign array_update_81867[9] = add_81474 == 32'h0000_0009 ? array_update_81865 : array_update_81854[9];
  assign array_index_81869 = array_update_72021[add_81866 > 32'h0000_0009 ? 4'h9 : add_81866[3:0]];
  assign array_index_81870 = array_update_81867[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_81874 = smul32b_32b_x_32b(array_index_81481[add_81866 > 32'h0000_0009 ? 4'h9 : add_81866[3:0]], array_index_81869[add_81747 > 32'h0000_0009 ? 4'h9 : add_81747[3:0]]);
  assign add_81876 = array_index_81870[add_81747 > 32'h0000_0009 ? 4'h9 : add_81747[3:0]] + smul_81874;
  assign array_update_81877[0] = add_81747 == 32'h0000_0000 ? add_81876 : array_index_81870[0];
  assign array_update_81877[1] = add_81747 == 32'h0000_0001 ? add_81876 : array_index_81870[1];
  assign array_update_81877[2] = add_81747 == 32'h0000_0002 ? add_81876 : array_index_81870[2];
  assign array_update_81877[3] = add_81747 == 32'h0000_0003 ? add_81876 : array_index_81870[3];
  assign array_update_81877[4] = add_81747 == 32'h0000_0004 ? add_81876 : array_index_81870[4];
  assign array_update_81877[5] = add_81747 == 32'h0000_0005 ? add_81876 : array_index_81870[5];
  assign array_update_81877[6] = add_81747 == 32'h0000_0006 ? add_81876 : array_index_81870[6];
  assign array_update_81877[7] = add_81747 == 32'h0000_0007 ? add_81876 : array_index_81870[7];
  assign array_update_81877[8] = add_81747 == 32'h0000_0008 ? add_81876 : array_index_81870[8];
  assign array_update_81877[9] = add_81747 == 32'h0000_0009 ? add_81876 : array_index_81870[9];
  assign array_update_81878[0] = add_81474 == 32'h0000_0000 ? array_update_81877 : array_update_81867[0];
  assign array_update_81878[1] = add_81474 == 32'h0000_0001 ? array_update_81877 : array_update_81867[1];
  assign array_update_81878[2] = add_81474 == 32'h0000_0002 ? array_update_81877 : array_update_81867[2];
  assign array_update_81878[3] = add_81474 == 32'h0000_0003 ? array_update_81877 : array_update_81867[3];
  assign array_update_81878[4] = add_81474 == 32'h0000_0004 ? array_update_81877 : array_update_81867[4];
  assign array_update_81878[5] = add_81474 == 32'h0000_0005 ? array_update_81877 : array_update_81867[5];
  assign array_update_81878[6] = add_81474 == 32'h0000_0006 ? array_update_81877 : array_update_81867[6];
  assign array_update_81878[7] = add_81474 == 32'h0000_0007 ? array_update_81877 : array_update_81867[7];
  assign array_update_81878[8] = add_81474 == 32'h0000_0008 ? array_update_81877 : array_update_81867[8];
  assign array_update_81878[9] = add_81474 == 32'h0000_0009 ? array_update_81877 : array_update_81867[9];
  assign array_index_81880 = array_update_81878[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign add_81882 = add_81747 + 32'h0000_0001;
  assign array_update_81883[0] = add_81882 == 32'h0000_0000 ? 32'h0000_0000 : array_index_81880[0];
  assign array_update_81883[1] = add_81882 == 32'h0000_0001 ? 32'h0000_0000 : array_index_81880[1];
  assign array_update_81883[2] = add_81882 == 32'h0000_0002 ? 32'h0000_0000 : array_index_81880[2];
  assign array_update_81883[3] = add_81882 == 32'h0000_0003 ? 32'h0000_0000 : array_index_81880[3];
  assign array_update_81883[4] = add_81882 == 32'h0000_0004 ? 32'h0000_0000 : array_index_81880[4];
  assign array_update_81883[5] = add_81882 == 32'h0000_0005 ? 32'h0000_0000 : array_index_81880[5];
  assign array_update_81883[6] = add_81882 == 32'h0000_0006 ? 32'h0000_0000 : array_index_81880[6];
  assign array_update_81883[7] = add_81882 == 32'h0000_0007 ? 32'h0000_0000 : array_index_81880[7];
  assign array_update_81883[8] = add_81882 == 32'h0000_0008 ? 32'h0000_0000 : array_index_81880[8];
  assign array_update_81883[9] = add_81882 == 32'h0000_0009 ? 32'h0000_0000 : array_index_81880[9];
  assign literal_81884 = 32'h0000_0000;
  assign array_update_81885[0] = add_81474 == 32'h0000_0000 ? array_update_81883 : array_update_81878[0];
  assign array_update_81885[1] = add_81474 == 32'h0000_0001 ? array_update_81883 : array_update_81878[1];
  assign array_update_81885[2] = add_81474 == 32'h0000_0002 ? array_update_81883 : array_update_81878[2];
  assign array_update_81885[3] = add_81474 == 32'h0000_0003 ? array_update_81883 : array_update_81878[3];
  assign array_update_81885[4] = add_81474 == 32'h0000_0004 ? array_update_81883 : array_update_81878[4];
  assign array_update_81885[5] = add_81474 == 32'h0000_0005 ? array_update_81883 : array_update_81878[5];
  assign array_update_81885[6] = add_81474 == 32'h0000_0006 ? array_update_81883 : array_update_81878[6];
  assign array_update_81885[7] = add_81474 == 32'h0000_0007 ? array_update_81883 : array_update_81878[7];
  assign array_update_81885[8] = add_81474 == 32'h0000_0008 ? array_update_81883 : array_update_81878[8];
  assign array_update_81885[9] = add_81474 == 32'h0000_0009 ? array_update_81883 : array_update_81878[9];
  assign array_index_81887 = array_update_72021[literal_81884 > 32'h0000_0009 ? 4'h9 : literal_81884[3:0]];
  assign array_index_81888 = array_update_81885[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_81892 = smul32b_32b_x_32b(array_index_81481[literal_81884 > 32'h0000_0009 ? 4'h9 : literal_81884[3:0]], array_index_81887[add_81882 > 32'h0000_0009 ? 4'h9 : add_81882[3:0]]);
  assign add_81894 = array_index_81888[add_81882 > 32'h0000_0009 ? 4'h9 : add_81882[3:0]] + smul_81892;
  assign array_update_81896[0] = add_81882 == 32'h0000_0000 ? add_81894 : array_index_81888[0];
  assign array_update_81896[1] = add_81882 == 32'h0000_0001 ? add_81894 : array_index_81888[1];
  assign array_update_81896[2] = add_81882 == 32'h0000_0002 ? add_81894 : array_index_81888[2];
  assign array_update_81896[3] = add_81882 == 32'h0000_0003 ? add_81894 : array_index_81888[3];
  assign array_update_81896[4] = add_81882 == 32'h0000_0004 ? add_81894 : array_index_81888[4];
  assign array_update_81896[5] = add_81882 == 32'h0000_0005 ? add_81894 : array_index_81888[5];
  assign array_update_81896[6] = add_81882 == 32'h0000_0006 ? add_81894 : array_index_81888[6];
  assign array_update_81896[7] = add_81882 == 32'h0000_0007 ? add_81894 : array_index_81888[7];
  assign array_update_81896[8] = add_81882 == 32'h0000_0008 ? add_81894 : array_index_81888[8];
  assign array_update_81896[9] = add_81882 == 32'h0000_0009 ? add_81894 : array_index_81888[9];
  assign add_81897 = literal_81884 + 32'h0000_0001;
  assign array_update_81898[0] = add_81474 == 32'h0000_0000 ? array_update_81896 : array_update_81885[0];
  assign array_update_81898[1] = add_81474 == 32'h0000_0001 ? array_update_81896 : array_update_81885[1];
  assign array_update_81898[2] = add_81474 == 32'h0000_0002 ? array_update_81896 : array_update_81885[2];
  assign array_update_81898[3] = add_81474 == 32'h0000_0003 ? array_update_81896 : array_update_81885[3];
  assign array_update_81898[4] = add_81474 == 32'h0000_0004 ? array_update_81896 : array_update_81885[4];
  assign array_update_81898[5] = add_81474 == 32'h0000_0005 ? array_update_81896 : array_update_81885[5];
  assign array_update_81898[6] = add_81474 == 32'h0000_0006 ? array_update_81896 : array_update_81885[6];
  assign array_update_81898[7] = add_81474 == 32'h0000_0007 ? array_update_81896 : array_update_81885[7];
  assign array_update_81898[8] = add_81474 == 32'h0000_0008 ? array_update_81896 : array_update_81885[8];
  assign array_update_81898[9] = add_81474 == 32'h0000_0009 ? array_update_81896 : array_update_81885[9];
  assign array_index_81900 = array_update_72021[add_81897 > 32'h0000_0009 ? 4'h9 : add_81897[3:0]];
  assign array_index_81901 = array_update_81898[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_81905 = smul32b_32b_x_32b(array_index_81481[add_81897 > 32'h0000_0009 ? 4'h9 : add_81897[3:0]], array_index_81900[add_81882 > 32'h0000_0009 ? 4'h9 : add_81882[3:0]]);
  assign add_81907 = array_index_81901[add_81882 > 32'h0000_0009 ? 4'h9 : add_81882[3:0]] + smul_81905;
  assign array_update_81909[0] = add_81882 == 32'h0000_0000 ? add_81907 : array_index_81901[0];
  assign array_update_81909[1] = add_81882 == 32'h0000_0001 ? add_81907 : array_index_81901[1];
  assign array_update_81909[2] = add_81882 == 32'h0000_0002 ? add_81907 : array_index_81901[2];
  assign array_update_81909[3] = add_81882 == 32'h0000_0003 ? add_81907 : array_index_81901[3];
  assign array_update_81909[4] = add_81882 == 32'h0000_0004 ? add_81907 : array_index_81901[4];
  assign array_update_81909[5] = add_81882 == 32'h0000_0005 ? add_81907 : array_index_81901[5];
  assign array_update_81909[6] = add_81882 == 32'h0000_0006 ? add_81907 : array_index_81901[6];
  assign array_update_81909[7] = add_81882 == 32'h0000_0007 ? add_81907 : array_index_81901[7];
  assign array_update_81909[8] = add_81882 == 32'h0000_0008 ? add_81907 : array_index_81901[8];
  assign array_update_81909[9] = add_81882 == 32'h0000_0009 ? add_81907 : array_index_81901[9];
  assign add_81910 = add_81897 + 32'h0000_0001;
  assign array_update_81911[0] = add_81474 == 32'h0000_0000 ? array_update_81909 : array_update_81898[0];
  assign array_update_81911[1] = add_81474 == 32'h0000_0001 ? array_update_81909 : array_update_81898[1];
  assign array_update_81911[2] = add_81474 == 32'h0000_0002 ? array_update_81909 : array_update_81898[2];
  assign array_update_81911[3] = add_81474 == 32'h0000_0003 ? array_update_81909 : array_update_81898[3];
  assign array_update_81911[4] = add_81474 == 32'h0000_0004 ? array_update_81909 : array_update_81898[4];
  assign array_update_81911[5] = add_81474 == 32'h0000_0005 ? array_update_81909 : array_update_81898[5];
  assign array_update_81911[6] = add_81474 == 32'h0000_0006 ? array_update_81909 : array_update_81898[6];
  assign array_update_81911[7] = add_81474 == 32'h0000_0007 ? array_update_81909 : array_update_81898[7];
  assign array_update_81911[8] = add_81474 == 32'h0000_0008 ? array_update_81909 : array_update_81898[8];
  assign array_update_81911[9] = add_81474 == 32'h0000_0009 ? array_update_81909 : array_update_81898[9];
  assign array_index_81913 = array_update_72021[add_81910 > 32'h0000_0009 ? 4'h9 : add_81910[3:0]];
  assign array_index_81914 = array_update_81911[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_81918 = smul32b_32b_x_32b(array_index_81481[add_81910 > 32'h0000_0009 ? 4'h9 : add_81910[3:0]], array_index_81913[add_81882 > 32'h0000_0009 ? 4'h9 : add_81882[3:0]]);
  assign add_81920 = array_index_81914[add_81882 > 32'h0000_0009 ? 4'h9 : add_81882[3:0]] + smul_81918;
  assign array_update_81922[0] = add_81882 == 32'h0000_0000 ? add_81920 : array_index_81914[0];
  assign array_update_81922[1] = add_81882 == 32'h0000_0001 ? add_81920 : array_index_81914[1];
  assign array_update_81922[2] = add_81882 == 32'h0000_0002 ? add_81920 : array_index_81914[2];
  assign array_update_81922[3] = add_81882 == 32'h0000_0003 ? add_81920 : array_index_81914[3];
  assign array_update_81922[4] = add_81882 == 32'h0000_0004 ? add_81920 : array_index_81914[4];
  assign array_update_81922[5] = add_81882 == 32'h0000_0005 ? add_81920 : array_index_81914[5];
  assign array_update_81922[6] = add_81882 == 32'h0000_0006 ? add_81920 : array_index_81914[6];
  assign array_update_81922[7] = add_81882 == 32'h0000_0007 ? add_81920 : array_index_81914[7];
  assign array_update_81922[8] = add_81882 == 32'h0000_0008 ? add_81920 : array_index_81914[8];
  assign array_update_81922[9] = add_81882 == 32'h0000_0009 ? add_81920 : array_index_81914[9];
  assign add_81923 = add_81910 + 32'h0000_0001;
  assign array_update_81924[0] = add_81474 == 32'h0000_0000 ? array_update_81922 : array_update_81911[0];
  assign array_update_81924[1] = add_81474 == 32'h0000_0001 ? array_update_81922 : array_update_81911[1];
  assign array_update_81924[2] = add_81474 == 32'h0000_0002 ? array_update_81922 : array_update_81911[2];
  assign array_update_81924[3] = add_81474 == 32'h0000_0003 ? array_update_81922 : array_update_81911[3];
  assign array_update_81924[4] = add_81474 == 32'h0000_0004 ? array_update_81922 : array_update_81911[4];
  assign array_update_81924[5] = add_81474 == 32'h0000_0005 ? array_update_81922 : array_update_81911[5];
  assign array_update_81924[6] = add_81474 == 32'h0000_0006 ? array_update_81922 : array_update_81911[6];
  assign array_update_81924[7] = add_81474 == 32'h0000_0007 ? array_update_81922 : array_update_81911[7];
  assign array_update_81924[8] = add_81474 == 32'h0000_0008 ? array_update_81922 : array_update_81911[8];
  assign array_update_81924[9] = add_81474 == 32'h0000_0009 ? array_update_81922 : array_update_81911[9];
  assign array_index_81926 = array_update_72021[add_81923 > 32'h0000_0009 ? 4'h9 : add_81923[3:0]];
  assign array_index_81927 = array_update_81924[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_81931 = smul32b_32b_x_32b(array_index_81481[add_81923 > 32'h0000_0009 ? 4'h9 : add_81923[3:0]], array_index_81926[add_81882 > 32'h0000_0009 ? 4'h9 : add_81882[3:0]]);
  assign add_81933 = array_index_81927[add_81882 > 32'h0000_0009 ? 4'h9 : add_81882[3:0]] + smul_81931;
  assign array_update_81935[0] = add_81882 == 32'h0000_0000 ? add_81933 : array_index_81927[0];
  assign array_update_81935[1] = add_81882 == 32'h0000_0001 ? add_81933 : array_index_81927[1];
  assign array_update_81935[2] = add_81882 == 32'h0000_0002 ? add_81933 : array_index_81927[2];
  assign array_update_81935[3] = add_81882 == 32'h0000_0003 ? add_81933 : array_index_81927[3];
  assign array_update_81935[4] = add_81882 == 32'h0000_0004 ? add_81933 : array_index_81927[4];
  assign array_update_81935[5] = add_81882 == 32'h0000_0005 ? add_81933 : array_index_81927[5];
  assign array_update_81935[6] = add_81882 == 32'h0000_0006 ? add_81933 : array_index_81927[6];
  assign array_update_81935[7] = add_81882 == 32'h0000_0007 ? add_81933 : array_index_81927[7];
  assign array_update_81935[8] = add_81882 == 32'h0000_0008 ? add_81933 : array_index_81927[8];
  assign array_update_81935[9] = add_81882 == 32'h0000_0009 ? add_81933 : array_index_81927[9];
  assign add_81936 = add_81923 + 32'h0000_0001;
  assign array_update_81937[0] = add_81474 == 32'h0000_0000 ? array_update_81935 : array_update_81924[0];
  assign array_update_81937[1] = add_81474 == 32'h0000_0001 ? array_update_81935 : array_update_81924[1];
  assign array_update_81937[2] = add_81474 == 32'h0000_0002 ? array_update_81935 : array_update_81924[2];
  assign array_update_81937[3] = add_81474 == 32'h0000_0003 ? array_update_81935 : array_update_81924[3];
  assign array_update_81937[4] = add_81474 == 32'h0000_0004 ? array_update_81935 : array_update_81924[4];
  assign array_update_81937[5] = add_81474 == 32'h0000_0005 ? array_update_81935 : array_update_81924[5];
  assign array_update_81937[6] = add_81474 == 32'h0000_0006 ? array_update_81935 : array_update_81924[6];
  assign array_update_81937[7] = add_81474 == 32'h0000_0007 ? array_update_81935 : array_update_81924[7];
  assign array_update_81937[8] = add_81474 == 32'h0000_0008 ? array_update_81935 : array_update_81924[8];
  assign array_update_81937[9] = add_81474 == 32'h0000_0009 ? array_update_81935 : array_update_81924[9];
  assign array_index_81939 = array_update_72021[add_81936 > 32'h0000_0009 ? 4'h9 : add_81936[3:0]];
  assign array_index_81940 = array_update_81937[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_81944 = smul32b_32b_x_32b(array_index_81481[add_81936 > 32'h0000_0009 ? 4'h9 : add_81936[3:0]], array_index_81939[add_81882 > 32'h0000_0009 ? 4'h9 : add_81882[3:0]]);
  assign add_81946 = array_index_81940[add_81882 > 32'h0000_0009 ? 4'h9 : add_81882[3:0]] + smul_81944;
  assign array_update_81948[0] = add_81882 == 32'h0000_0000 ? add_81946 : array_index_81940[0];
  assign array_update_81948[1] = add_81882 == 32'h0000_0001 ? add_81946 : array_index_81940[1];
  assign array_update_81948[2] = add_81882 == 32'h0000_0002 ? add_81946 : array_index_81940[2];
  assign array_update_81948[3] = add_81882 == 32'h0000_0003 ? add_81946 : array_index_81940[3];
  assign array_update_81948[4] = add_81882 == 32'h0000_0004 ? add_81946 : array_index_81940[4];
  assign array_update_81948[5] = add_81882 == 32'h0000_0005 ? add_81946 : array_index_81940[5];
  assign array_update_81948[6] = add_81882 == 32'h0000_0006 ? add_81946 : array_index_81940[6];
  assign array_update_81948[7] = add_81882 == 32'h0000_0007 ? add_81946 : array_index_81940[7];
  assign array_update_81948[8] = add_81882 == 32'h0000_0008 ? add_81946 : array_index_81940[8];
  assign array_update_81948[9] = add_81882 == 32'h0000_0009 ? add_81946 : array_index_81940[9];
  assign add_81949 = add_81936 + 32'h0000_0001;
  assign array_update_81950[0] = add_81474 == 32'h0000_0000 ? array_update_81948 : array_update_81937[0];
  assign array_update_81950[1] = add_81474 == 32'h0000_0001 ? array_update_81948 : array_update_81937[1];
  assign array_update_81950[2] = add_81474 == 32'h0000_0002 ? array_update_81948 : array_update_81937[2];
  assign array_update_81950[3] = add_81474 == 32'h0000_0003 ? array_update_81948 : array_update_81937[3];
  assign array_update_81950[4] = add_81474 == 32'h0000_0004 ? array_update_81948 : array_update_81937[4];
  assign array_update_81950[5] = add_81474 == 32'h0000_0005 ? array_update_81948 : array_update_81937[5];
  assign array_update_81950[6] = add_81474 == 32'h0000_0006 ? array_update_81948 : array_update_81937[6];
  assign array_update_81950[7] = add_81474 == 32'h0000_0007 ? array_update_81948 : array_update_81937[7];
  assign array_update_81950[8] = add_81474 == 32'h0000_0008 ? array_update_81948 : array_update_81937[8];
  assign array_update_81950[9] = add_81474 == 32'h0000_0009 ? array_update_81948 : array_update_81937[9];
  assign array_index_81952 = array_update_72021[add_81949 > 32'h0000_0009 ? 4'h9 : add_81949[3:0]];
  assign array_index_81953 = array_update_81950[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_81957 = smul32b_32b_x_32b(array_index_81481[add_81949 > 32'h0000_0009 ? 4'h9 : add_81949[3:0]], array_index_81952[add_81882 > 32'h0000_0009 ? 4'h9 : add_81882[3:0]]);
  assign add_81959 = array_index_81953[add_81882 > 32'h0000_0009 ? 4'h9 : add_81882[3:0]] + smul_81957;
  assign array_update_81961[0] = add_81882 == 32'h0000_0000 ? add_81959 : array_index_81953[0];
  assign array_update_81961[1] = add_81882 == 32'h0000_0001 ? add_81959 : array_index_81953[1];
  assign array_update_81961[2] = add_81882 == 32'h0000_0002 ? add_81959 : array_index_81953[2];
  assign array_update_81961[3] = add_81882 == 32'h0000_0003 ? add_81959 : array_index_81953[3];
  assign array_update_81961[4] = add_81882 == 32'h0000_0004 ? add_81959 : array_index_81953[4];
  assign array_update_81961[5] = add_81882 == 32'h0000_0005 ? add_81959 : array_index_81953[5];
  assign array_update_81961[6] = add_81882 == 32'h0000_0006 ? add_81959 : array_index_81953[6];
  assign array_update_81961[7] = add_81882 == 32'h0000_0007 ? add_81959 : array_index_81953[7];
  assign array_update_81961[8] = add_81882 == 32'h0000_0008 ? add_81959 : array_index_81953[8];
  assign array_update_81961[9] = add_81882 == 32'h0000_0009 ? add_81959 : array_index_81953[9];
  assign add_81962 = add_81949 + 32'h0000_0001;
  assign array_update_81963[0] = add_81474 == 32'h0000_0000 ? array_update_81961 : array_update_81950[0];
  assign array_update_81963[1] = add_81474 == 32'h0000_0001 ? array_update_81961 : array_update_81950[1];
  assign array_update_81963[2] = add_81474 == 32'h0000_0002 ? array_update_81961 : array_update_81950[2];
  assign array_update_81963[3] = add_81474 == 32'h0000_0003 ? array_update_81961 : array_update_81950[3];
  assign array_update_81963[4] = add_81474 == 32'h0000_0004 ? array_update_81961 : array_update_81950[4];
  assign array_update_81963[5] = add_81474 == 32'h0000_0005 ? array_update_81961 : array_update_81950[5];
  assign array_update_81963[6] = add_81474 == 32'h0000_0006 ? array_update_81961 : array_update_81950[6];
  assign array_update_81963[7] = add_81474 == 32'h0000_0007 ? array_update_81961 : array_update_81950[7];
  assign array_update_81963[8] = add_81474 == 32'h0000_0008 ? array_update_81961 : array_update_81950[8];
  assign array_update_81963[9] = add_81474 == 32'h0000_0009 ? array_update_81961 : array_update_81950[9];
  assign array_index_81965 = array_update_72021[add_81962 > 32'h0000_0009 ? 4'h9 : add_81962[3:0]];
  assign array_index_81966 = array_update_81963[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_81970 = smul32b_32b_x_32b(array_index_81481[add_81962 > 32'h0000_0009 ? 4'h9 : add_81962[3:0]], array_index_81965[add_81882 > 32'h0000_0009 ? 4'h9 : add_81882[3:0]]);
  assign add_81972 = array_index_81966[add_81882 > 32'h0000_0009 ? 4'h9 : add_81882[3:0]] + smul_81970;
  assign array_update_81974[0] = add_81882 == 32'h0000_0000 ? add_81972 : array_index_81966[0];
  assign array_update_81974[1] = add_81882 == 32'h0000_0001 ? add_81972 : array_index_81966[1];
  assign array_update_81974[2] = add_81882 == 32'h0000_0002 ? add_81972 : array_index_81966[2];
  assign array_update_81974[3] = add_81882 == 32'h0000_0003 ? add_81972 : array_index_81966[3];
  assign array_update_81974[4] = add_81882 == 32'h0000_0004 ? add_81972 : array_index_81966[4];
  assign array_update_81974[5] = add_81882 == 32'h0000_0005 ? add_81972 : array_index_81966[5];
  assign array_update_81974[6] = add_81882 == 32'h0000_0006 ? add_81972 : array_index_81966[6];
  assign array_update_81974[7] = add_81882 == 32'h0000_0007 ? add_81972 : array_index_81966[7];
  assign array_update_81974[8] = add_81882 == 32'h0000_0008 ? add_81972 : array_index_81966[8];
  assign array_update_81974[9] = add_81882 == 32'h0000_0009 ? add_81972 : array_index_81966[9];
  assign add_81975 = add_81962 + 32'h0000_0001;
  assign array_update_81976[0] = add_81474 == 32'h0000_0000 ? array_update_81974 : array_update_81963[0];
  assign array_update_81976[1] = add_81474 == 32'h0000_0001 ? array_update_81974 : array_update_81963[1];
  assign array_update_81976[2] = add_81474 == 32'h0000_0002 ? array_update_81974 : array_update_81963[2];
  assign array_update_81976[3] = add_81474 == 32'h0000_0003 ? array_update_81974 : array_update_81963[3];
  assign array_update_81976[4] = add_81474 == 32'h0000_0004 ? array_update_81974 : array_update_81963[4];
  assign array_update_81976[5] = add_81474 == 32'h0000_0005 ? array_update_81974 : array_update_81963[5];
  assign array_update_81976[6] = add_81474 == 32'h0000_0006 ? array_update_81974 : array_update_81963[6];
  assign array_update_81976[7] = add_81474 == 32'h0000_0007 ? array_update_81974 : array_update_81963[7];
  assign array_update_81976[8] = add_81474 == 32'h0000_0008 ? array_update_81974 : array_update_81963[8];
  assign array_update_81976[9] = add_81474 == 32'h0000_0009 ? array_update_81974 : array_update_81963[9];
  assign array_index_81978 = array_update_72021[add_81975 > 32'h0000_0009 ? 4'h9 : add_81975[3:0]];
  assign array_index_81979 = array_update_81976[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_81983 = smul32b_32b_x_32b(array_index_81481[add_81975 > 32'h0000_0009 ? 4'h9 : add_81975[3:0]], array_index_81978[add_81882 > 32'h0000_0009 ? 4'h9 : add_81882[3:0]]);
  assign add_81985 = array_index_81979[add_81882 > 32'h0000_0009 ? 4'h9 : add_81882[3:0]] + smul_81983;
  assign array_update_81987[0] = add_81882 == 32'h0000_0000 ? add_81985 : array_index_81979[0];
  assign array_update_81987[1] = add_81882 == 32'h0000_0001 ? add_81985 : array_index_81979[1];
  assign array_update_81987[2] = add_81882 == 32'h0000_0002 ? add_81985 : array_index_81979[2];
  assign array_update_81987[3] = add_81882 == 32'h0000_0003 ? add_81985 : array_index_81979[3];
  assign array_update_81987[4] = add_81882 == 32'h0000_0004 ? add_81985 : array_index_81979[4];
  assign array_update_81987[5] = add_81882 == 32'h0000_0005 ? add_81985 : array_index_81979[5];
  assign array_update_81987[6] = add_81882 == 32'h0000_0006 ? add_81985 : array_index_81979[6];
  assign array_update_81987[7] = add_81882 == 32'h0000_0007 ? add_81985 : array_index_81979[7];
  assign array_update_81987[8] = add_81882 == 32'h0000_0008 ? add_81985 : array_index_81979[8];
  assign array_update_81987[9] = add_81882 == 32'h0000_0009 ? add_81985 : array_index_81979[9];
  assign add_81988 = add_81975 + 32'h0000_0001;
  assign array_update_81989[0] = add_81474 == 32'h0000_0000 ? array_update_81987 : array_update_81976[0];
  assign array_update_81989[1] = add_81474 == 32'h0000_0001 ? array_update_81987 : array_update_81976[1];
  assign array_update_81989[2] = add_81474 == 32'h0000_0002 ? array_update_81987 : array_update_81976[2];
  assign array_update_81989[3] = add_81474 == 32'h0000_0003 ? array_update_81987 : array_update_81976[3];
  assign array_update_81989[4] = add_81474 == 32'h0000_0004 ? array_update_81987 : array_update_81976[4];
  assign array_update_81989[5] = add_81474 == 32'h0000_0005 ? array_update_81987 : array_update_81976[5];
  assign array_update_81989[6] = add_81474 == 32'h0000_0006 ? array_update_81987 : array_update_81976[6];
  assign array_update_81989[7] = add_81474 == 32'h0000_0007 ? array_update_81987 : array_update_81976[7];
  assign array_update_81989[8] = add_81474 == 32'h0000_0008 ? array_update_81987 : array_update_81976[8];
  assign array_update_81989[9] = add_81474 == 32'h0000_0009 ? array_update_81987 : array_update_81976[9];
  assign array_index_81991 = array_update_72021[add_81988 > 32'h0000_0009 ? 4'h9 : add_81988[3:0]];
  assign array_index_81992 = array_update_81989[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_81996 = smul32b_32b_x_32b(array_index_81481[add_81988 > 32'h0000_0009 ? 4'h9 : add_81988[3:0]], array_index_81991[add_81882 > 32'h0000_0009 ? 4'h9 : add_81882[3:0]]);
  assign add_81998 = array_index_81992[add_81882 > 32'h0000_0009 ? 4'h9 : add_81882[3:0]] + smul_81996;
  assign array_update_82000[0] = add_81882 == 32'h0000_0000 ? add_81998 : array_index_81992[0];
  assign array_update_82000[1] = add_81882 == 32'h0000_0001 ? add_81998 : array_index_81992[1];
  assign array_update_82000[2] = add_81882 == 32'h0000_0002 ? add_81998 : array_index_81992[2];
  assign array_update_82000[3] = add_81882 == 32'h0000_0003 ? add_81998 : array_index_81992[3];
  assign array_update_82000[4] = add_81882 == 32'h0000_0004 ? add_81998 : array_index_81992[4];
  assign array_update_82000[5] = add_81882 == 32'h0000_0005 ? add_81998 : array_index_81992[5];
  assign array_update_82000[6] = add_81882 == 32'h0000_0006 ? add_81998 : array_index_81992[6];
  assign array_update_82000[7] = add_81882 == 32'h0000_0007 ? add_81998 : array_index_81992[7];
  assign array_update_82000[8] = add_81882 == 32'h0000_0008 ? add_81998 : array_index_81992[8];
  assign array_update_82000[9] = add_81882 == 32'h0000_0009 ? add_81998 : array_index_81992[9];
  assign add_82001 = add_81988 + 32'h0000_0001;
  assign array_update_82002[0] = add_81474 == 32'h0000_0000 ? array_update_82000 : array_update_81989[0];
  assign array_update_82002[1] = add_81474 == 32'h0000_0001 ? array_update_82000 : array_update_81989[1];
  assign array_update_82002[2] = add_81474 == 32'h0000_0002 ? array_update_82000 : array_update_81989[2];
  assign array_update_82002[3] = add_81474 == 32'h0000_0003 ? array_update_82000 : array_update_81989[3];
  assign array_update_82002[4] = add_81474 == 32'h0000_0004 ? array_update_82000 : array_update_81989[4];
  assign array_update_82002[5] = add_81474 == 32'h0000_0005 ? array_update_82000 : array_update_81989[5];
  assign array_update_82002[6] = add_81474 == 32'h0000_0006 ? array_update_82000 : array_update_81989[6];
  assign array_update_82002[7] = add_81474 == 32'h0000_0007 ? array_update_82000 : array_update_81989[7];
  assign array_update_82002[8] = add_81474 == 32'h0000_0008 ? array_update_82000 : array_update_81989[8];
  assign array_update_82002[9] = add_81474 == 32'h0000_0009 ? array_update_82000 : array_update_81989[9];
  assign array_index_82004 = array_update_72021[add_82001 > 32'h0000_0009 ? 4'h9 : add_82001[3:0]];
  assign array_index_82005 = array_update_82002[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_82009 = smul32b_32b_x_32b(array_index_81481[add_82001 > 32'h0000_0009 ? 4'h9 : add_82001[3:0]], array_index_82004[add_81882 > 32'h0000_0009 ? 4'h9 : add_81882[3:0]]);
  assign add_82011 = array_index_82005[add_81882 > 32'h0000_0009 ? 4'h9 : add_81882[3:0]] + smul_82009;
  assign array_update_82012[0] = add_81882 == 32'h0000_0000 ? add_82011 : array_index_82005[0];
  assign array_update_82012[1] = add_81882 == 32'h0000_0001 ? add_82011 : array_index_82005[1];
  assign array_update_82012[2] = add_81882 == 32'h0000_0002 ? add_82011 : array_index_82005[2];
  assign array_update_82012[3] = add_81882 == 32'h0000_0003 ? add_82011 : array_index_82005[3];
  assign array_update_82012[4] = add_81882 == 32'h0000_0004 ? add_82011 : array_index_82005[4];
  assign array_update_82012[5] = add_81882 == 32'h0000_0005 ? add_82011 : array_index_82005[5];
  assign array_update_82012[6] = add_81882 == 32'h0000_0006 ? add_82011 : array_index_82005[6];
  assign array_update_82012[7] = add_81882 == 32'h0000_0007 ? add_82011 : array_index_82005[7];
  assign array_update_82012[8] = add_81882 == 32'h0000_0008 ? add_82011 : array_index_82005[8];
  assign array_update_82012[9] = add_81882 == 32'h0000_0009 ? add_82011 : array_index_82005[9];
  assign array_update_82013[0] = add_81474 == 32'h0000_0000 ? array_update_82012 : array_update_82002[0];
  assign array_update_82013[1] = add_81474 == 32'h0000_0001 ? array_update_82012 : array_update_82002[1];
  assign array_update_82013[2] = add_81474 == 32'h0000_0002 ? array_update_82012 : array_update_82002[2];
  assign array_update_82013[3] = add_81474 == 32'h0000_0003 ? array_update_82012 : array_update_82002[3];
  assign array_update_82013[4] = add_81474 == 32'h0000_0004 ? array_update_82012 : array_update_82002[4];
  assign array_update_82013[5] = add_81474 == 32'h0000_0005 ? array_update_82012 : array_update_82002[5];
  assign array_update_82013[6] = add_81474 == 32'h0000_0006 ? array_update_82012 : array_update_82002[6];
  assign array_update_82013[7] = add_81474 == 32'h0000_0007 ? array_update_82012 : array_update_82002[7];
  assign array_update_82013[8] = add_81474 == 32'h0000_0008 ? array_update_82012 : array_update_82002[8];
  assign array_update_82013[9] = add_81474 == 32'h0000_0009 ? array_update_82012 : array_update_82002[9];
  assign array_index_82015 = array_update_82013[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign add_82017 = add_81882 + 32'h0000_0001;
  assign array_update_82018[0] = add_82017 == 32'h0000_0000 ? 32'h0000_0000 : array_index_82015[0];
  assign array_update_82018[1] = add_82017 == 32'h0000_0001 ? 32'h0000_0000 : array_index_82015[1];
  assign array_update_82018[2] = add_82017 == 32'h0000_0002 ? 32'h0000_0000 : array_index_82015[2];
  assign array_update_82018[3] = add_82017 == 32'h0000_0003 ? 32'h0000_0000 : array_index_82015[3];
  assign array_update_82018[4] = add_82017 == 32'h0000_0004 ? 32'h0000_0000 : array_index_82015[4];
  assign array_update_82018[5] = add_82017 == 32'h0000_0005 ? 32'h0000_0000 : array_index_82015[5];
  assign array_update_82018[6] = add_82017 == 32'h0000_0006 ? 32'h0000_0000 : array_index_82015[6];
  assign array_update_82018[7] = add_82017 == 32'h0000_0007 ? 32'h0000_0000 : array_index_82015[7];
  assign array_update_82018[8] = add_82017 == 32'h0000_0008 ? 32'h0000_0000 : array_index_82015[8];
  assign array_update_82018[9] = add_82017 == 32'h0000_0009 ? 32'h0000_0000 : array_index_82015[9];
  assign literal_82019 = 32'h0000_0000;
  assign array_update_82020[0] = add_81474 == 32'h0000_0000 ? array_update_82018 : array_update_82013[0];
  assign array_update_82020[1] = add_81474 == 32'h0000_0001 ? array_update_82018 : array_update_82013[1];
  assign array_update_82020[2] = add_81474 == 32'h0000_0002 ? array_update_82018 : array_update_82013[2];
  assign array_update_82020[3] = add_81474 == 32'h0000_0003 ? array_update_82018 : array_update_82013[3];
  assign array_update_82020[4] = add_81474 == 32'h0000_0004 ? array_update_82018 : array_update_82013[4];
  assign array_update_82020[5] = add_81474 == 32'h0000_0005 ? array_update_82018 : array_update_82013[5];
  assign array_update_82020[6] = add_81474 == 32'h0000_0006 ? array_update_82018 : array_update_82013[6];
  assign array_update_82020[7] = add_81474 == 32'h0000_0007 ? array_update_82018 : array_update_82013[7];
  assign array_update_82020[8] = add_81474 == 32'h0000_0008 ? array_update_82018 : array_update_82013[8];
  assign array_update_82020[9] = add_81474 == 32'h0000_0009 ? array_update_82018 : array_update_82013[9];
  assign array_index_82022 = array_update_72021[literal_82019 > 32'h0000_0009 ? 4'h9 : literal_82019[3:0]];
  assign array_index_82023 = array_update_82020[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_82027 = smul32b_32b_x_32b(array_index_81481[literal_82019 > 32'h0000_0009 ? 4'h9 : literal_82019[3:0]], array_index_82022[add_82017 > 32'h0000_0009 ? 4'h9 : add_82017[3:0]]);
  assign add_82029 = array_index_82023[add_82017 > 32'h0000_0009 ? 4'h9 : add_82017[3:0]] + smul_82027;
  assign array_update_82031[0] = add_82017 == 32'h0000_0000 ? add_82029 : array_index_82023[0];
  assign array_update_82031[1] = add_82017 == 32'h0000_0001 ? add_82029 : array_index_82023[1];
  assign array_update_82031[2] = add_82017 == 32'h0000_0002 ? add_82029 : array_index_82023[2];
  assign array_update_82031[3] = add_82017 == 32'h0000_0003 ? add_82029 : array_index_82023[3];
  assign array_update_82031[4] = add_82017 == 32'h0000_0004 ? add_82029 : array_index_82023[4];
  assign array_update_82031[5] = add_82017 == 32'h0000_0005 ? add_82029 : array_index_82023[5];
  assign array_update_82031[6] = add_82017 == 32'h0000_0006 ? add_82029 : array_index_82023[6];
  assign array_update_82031[7] = add_82017 == 32'h0000_0007 ? add_82029 : array_index_82023[7];
  assign array_update_82031[8] = add_82017 == 32'h0000_0008 ? add_82029 : array_index_82023[8];
  assign array_update_82031[9] = add_82017 == 32'h0000_0009 ? add_82029 : array_index_82023[9];
  assign add_82032 = literal_82019 + 32'h0000_0001;
  assign array_update_82033[0] = add_81474 == 32'h0000_0000 ? array_update_82031 : array_update_82020[0];
  assign array_update_82033[1] = add_81474 == 32'h0000_0001 ? array_update_82031 : array_update_82020[1];
  assign array_update_82033[2] = add_81474 == 32'h0000_0002 ? array_update_82031 : array_update_82020[2];
  assign array_update_82033[3] = add_81474 == 32'h0000_0003 ? array_update_82031 : array_update_82020[3];
  assign array_update_82033[4] = add_81474 == 32'h0000_0004 ? array_update_82031 : array_update_82020[4];
  assign array_update_82033[5] = add_81474 == 32'h0000_0005 ? array_update_82031 : array_update_82020[5];
  assign array_update_82033[6] = add_81474 == 32'h0000_0006 ? array_update_82031 : array_update_82020[6];
  assign array_update_82033[7] = add_81474 == 32'h0000_0007 ? array_update_82031 : array_update_82020[7];
  assign array_update_82033[8] = add_81474 == 32'h0000_0008 ? array_update_82031 : array_update_82020[8];
  assign array_update_82033[9] = add_81474 == 32'h0000_0009 ? array_update_82031 : array_update_82020[9];
  assign array_index_82035 = array_update_72021[add_82032 > 32'h0000_0009 ? 4'h9 : add_82032[3:0]];
  assign array_index_82036 = array_update_82033[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_82040 = smul32b_32b_x_32b(array_index_81481[add_82032 > 32'h0000_0009 ? 4'h9 : add_82032[3:0]], array_index_82035[add_82017 > 32'h0000_0009 ? 4'h9 : add_82017[3:0]]);
  assign add_82042 = array_index_82036[add_82017 > 32'h0000_0009 ? 4'h9 : add_82017[3:0]] + smul_82040;
  assign array_update_82044[0] = add_82017 == 32'h0000_0000 ? add_82042 : array_index_82036[0];
  assign array_update_82044[1] = add_82017 == 32'h0000_0001 ? add_82042 : array_index_82036[1];
  assign array_update_82044[2] = add_82017 == 32'h0000_0002 ? add_82042 : array_index_82036[2];
  assign array_update_82044[3] = add_82017 == 32'h0000_0003 ? add_82042 : array_index_82036[3];
  assign array_update_82044[4] = add_82017 == 32'h0000_0004 ? add_82042 : array_index_82036[4];
  assign array_update_82044[5] = add_82017 == 32'h0000_0005 ? add_82042 : array_index_82036[5];
  assign array_update_82044[6] = add_82017 == 32'h0000_0006 ? add_82042 : array_index_82036[6];
  assign array_update_82044[7] = add_82017 == 32'h0000_0007 ? add_82042 : array_index_82036[7];
  assign array_update_82044[8] = add_82017 == 32'h0000_0008 ? add_82042 : array_index_82036[8];
  assign array_update_82044[9] = add_82017 == 32'h0000_0009 ? add_82042 : array_index_82036[9];
  assign add_82045 = add_82032 + 32'h0000_0001;
  assign array_update_82046[0] = add_81474 == 32'h0000_0000 ? array_update_82044 : array_update_82033[0];
  assign array_update_82046[1] = add_81474 == 32'h0000_0001 ? array_update_82044 : array_update_82033[1];
  assign array_update_82046[2] = add_81474 == 32'h0000_0002 ? array_update_82044 : array_update_82033[2];
  assign array_update_82046[3] = add_81474 == 32'h0000_0003 ? array_update_82044 : array_update_82033[3];
  assign array_update_82046[4] = add_81474 == 32'h0000_0004 ? array_update_82044 : array_update_82033[4];
  assign array_update_82046[5] = add_81474 == 32'h0000_0005 ? array_update_82044 : array_update_82033[5];
  assign array_update_82046[6] = add_81474 == 32'h0000_0006 ? array_update_82044 : array_update_82033[6];
  assign array_update_82046[7] = add_81474 == 32'h0000_0007 ? array_update_82044 : array_update_82033[7];
  assign array_update_82046[8] = add_81474 == 32'h0000_0008 ? array_update_82044 : array_update_82033[8];
  assign array_update_82046[9] = add_81474 == 32'h0000_0009 ? array_update_82044 : array_update_82033[9];
  assign array_index_82048 = array_update_72021[add_82045 > 32'h0000_0009 ? 4'h9 : add_82045[3:0]];
  assign array_index_82049 = array_update_82046[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_82053 = smul32b_32b_x_32b(array_index_81481[add_82045 > 32'h0000_0009 ? 4'h9 : add_82045[3:0]], array_index_82048[add_82017 > 32'h0000_0009 ? 4'h9 : add_82017[3:0]]);
  assign add_82055 = array_index_82049[add_82017 > 32'h0000_0009 ? 4'h9 : add_82017[3:0]] + smul_82053;
  assign array_update_82057[0] = add_82017 == 32'h0000_0000 ? add_82055 : array_index_82049[0];
  assign array_update_82057[1] = add_82017 == 32'h0000_0001 ? add_82055 : array_index_82049[1];
  assign array_update_82057[2] = add_82017 == 32'h0000_0002 ? add_82055 : array_index_82049[2];
  assign array_update_82057[3] = add_82017 == 32'h0000_0003 ? add_82055 : array_index_82049[3];
  assign array_update_82057[4] = add_82017 == 32'h0000_0004 ? add_82055 : array_index_82049[4];
  assign array_update_82057[5] = add_82017 == 32'h0000_0005 ? add_82055 : array_index_82049[5];
  assign array_update_82057[6] = add_82017 == 32'h0000_0006 ? add_82055 : array_index_82049[6];
  assign array_update_82057[7] = add_82017 == 32'h0000_0007 ? add_82055 : array_index_82049[7];
  assign array_update_82057[8] = add_82017 == 32'h0000_0008 ? add_82055 : array_index_82049[8];
  assign array_update_82057[9] = add_82017 == 32'h0000_0009 ? add_82055 : array_index_82049[9];
  assign add_82058 = add_82045 + 32'h0000_0001;
  assign array_update_82059[0] = add_81474 == 32'h0000_0000 ? array_update_82057 : array_update_82046[0];
  assign array_update_82059[1] = add_81474 == 32'h0000_0001 ? array_update_82057 : array_update_82046[1];
  assign array_update_82059[2] = add_81474 == 32'h0000_0002 ? array_update_82057 : array_update_82046[2];
  assign array_update_82059[3] = add_81474 == 32'h0000_0003 ? array_update_82057 : array_update_82046[3];
  assign array_update_82059[4] = add_81474 == 32'h0000_0004 ? array_update_82057 : array_update_82046[4];
  assign array_update_82059[5] = add_81474 == 32'h0000_0005 ? array_update_82057 : array_update_82046[5];
  assign array_update_82059[6] = add_81474 == 32'h0000_0006 ? array_update_82057 : array_update_82046[6];
  assign array_update_82059[7] = add_81474 == 32'h0000_0007 ? array_update_82057 : array_update_82046[7];
  assign array_update_82059[8] = add_81474 == 32'h0000_0008 ? array_update_82057 : array_update_82046[8];
  assign array_update_82059[9] = add_81474 == 32'h0000_0009 ? array_update_82057 : array_update_82046[9];
  assign array_index_82061 = array_update_72021[add_82058 > 32'h0000_0009 ? 4'h9 : add_82058[3:0]];
  assign array_index_82062 = array_update_82059[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_82066 = smul32b_32b_x_32b(array_index_81481[add_82058 > 32'h0000_0009 ? 4'h9 : add_82058[3:0]], array_index_82061[add_82017 > 32'h0000_0009 ? 4'h9 : add_82017[3:0]]);
  assign add_82068 = array_index_82062[add_82017 > 32'h0000_0009 ? 4'h9 : add_82017[3:0]] + smul_82066;
  assign array_update_82070[0] = add_82017 == 32'h0000_0000 ? add_82068 : array_index_82062[0];
  assign array_update_82070[1] = add_82017 == 32'h0000_0001 ? add_82068 : array_index_82062[1];
  assign array_update_82070[2] = add_82017 == 32'h0000_0002 ? add_82068 : array_index_82062[2];
  assign array_update_82070[3] = add_82017 == 32'h0000_0003 ? add_82068 : array_index_82062[3];
  assign array_update_82070[4] = add_82017 == 32'h0000_0004 ? add_82068 : array_index_82062[4];
  assign array_update_82070[5] = add_82017 == 32'h0000_0005 ? add_82068 : array_index_82062[5];
  assign array_update_82070[6] = add_82017 == 32'h0000_0006 ? add_82068 : array_index_82062[6];
  assign array_update_82070[7] = add_82017 == 32'h0000_0007 ? add_82068 : array_index_82062[7];
  assign array_update_82070[8] = add_82017 == 32'h0000_0008 ? add_82068 : array_index_82062[8];
  assign array_update_82070[9] = add_82017 == 32'h0000_0009 ? add_82068 : array_index_82062[9];
  assign add_82071 = add_82058 + 32'h0000_0001;
  assign array_update_82072[0] = add_81474 == 32'h0000_0000 ? array_update_82070 : array_update_82059[0];
  assign array_update_82072[1] = add_81474 == 32'h0000_0001 ? array_update_82070 : array_update_82059[1];
  assign array_update_82072[2] = add_81474 == 32'h0000_0002 ? array_update_82070 : array_update_82059[2];
  assign array_update_82072[3] = add_81474 == 32'h0000_0003 ? array_update_82070 : array_update_82059[3];
  assign array_update_82072[4] = add_81474 == 32'h0000_0004 ? array_update_82070 : array_update_82059[4];
  assign array_update_82072[5] = add_81474 == 32'h0000_0005 ? array_update_82070 : array_update_82059[5];
  assign array_update_82072[6] = add_81474 == 32'h0000_0006 ? array_update_82070 : array_update_82059[6];
  assign array_update_82072[7] = add_81474 == 32'h0000_0007 ? array_update_82070 : array_update_82059[7];
  assign array_update_82072[8] = add_81474 == 32'h0000_0008 ? array_update_82070 : array_update_82059[8];
  assign array_update_82072[9] = add_81474 == 32'h0000_0009 ? array_update_82070 : array_update_82059[9];
  assign array_index_82074 = array_update_72021[add_82071 > 32'h0000_0009 ? 4'h9 : add_82071[3:0]];
  assign array_index_82075 = array_update_82072[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_82079 = smul32b_32b_x_32b(array_index_81481[add_82071 > 32'h0000_0009 ? 4'h9 : add_82071[3:0]], array_index_82074[add_82017 > 32'h0000_0009 ? 4'h9 : add_82017[3:0]]);
  assign add_82081 = array_index_82075[add_82017 > 32'h0000_0009 ? 4'h9 : add_82017[3:0]] + smul_82079;
  assign array_update_82083[0] = add_82017 == 32'h0000_0000 ? add_82081 : array_index_82075[0];
  assign array_update_82083[1] = add_82017 == 32'h0000_0001 ? add_82081 : array_index_82075[1];
  assign array_update_82083[2] = add_82017 == 32'h0000_0002 ? add_82081 : array_index_82075[2];
  assign array_update_82083[3] = add_82017 == 32'h0000_0003 ? add_82081 : array_index_82075[3];
  assign array_update_82083[4] = add_82017 == 32'h0000_0004 ? add_82081 : array_index_82075[4];
  assign array_update_82083[5] = add_82017 == 32'h0000_0005 ? add_82081 : array_index_82075[5];
  assign array_update_82083[6] = add_82017 == 32'h0000_0006 ? add_82081 : array_index_82075[6];
  assign array_update_82083[7] = add_82017 == 32'h0000_0007 ? add_82081 : array_index_82075[7];
  assign array_update_82083[8] = add_82017 == 32'h0000_0008 ? add_82081 : array_index_82075[8];
  assign array_update_82083[9] = add_82017 == 32'h0000_0009 ? add_82081 : array_index_82075[9];
  assign add_82084 = add_82071 + 32'h0000_0001;
  assign array_update_82085[0] = add_81474 == 32'h0000_0000 ? array_update_82083 : array_update_82072[0];
  assign array_update_82085[1] = add_81474 == 32'h0000_0001 ? array_update_82083 : array_update_82072[1];
  assign array_update_82085[2] = add_81474 == 32'h0000_0002 ? array_update_82083 : array_update_82072[2];
  assign array_update_82085[3] = add_81474 == 32'h0000_0003 ? array_update_82083 : array_update_82072[3];
  assign array_update_82085[4] = add_81474 == 32'h0000_0004 ? array_update_82083 : array_update_82072[4];
  assign array_update_82085[5] = add_81474 == 32'h0000_0005 ? array_update_82083 : array_update_82072[5];
  assign array_update_82085[6] = add_81474 == 32'h0000_0006 ? array_update_82083 : array_update_82072[6];
  assign array_update_82085[7] = add_81474 == 32'h0000_0007 ? array_update_82083 : array_update_82072[7];
  assign array_update_82085[8] = add_81474 == 32'h0000_0008 ? array_update_82083 : array_update_82072[8];
  assign array_update_82085[9] = add_81474 == 32'h0000_0009 ? array_update_82083 : array_update_82072[9];
  assign array_index_82087 = array_update_72021[add_82084 > 32'h0000_0009 ? 4'h9 : add_82084[3:0]];
  assign array_index_82088 = array_update_82085[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_82092 = smul32b_32b_x_32b(array_index_81481[add_82084 > 32'h0000_0009 ? 4'h9 : add_82084[3:0]], array_index_82087[add_82017 > 32'h0000_0009 ? 4'h9 : add_82017[3:0]]);
  assign add_82094 = array_index_82088[add_82017 > 32'h0000_0009 ? 4'h9 : add_82017[3:0]] + smul_82092;
  assign array_update_82096[0] = add_82017 == 32'h0000_0000 ? add_82094 : array_index_82088[0];
  assign array_update_82096[1] = add_82017 == 32'h0000_0001 ? add_82094 : array_index_82088[1];
  assign array_update_82096[2] = add_82017 == 32'h0000_0002 ? add_82094 : array_index_82088[2];
  assign array_update_82096[3] = add_82017 == 32'h0000_0003 ? add_82094 : array_index_82088[3];
  assign array_update_82096[4] = add_82017 == 32'h0000_0004 ? add_82094 : array_index_82088[4];
  assign array_update_82096[5] = add_82017 == 32'h0000_0005 ? add_82094 : array_index_82088[5];
  assign array_update_82096[6] = add_82017 == 32'h0000_0006 ? add_82094 : array_index_82088[6];
  assign array_update_82096[7] = add_82017 == 32'h0000_0007 ? add_82094 : array_index_82088[7];
  assign array_update_82096[8] = add_82017 == 32'h0000_0008 ? add_82094 : array_index_82088[8];
  assign array_update_82096[9] = add_82017 == 32'h0000_0009 ? add_82094 : array_index_82088[9];
  assign add_82097 = add_82084 + 32'h0000_0001;
  assign array_update_82098[0] = add_81474 == 32'h0000_0000 ? array_update_82096 : array_update_82085[0];
  assign array_update_82098[1] = add_81474 == 32'h0000_0001 ? array_update_82096 : array_update_82085[1];
  assign array_update_82098[2] = add_81474 == 32'h0000_0002 ? array_update_82096 : array_update_82085[2];
  assign array_update_82098[3] = add_81474 == 32'h0000_0003 ? array_update_82096 : array_update_82085[3];
  assign array_update_82098[4] = add_81474 == 32'h0000_0004 ? array_update_82096 : array_update_82085[4];
  assign array_update_82098[5] = add_81474 == 32'h0000_0005 ? array_update_82096 : array_update_82085[5];
  assign array_update_82098[6] = add_81474 == 32'h0000_0006 ? array_update_82096 : array_update_82085[6];
  assign array_update_82098[7] = add_81474 == 32'h0000_0007 ? array_update_82096 : array_update_82085[7];
  assign array_update_82098[8] = add_81474 == 32'h0000_0008 ? array_update_82096 : array_update_82085[8];
  assign array_update_82098[9] = add_81474 == 32'h0000_0009 ? array_update_82096 : array_update_82085[9];
  assign array_index_82100 = array_update_72021[add_82097 > 32'h0000_0009 ? 4'h9 : add_82097[3:0]];
  assign array_index_82101 = array_update_82098[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_82105 = smul32b_32b_x_32b(array_index_81481[add_82097 > 32'h0000_0009 ? 4'h9 : add_82097[3:0]], array_index_82100[add_82017 > 32'h0000_0009 ? 4'h9 : add_82017[3:0]]);
  assign add_82107 = array_index_82101[add_82017 > 32'h0000_0009 ? 4'h9 : add_82017[3:0]] + smul_82105;
  assign array_update_82109[0] = add_82017 == 32'h0000_0000 ? add_82107 : array_index_82101[0];
  assign array_update_82109[1] = add_82017 == 32'h0000_0001 ? add_82107 : array_index_82101[1];
  assign array_update_82109[2] = add_82017 == 32'h0000_0002 ? add_82107 : array_index_82101[2];
  assign array_update_82109[3] = add_82017 == 32'h0000_0003 ? add_82107 : array_index_82101[3];
  assign array_update_82109[4] = add_82017 == 32'h0000_0004 ? add_82107 : array_index_82101[4];
  assign array_update_82109[5] = add_82017 == 32'h0000_0005 ? add_82107 : array_index_82101[5];
  assign array_update_82109[6] = add_82017 == 32'h0000_0006 ? add_82107 : array_index_82101[6];
  assign array_update_82109[7] = add_82017 == 32'h0000_0007 ? add_82107 : array_index_82101[7];
  assign array_update_82109[8] = add_82017 == 32'h0000_0008 ? add_82107 : array_index_82101[8];
  assign array_update_82109[9] = add_82017 == 32'h0000_0009 ? add_82107 : array_index_82101[9];
  assign add_82110 = add_82097 + 32'h0000_0001;
  assign array_update_82111[0] = add_81474 == 32'h0000_0000 ? array_update_82109 : array_update_82098[0];
  assign array_update_82111[1] = add_81474 == 32'h0000_0001 ? array_update_82109 : array_update_82098[1];
  assign array_update_82111[2] = add_81474 == 32'h0000_0002 ? array_update_82109 : array_update_82098[2];
  assign array_update_82111[3] = add_81474 == 32'h0000_0003 ? array_update_82109 : array_update_82098[3];
  assign array_update_82111[4] = add_81474 == 32'h0000_0004 ? array_update_82109 : array_update_82098[4];
  assign array_update_82111[5] = add_81474 == 32'h0000_0005 ? array_update_82109 : array_update_82098[5];
  assign array_update_82111[6] = add_81474 == 32'h0000_0006 ? array_update_82109 : array_update_82098[6];
  assign array_update_82111[7] = add_81474 == 32'h0000_0007 ? array_update_82109 : array_update_82098[7];
  assign array_update_82111[8] = add_81474 == 32'h0000_0008 ? array_update_82109 : array_update_82098[8];
  assign array_update_82111[9] = add_81474 == 32'h0000_0009 ? array_update_82109 : array_update_82098[9];
  assign array_index_82113 = array_update_72021[add_82110 > 32'h0000_0009 ? 4'h9 : add_82110[3:0]];
  assign array_index_82114 = array_update_82111[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_82118 = smul32b_32b_x_32b(array_index_81481[add_82110 > 32'h0000_0009 ? 4'h9 : add_82110[3:0]], array_index_82113[add_82017 > 32'h0000_0009 ? 4'h9 : add_82017[3:0]]);
  assign add_82120 = array_index_82114[add_82017 > 32'h0000_0009 ? 4'h9 : add_82017[3:0]] + smul_82118;
  assign array_update_82122[0] = add_82017 == 32'h0000_0000 ? add_82120 : array_index_82114[0];
  assign array_update_82122[1] = add_82017 == 32'h0000_0001 ? add_82120 : array_index_82114[1];
  assign array_update_82122[2] = add_82017 == 32'h0000_0002 ? add_82120 : array_index_82114[2];
  assign array_update_82122[3] = add_82017 == 32'h0000_0003 ? add_82120 : array_index_82114[3];
  assign array_update_82122[4] = add_82017 == 32'h0000_0004 ? add_82120 : array_index_82114[4];
  assign array_update_82122[5] = add_82017 == 32'h0000_0005 ? add_82120 : array_index_82114[5];
  assign array_update_82122[6] = add_82017 == 32'h0000_0006 ? add_82120 : array_index_82114[6];
  assign array_update_82122[7] = add_82017 == 32'h0000_0007 ? add_82120 : array_index_82114[7];
  assign array_update_82122[8] = add_82017 == 32'h0000_0008 ? add_82120 : array_index_82114[8];
  assign array_update_82122[9] = add_82017 == 32'h0000_0009 ? add_82120 : array_index_82114[9];
  assign add_82123 = add_82110 + 32'h0000_0001;
  assign array_update_82124[0] = add_81474 == 32'h0000_0000 ? array_update_82122 : array_update_82111[0];
  assign array_update_82124[1] = add_81474 == 32'h0000_0001 ? array_update_82122 : array_update_82111[1];
  assign array_update_82124[2] = add_81474 == 32'h0000_0002 ? array_update_82122 : array_update_82111[2];
  assign array_update_82124[3] = add_81474 == 32'h0000_0003 ? array_update_82122 : array_update_82111[3];
  assign array_update_82124[4] = add_81474 == 32'h0000_0004 ? array_update_82122 : array_update_82111[4];
  assign array_update_82124[5] = add_81474 == 32'h0000_0005 ? array_update_82122 : array_update_82111[5];
  assign array_update_82124[6] = add_81474 == 32'h0000_0006 ? array_update_82122 : array_update_82111[6];
  assign array_update_82124[7] = add_81474 == 32'h0000_0007 ? array_update_82122 : array_update_82111[7];
  assign array_update_82124[8] = add_81474 == 32'h0000_0008 ? array_update_82122 : array_update_82111[8];
  assign array_update_82124[9] = add_81474 == 32'h0000_0009 ? array_update_82122 : array_update_82111[9];
  assign array_index_82126 = array_update_72021[add_82123 > 32'h0000_0009 ? 4'h9 : add_82123[3:0]];
  assign array_index_82127 = array_update_82124[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_82131 = smul32b_32b_x_32b(array_index_81481[add_82123 > 32'h0000_0009 ? 4'h9 : add_82123[3:0]], array_index_82126[add_82017 > 32'h0000_0009 ? 4'h9 : add_82017[3:0]]);
  assign add_82133 = array_index_82127[add_82017 > 32'h0000_0009 ? 4'h9 : add_82017[3:0]] + smul_82131;
  assign array_update_82135[0] = add_82017 == 32'h0000_0000 ? add_82133 : array_index_82127[0];
  assign array_update_82135[1] = add_82017 == 32'h0000_0001 ? add_82133 : array_index_82127[1];
  assign array_update_82135[2] = add_82017 == 32'h0000_0002 ? add_82133 : array_index_82127[2];
  assign array_update_82135[3] = add_82017 == 32'h0000_0003 ? add_82133 : array_index_82127[3];
  assign array_update_82135[4] = add_82017 == 32'h0000_0004 ? add_82133 : array_index_82127[4];
  assign array_update_82135[5] = add_82017 == 32'h0000_0005 ? add_82133 : array_index_82127[5];
  assign array_update_82135[6] = add_82017 == 32'h0000_0006 ? add_82133 : array_index_82127[6];
  assign array_update_82135[7] = add_82017 == 32'h0000_0007 ? add_82133 : array_index_82127[7];
  assign array_update_82135[8] = add_82017 == 32'h0000_0008 ? add_82133 : array_index_82127[8];
  assign array_update_82135[9] = add_82017 == 32'h0000_0009 ? add_82133 : array_index_82127[9];
  assign add_82136 = add_82123 + 32'h0000_0001;
  assign array_update_82137[0] = add_81474 == 32'h0000_0000 ? array_update_82135 : array_update_82124[0];
  assign array_update_82137[1] = add_81474 == 32'h0000_0001 ? array_update_82135 : array_update_82124[1];
  assign array_update_82137[2] = add_81474 == 32'h0000_0002 ? array_update_82135 : array_update_82124[2];
  assign array_update_82137[3] = add_81474 == 32'h0000_0003 ? array_update_82135 : array_update_82124[3];
  assign array_update_82137[4] = add_81474 == 32'h0000_0004 ? array_update_82135 : array_update_82124[4];
  assign array_update_82137[5] = add_81474 == 32'h0000_0005 ? array_update_82135 : array_update_82124[5];
  assign array_update_82137[6] = add_81474 == 32'h0000_0006 ? array_update_82135 : array_update_82124[6];
  assign array_update_82137[7] = add_81474 == 32'h0000_0007 ? array_update_82135 : array_update_82124[7];
  assign array_update_82137[8] = add_81474 == 32'h0000_0008 ? array_update_82135 : array_update_82124[8];
  assign array_update_82137[9] = add_81474 == 32'h0000_0009 ? array_update_82135 : array_update_82124[9];
  assign array_index_82139 = array_update_72021[add_82136 > 32'h0000_0009 ? 4'h9 : add_82136[3:0]];
  assign array_index_82140 = array_update_82137[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_82144 = smul32b_32b_x_32b(array_index_81481[add_82136 > 32'h0000_0009 ? 4'h9 : add_82136[3:0]], array_index_82139[add_82017 > 32'h0000_0009 ? 4'h9 : add_82017[3:0]]);
  assign add_82146 = array_index_82140[add_82017 > 32'h0000_0009 ? 4'h9 : add_82017[3:0]] + smul_82144;
  assign array_update_82147[0] = add_82017 == 32'h0000_0000 ? add_82146 : array_index_82140[0];
  assign array_update_82147[1] = add_82017 == 32'h0000_0001 ? add_82146 : array_index_82140[1];
  assign array_update_82147[2] = add_82017 == 32'h0000_0002 ? add_82146 : array_index_82140[2];
  assign array_update_82147[3] = add_82017 == 32'h0000_0003 ? add_82146 : array_index_82140[3];
  assign array_update_82147[4] = add_82017 == 32'h0000_0004 ? add_82146 : array_index_82140[4];
  assign array_update_82147[5] = add_82017 == 32'h0000_0005 ? add_82146 : array_index_82140[5];
  assign array_update_82147[6] = add_82017 == 32'h0000_0006 ? add_82146 : array_index_82140[6];
  assign array_update_82147[7] = add_82017 == 32'h0000_0007 ? add_82146 : array_index_82140[7];
  assign array_update_82147[8] = add_82017 == 32'h0000_0008 ? add_82146 : array_index_82140[8];
  assign array_update_82147[9] = add_82017 == 32'h0000_0009 ? add_82146 : array_index_82140[9];
  assign array_update_82148[0] = add_81474 == 32'h0000_0000 ? array_update_82147 : array_update_82137[0];
  assign array_update_82148[1] = add_81474 == 32'h0000_0001 ? array_update_82147 : array_update_82137[1];
  assign array_update_82148[2] = add_81474 == 32'h0000_0002 ? array_update_82147 : array_update_82137[2];
  assign array_update_82148[3] = add_81474 == 32'h0000_0003 ? array_update_82147 : array_update_82137[3];
  assign array_update_82148[4] = add_81474 == 32'h0000_0004 ? array_update_82147 : array_update_82137[4];
  assign array_update_82148[5] = add_81474 == 32'h0000_0005 ? array_update_82147 : array_update_82137[5];
  assign array_update_82148[6] = add_81474 == 32'h0000_0006 ? array_update_82147 : array_update_82137[6];
  assign array_update_82148[7] = add_81474 == 32'h0000_0007 ? array_update_82147 : array_update_82137[7];
  assign array_update_82148[8] = add_81474 == 32'h0000_0008 ? array_update_82147 : array_update_82137[8];
  assign array_update_82148[9] = add_81474 == 32'h0000_0009 ? array_update_82147 : array_update_82137[9];
  assign array_index_82150 = array_update_82148[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign add_82152 = add_82017 + 32'h0000_0001;
  assign array_update_82153[0] = add_82152 == 32'h0000_0000 ? 32'h0000_0000 : array_index_82150[0];
  assign array_update_82153[1] = add_82152 == 32'h0000_0001 ? 32'h0000_0000 : array_index_82150[1];
  assign array_update_82153[2] = add_82152 == 32'h0000_0002 ? 32'h0000_0000 : array_index_82150[2];
  assign array_update_82153[3] = add_82152 == 32'h0000_0003 ? 32'h0000_0000 : array_index_82150[3];
  assign array_update_82153[4] = add_82152 == 32'h0000_0004 ? 32'h0000_0000 : array_index_82150[4];
  assign array_update_82153[5] = add_82152 == 32'h0000_0005 ? 32'h0000_0000 : array_index_82150[5];
  assign array_update_82153[6] = add_82152 == 32'h0000_0006 ? 32'h0000_0000 : array_index_82150[6];
  assign array_update_82153[7] = add_82152 == 32'h0000_0007 ? 32'h0000_0000 : array_index_82150[7];
  assign array_update_82153[8] = add_82152 == 32'h0000_0008 ? 32'h0000_0000 : array_index_82150[8];
  assign array_update_82153[9] = add_82152 == 32'h0000_0009 ? 32'h0000_0000 : array_index_82150[9];
  assign literal_82154 = 32'h0000_0000;
  assign array_update_82155[0] = add_81474 == 32'h0000_0000 ? array_update_82153 : array_update_82148[0];
  assign array_update_82155[1] = add_81474 == 32'h0000_0001 ? array_update_82153 : array_update_82148[1];
  assign array_update_82155[2] = add_81474 == 32'h0000_0002 ? array_update_82153 : array_update_82148[2];
  assign array_update_82155[3] = add_81474 == 32'h0000_0003 ? array_update_82153 : array_update_82148[3];
  assign array_update_82155[4] = add_81474 == 32'h0000_0004 ? array_update_82153 : array_update_82148[4];
  assign array_update_82155[5] = add_81474 == 32'h0000_0005 ? array_update_82153 : array_update_82148[5];
  assign array_update_82155[6] = add_81474 == 32'h0000_0006 ? array_update_82153 : array_update_82148[6];
  assign array_update_82155[7] = add_81474 == 32'h0000_0007 ? array_update_82153 : array_update_82148[7];
  assign array_update_82155[8] = add_81474 == 32'h0000_0008 ? array_update_82153 : array_update_82148[8];
  assign array_update_82155[9] = add_81474 == 32'h0000_0009 ? array_update_82153 : array_update_82148[9];
  assign array_index_82157 = array_update_72021[literal_82154 > 32'h0000_0009 ? 4'h9 : literal_82154[3:0]];
  assign array_index_82158 = array_update_82155[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_82162 = smul32b_32b_x_32b(array_index_81481[literal_82154 > 32'h0000_0009 ? 4'h9 : literal_82154[3:0]], array_index_82157[add_82152 > 32'h0000_0009 ? 4'h9 : add_82152[3:0]]);
  assign add_82164 = array_index_82158[add_82152 > 32'h0000_0009 ? 4'h9 : add_82152[3:0]] + smul_82162;
  assign array_update_82166[0] = add_82152 == 32'h0000_0000 ? add_82164 : array_index_82158[0];
  assign array_update_82166[1] = add_82152 == 32'h0000_0001 ? add_82164 : array_index_82158[1];
  assign array_update_82166[2] = add_82152 == 32'h0000_0002 ? add_82164 : array_index_82158[2];
  assign array_update_82166[3] = add_82152 == 32'h0000_0003 ? add_82164 : array_index_82158[3];
  assign array_update_82166[4] = add_82152 == 32'h0000_0004 ? add_82164 : array_index_82158[4];
  assign array_update_82166[5] = add_82152 == 32'h0000_0005 ? add_82164 : array_index_82158[5];
  assign array_update_82166[6] = add_82152 == 32'h0000_0006 ? add_82164 : array_index_82158[6];
  assign array_update_82166[7] = add_82152 == 32'h0000_0007 ? add_82164 : array_index_82158[7];
  assign array_update_82166[8] = add_82152 == 32'h0000_0008 ? add_82164 : array_index_82158[8];
  assign array_update_82166[9] = add_82152 == 32'h0000_0009 ? add_82164 : array_index_82158[9];
  assign add_82167 = literal_82154 + 32'h0000_0001;
  assign array_update_82168[0] = add_81474 == 32'h0000_0000 ? array_update_82166 : array_update_82155[0];
  assign array_update_82168[1] = add_81474 == 32'h0000_0001 ? array_update_82166 : array_update_82155[1];
  assign array_update_82168[2] = add_81474 == 32'h0000_0002 ? array_update_82166 : array_update_82155[2];
  assign array_update_82168[3] = add_81474 == 32'h0000_0003 ? array_update_82166 : array_update_82155[3];
  assign array_update_82168[4] = add_81474 == 32'h0000_0004 ? array_update_82166 : array_update_82155[4];
  assign array_update_82168[5] = add_81474 == 32'h0000_0005 ? array_update_82166 : array_update_82155[5];
  assign array_update_82168[6] = add_81474 == 32'h0000_0006 ? array_update_82166 : array_update_82155[6];
  assign array_update_82168[7] = add_81474 == 32'h0000_0007 ? array_update_82166 : array_update_82155[7];
  assign array_update_82168[8] = add_81474 == 32'h0000_0008 ? array_update_82166 : array_update_82155[8];
  assign array_update_82168[9] = add_81474 == 32'h0000_0009 ? array_update_82166 : array_update_82155[9];
  assign array_index_82170 = array_update_72021[add_82167 > 32'h0000_0009 ? 4'h9 : add_82167[3:0]];
  assign array_index_82171 = array_update_82168[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_82175 = smul32b_32b_x_32b(array_index_81481[add_82167 > 32'h0000_0009 ? 4'h9 : add_82167[3:0]], array_index_82170[add_82152 > 32'h0000_0009 ? 4'h9 : add_82152[3:0]]);
  assign add_82177 = array_index_82171[add_82152 > 32'h0000_0009 ? 4'h9 : add_82152[3:0]] + smul_82175;
  assign array_update_82179[0] = add_82152 == 32'h0000_0000 ? add_82177 : array_index_82171[0];
  assign array_update_82179[1] = add_82152 == 32'h0000_0001 ? add_82177 : array_index_82171[1];
  assign array_update_82179[2] = add_82152 == 32'h0000_0002 ? add_82177 : array_index_82171[2];
  assign array_update_82179[3] = add_82152 == 32'h0000_0003 ? add_82177 : array_index_82171[3];
  assign array_update_82179[4] = add_82152 == 32'h0000_0004 ? add_82177 : array_index_82171[4];
  assign array_update_82179[5] = add_82152 == 32'h0000_0005 ? add_82177 : array_index_82171[5];
  assign array_update_82179[6] = add_82152 == 32'h0000_0006 ? add_82177 : array_index_82171[6];
  assign array_update_82179[7] = add_82152 == 32'h0000_0007 ? add_82177 : array_index_82171[7];
  assign array_update_82179[8] = add_82152 == 32'h0000_0008 ? add_82177 : array_index_82171[8];
  assign array_update_82179[9] = add_82152 == 32'h0000_0009 ? add_82177 : array_index_82171[9];
  assign add_82180 = add_82167 + 32'h0000_0001;
  assign array_update_82181[0] = add_81474 == 32'h0000_0000 ? array_update_82179 : array_update_82168[0];
  assign array_update_82181[1] = add_81474 == 32'h0000_0001 ? array_update_82179 : array_update_82168[1];
  assign array_update_82181[2] = add_81474 == 32'h0000_0002 ? array_update_82179 : array_update_82168[2];
  assign array_update_82181[3] = add_81474 == 32'h0000_0003 ? array_update_82179 : array_update_82168[3];
  assign array_update_82181[4] = add_81474 == 32'h0000_0004 ? array_update_82179 : array_update_82168[4];
  assign array_update_82181[5] = add_81474 == 32'h0000_0005 ? array_update_82179 : array_update_82168[5];
  assign array_update_82181[6] = add_81474 == 32'h0000_0006 ? array_update_82179 : array_update_82168[6];
  assign array_update_82181[7] = add_81474 == 32'h0000_0007 ? array_update_82179 : array_update_82168[7];
  assign array_update_82181[8] = add_81474 == 32'h0000_0008 ? array_update_82179 : array_update_82168[8];
  assign array_update_82181[9] = add_81474 == 32'h0000_0009 ? array_update_82179 : array_update_82168[9];
  assign array_index_82183 = array_update_72021[add_82180 > 32'h0000_0009 ? 4'h9 : add_82180[3:0]];
  assign array_index_82184 = array_update_82181[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_82188 = smul32b_32b_x_32b(array_index_81481[add_82180 > 32'h0000_0009 ? 4'h9 : add_82180[3:0]], array_index_82183[add_82152 > 32'h0000_0009 ? 4'h9 : add_82152[3:0]]);
  assign add_82190 = array_index_82184[add_82152 > 32'h0000_0009 ? 4'h9 : add_82152[3:0]] + smul_82188;
  assign array_update_82192[0] = add_82152 == 32'h0000_0000 ? add_82190 : array_index_82184[0];
  assign array_update_82192[1] = add_82152 == 32'h0000_0001 ? add_82190 : array_index_82184[1];
  assign array_update_82192[2] = add_82152 == 32'h0000_0002 ? add_82190 : array_index_82184[2];
  assign array_update_82192[3] = add_82152 == 32'h0000_0003 ? add_82190 : array_index_82184[3];
  assign array_update_82192[4] = add_82152 == 32'h0000_0004 ? add_82190 : array_index_82184[4];
  assign array_update_82192[5] = add_82152 == 32'h0000_0005 ? add_82190 : array_index_82184[5];
  assign array_update_82192[6] = add_82152 == 32'h0000_0006 ? add_82190 : array_index_82184[6];
  assign array_update_82192[7] = add_82152 == 32'h0000_0007 ? add_82190 : array_index_82184[7];
  assign array_update_82192[8] = add_82152 == 32'h0000_0008 ? add_82190 : array_index_82184[8];
  assign array_update_82192[9] = add_82152 == 32'h0000_0009 ? add_82190 : array_index_82184[9];
  assign add_82193 = add_82180 + 32'h0000_0001;
  assign array_update_82194[0] = add_81474 == 32'h0000_0000 ? array_update_82192 : array_update_82181[0];
  assign array_update_82194[1] = add_81474 == 32'h0000_0001 ? array_update_82192 : array_update_82181[1];
  assign array_update_82194[2] = add_81474 == 32'h0000_0002 ? array_update_82192 : array_update_82181[2];
  assign array_update_82194[3] = add_81474 == 32'h0000_0003 ? array_update_82192 : array_update_82181[3];
  assign array_update_82194[4] = add_81474 == 32'h0000_0004 ? array_update_82192 : array_update_82181[4];
  assign array_update_82194[5] = add_81474 == 32'h0000_0005 ? array_update_82192 : array_update_82181[5];
  assign array_update_82194[6] = add_81474 == 32'h0000_0006 ? array_update_82192 : array_update_82181[6];
  assign array_update_82194[7] = add_81474 == 32'h0000_0007 ? array_update_82192 : array_update_82181[7];
  assign array_update_82194[8] = add_81474 == 32'h0000_0008 ? array_update_82192 : array_update_82181[8];
  assign array_update_82194[9] = add_81474 == 32'h0000_0009 ? array_update_82192 : array_update_82181[9];
  assign array_index_82196 = array_update_72021[add_82193 > 32'h0000_0009 ? 4'h9 : add_82193[3:0]];
  assign array_index_82197 = array_update_82194[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_82201 = smul32b_32b_x_32b(array_index_81481[add_82193 > 32'h0000_0009 ? 4'h9 : add_82193[3:0]], array_index_82196[add_82152 > 32'h0000_0009 ? 4'h9 : add_82152[3:0]]);
  assign add_82203 = array_index_82197[add_82152 > 32'h0000_0009 ? 4'h9 : add_82152[3:0]] + smul_82201;
  assign array_update_82205[0] = add_82152 == 32'h0000_0000 ? add_82203 : array_index_82197[0];
  assign array_update_82205[1] = add_82152 == 32'h0000_0001 ? add_82203 : array_index_82197[1];
  assign array_update_82205[2] = add_82152 == 32'h0000_0002 ? add_82203 : array_index_82197[2];
  assign array_update_82205[3] = add_82152 == 32'h0000_0003 ? add_82203 : array_index_82197[3];
  assign array_update_82205[4] = add_82152 == 32'h0000_0004 ? add_82203 : array_index_82197[4];
  assign array_update_82205[5] = add_82152 == 32'h0000_0005 ? add_82203 : array_index_82197[5];
  assign array_update_82205[6] = add_82152 == 32'h0000_0006 ? add_82203 : array_index_82197[6];
  assign array_update_82205[7] = add_82152 == 32'h0000_0007 ? add_82203 : array_index_82197[7];
  assign array_update_82205[8] = add_82152 == 32'h0000_0008 ? add_82203 : array_index_82197[8];
  assign array_update_82205[9] = add_82152 == 32'h0000_0009 ? add_82203 : array_index_82197[9];
  assign add_82206 = add_82193 + 32'h0000_0001;
  assign array_update_82207[0] = add_81474 == 32'h0000_0000 ? array_update_82205 : array_update_82194[0];
  assign array_update_82207[1] = add_81474 == 32'h0000_0001 ? array_update_82205 : array_update_82194[1];
  assign array_update_82207[2] = add_81474 == 32'h0000_0002 ? array_update_82205 : array_update_82194[2];
  assign array_update_82207[3] = add_81474 == 32'h0000_0003 ? array_update_82205 : array_update_82194[3];
  assign array_update_82207[4] = add_81474 == 32'h0000_0004 ? array_update_82205 : array_update_82194[4];
  assign array_update_82207[5] = add_81474 == 32'h0000_0005 ? array_update_82205 : array_update_82194[5];
  assign array_update_82207[6] = add_81474 == 32'h0000_0006 ? array_update_82205 : array_update_82194[6];
  assign array_update_82207[7] = add_81474 == 32'h0000_0007 ? array_update_82205 : array_update_82194[7];
  assign array_update_82207[8] = add_81474 == 32'h0000_0008 ? array_update_82205 : array_update_82194[8];
  assign array_update_82207[9] = add_81474 == 32'h0000_0009 ? array_update_82205 : array_update_82194[9];
  assign array_index_82209 = array_update_72021[add_82206 > 32'h0000_0009 ? 4'h9 : add_82206[3:0]];
  assign array_index_82210 = array_update_82207[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_82214 = smul32b_32b_x_32b(array_index_81481[add_82206 > 32'h0000_0009 ? 4'h9 : add_82206[3:0]], array_index_82209[add_82152 > 32'h0000_0009 ? 4'h9 : add_82152[3:0]]);
  assign add_82216 = array_index_82210[add_82152 > 32'h0000_0009 ? 4'h9 : add_82152[3:0]] + smul_82214;
  assign array_update_82218[0] = add_82152 == 32'h0000_0000 ? add_82216 : array_index_82210[0];
  assign array_update_82218[1] = add_82152 == 32'h0000_0001 ? add_82216 : array_index_82210[1];
  assign array_update_82218[2] = add_82152 == 32'h0000_0002 ? add_82216 : array_index_82210[2];
  assign array_update_82218[3] = add_82152 == 32'h0000_0003 ? add_82216 : array_index_82210[3];
  assign array_update_82218[4] = add_82152 == 32'h0000_0004 ? add_82216 : array_index_82210[4];
  assign array_update_82218[5] = add_82152 == 32'h0000_0005 ? add_82216 : array_index_82210[5];
  assign array_update_82218[6] = add_82152 == 32'h0000_0006 ? add_82216 : array_index_82210[6];
  assign array_update_82218[7] = add_82152 == 32'h0000_0007 ? add_82216 : array_index_82210[7];
  assign array_update_82218[8] = add_82152 == 32'h0000_0008 ? add_82216 : array_index_82210[8];
  assign array_update_82218[9] = add_82152 == 32'h0000_0009 ? add_82216 : array_index_82210[9];
  assign add_82219 = add_82206 + 32'h0000_0001;
  assign array_update_82220[0] = add_81474 == 32'h0000_0000 ? array_update_82218 : array_update_82207[0];
  assign array_update_82220[1] = add_81474 == 32'h0000_0001 ? array_update_82218 : array_update_82207[1];
  assign array_update_82220[2] = add_81474 == 32'h0000_0002 ? array_update_82218 : array_update_82207[2];
  assign array_update_82220[3] = add_81474 == 32'h0000_0003 ? array_update_82218 : array_update_82207[3];
  assign array_update_82220[4] = add_81474 == 32'h0000_0004 ? array_update_82218 : array_update_82207[4];
  assign array_update_82220[5] = add_81474 == 32'h0000_0005 ? array_update_82218 : array_update_82207[5];
  assign array_update_82220[6] = add_81474 == 32'h0000_0006 ? array_update_82218 : array_update_82207[6];
  assign array_update_82220[7] = add_81474 == 32'h0000_0007 ? array_update_82218 : array_update_82207[7];
  assign array_update_82220[8] = add_81474 == 32'h0000_0008 ? array_update_82218 : array_update_82207[8];
  assign array_update_82220[9] = add_81474 == 32'h0000_0009 ? array_update_82218 : array_update_82207[9];
  assign array_index_82222 = array_update_72021[add_82219 > 32'h0000_0009 ? 4'h9 : add_82219[3:0]];
  assign array_index_82223 = array_update_82220[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_82227 = smul32b_32b_x_32b(array_index_81481[add_82219 > 32'h0000_0009 ? 4'h9 : add_82219[3:0]], array_index_82222[add_82152 > 32'h0000_0009 ? 4'h9 : add_82152[3:0]]);
  assign add_82229 = array_index_82223[add_82152 > 32'h0000_0009 ? 4'h9 : add_82152[3:0]] + smul_82227;
  assign array_update_82231[0] = add_82152 == 32'h0000_0000 ? add_82229 : array_index_82223[0];
  assign array_update_82231[1] = add_82152 == 32'h0000_0001 ? add_82229 : array_index_82223[1];
  assign array_update_82231[2] = add_82152 == 32'h0000_0002 ? add_82229 : array_index_82223[2];
  assign array_update_82231[3] = add_82152 == 32'h0000_0003 ? add_82229 : array_index_82223[3];
  assign array_update_82231[4] = add_82152 == 32'h0000_0004 ? add_82229 : array_index_82223[4];
  assign array_update_82231[5] = add_82152 == 32'h0000_0005 ? add_82229 : array_index_82223[5];
  assign array_update_82231[6] = add_82152 == 32'h0000_0006 ? add_82229 : array_index_82223[6];
  assign array_update_82231[7] = add_82152 == 32'h0000_0007 ? add_82229 : array_index_82223[7];
  assign array_update_82231[8] = add_82152 == 32'h0000_0008 ? add_82229 : array_index_82223[8];
  assign array_update_82231[9] = add_82152 == 32'h0000_0009 ? add_82229 : array_index_82223[9];
  assign add_82232 = add_82219 + 32'h0000_0001;
  assign array_update_82233[0] = add_81474 == 32'h0000_0000 ? array_update_82231 : array_update_82220[0];
  assign array_update_82233[1] = add_81474 == 32'h0000_0001 ? array_update_82231 : array_update_82220[1];
  assign array_update_82233[2] = add_81474 == 32'h0000_0002 ? array_update_82231 : array_update_82220[2];
  assign array_update_82233[3] = add_81474 == 32'h0000_0003 ? array_update_82231 : array_update_82220[3];
  assign array_update_82233[4] = add_81474 == 32'h0000_0004 ? array_update_82231 : array_update_82220[4];
  assign array_update_82233[5] = add_81474 == 32'h0000_0005 ? array_update_82231 : array_update_82220[5];
  assign array_update_82233[6] = add_81474 == 32'h0000_0006 ? array_update_82231 : array_update_82220[6];
  assign array_update_82233[7] = add_81474 == 32'h0000_0007 ? array_update_82231 : array_update_82220[7];
  assign array_update_82233[8] = add_81474 == 32'h0000_0008 ? array_update_82231 : array_update_82220[8];
  assign array_update_82233[9] = add_81474 == 32'h0000_0009 ? array_update_82231 : array_update_82220[9];
  assign array_index_82235 = array_update_72021[add_82232 > 32'h0000_0009 ? 4'h9 : add_82232[3:0]];
  assign array_index_82236 = array_update_82233[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_82240 = smul32b_32b_x_32b(array_index_81481[add_82232 > 32'h0000_0009 ? 4'h9 : add_82232[3:0]], array_index_82235[add_82152 > 32'h0000_0009 ? 4'h9 : add_82152[3:0]]);
  assign add_82242 = array_index_82236[add_82152 > 32'h0000_0009 ? 4'h9 : add_82152[3:0]] + smul_82240;
  assign array_update_82244[0] = add_82152 == 32'h0000_0000 ? add_82242 : array_index_82236[0];
  assign array_update_82244[1] = add_82152 == 32'h0000_0001 ? add_82242 : array_index_82236[1];
  assign array_update_82244[2] = add_82152 == 32'h0000_0002 ? add_82242 : array_index_82236[2];
  assign array_update_82244[3] = add_82152 == 32'h0000_0003 ? add_82242 : array_index_82236[3];
  assign array_update_82244[4] = add_82152 == 32'h0000_0004 ? add_82242 : array_index_82236[4];
  assign array_update_82244[5] = add_82152 == 32'h0000_0005 ? add_82242 : array_index_82236[5];
  assign array_update_82244[6] = add_82152 == 32'h0000_0006 ? add_82242 : array_index_82236[6];
  assign array_update_82244[7] = add_82152 == 32'h0000_0007 ? add_82242 : array_index_82236[7];
  assign array_update_82244[8] = add_82152 == 32'h0000_0008 ? add_82242 : array_index_82236[8];
  assign array_update_82244[9] = add_82152 == 32'h0000_0009 ? add_82242 : array_index_82236[9];
  assign add_82245 = add_82232 + 32'h0000_0001;
  assign array_update_82246[0] = add_81474 == 32'h0000_0000 ? array_update_82244 : array_update_82233[0];
  assign array_update_82246[1] = add_81474 == 32'h0000_0001 ? array_update_82244 : array_update_82233[1];
  assign array_update_82246[2] = add_81474 == 32'h0000_0002 ? array_update_82244 : array_update_82233[2];
  assign array_update_82246[3] = add_81474 == 32'h0000_0003 ? array_update_82244 : array_update_82233[3];
  assign array_update_82246[4] = add_81474 == 32'h0000_0004 ? array_update_82244 : array_update_82233[4];
  assign array_update_82246[5] = add_81474 == 32'h0000_0005 ? array_update_82244 : array_update_82233[5];
  assign array_update_82246[6] = add_81474 == 32'h0000_0006 ? array_update_82244 : array_update_82233[6];
  assign array_update_82246[7] = add_81474 == 32'h0000_0007 ? array_update_82244 : array_update_82233[7];
  assign array_update_82246[8] = add_81474 == 32'h0000_0008 ? array_update_82244 : array_update_82233[8];
  assign array_update_82246[9] = add_81474 == 32'h0000_0009 ? array_update_82244 : array_update_82233[9];
  assign array_index_82248 = array_update_72021[add_82245 > 32'h0000_0009 ? 4'h9 : add_82245[3:0]];
  assign array_index_82249 = array_update_82246[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_82253 = smul32b_32b_x_32b(array_index_81481[add_82245 > 32'h0000_0009 ? 4'h9 : add_82245[3:0]], array_index_82248[add_82152 > 32'h0000_0009 ? 4'h9 : add_82152[3:0]]);
  assign add_82255 = array_index_82249[add_82152 > 32'h0000_0009 ? 4'h9 : add_82152[3:0]] + smul_82253;
  assign array_update_82257[0] = add_82152 == 32'h0000_0000 ? add_82255 : array_index_82249[0];
  assign array_update_82257[1] = add_82152 == 32'h0000_0001 ? add_82255 : array_index_82249[1];
  assign array_update_82257[2] = add_82152 == 32'h0000_0002 ? add_82255 : array_index_82249[2];
  assign array_update_82257[3] = add_82152 == 32'h0000_0003 ? add_82255 : array_index_82249[3];
  assign array_update_82257[4] = add_82152 == 32'h0000_0004 ? add_82255 : array_index_82249[4];
  assign array_update_82257[5] = add_82152 == 32'h0000_0005 ? add_82255 : array_index_82249[5];
  assign array_update_82257[6] = add_82152 == 32'h0000_0006 ? add_82255 : array_index_82249[6];
  assign array_update_82257[7] = add_82152 == 32'h0000_0007 ? add_82255 : array_index_82249[7];
  assign array_update_82257[8] = add_82152 == 32'h0000_0008 ? add_82255 : array_index_82249[8];
  assign array_update_82257[9] = add_82152 == 32'h0000_0009 ? add_82255 : array_index_82249[9];
  assign add_82258 = add_82245 + 32'h0000_0001;
  assign array_update_82259[0] = add_81474 == 32'h0000_0000 ? array_update_82257 : array_update_82246[0];
  assign array_update_82259[1] = add_81474 == 32'h0000_0001 ? array_update_82257 : array_update_82246[1];
  assign array_update_82259[2] = add_81474 == 32'h0000_0002 ? array_update_82257 : array_update_82246[2];
  assign array_update_82259[3] = add_81474 == 32'h0000_0003 ? array_update_82257 : array_update_82246[3];
  assign array_update_82259[4] = add_81474 == 32'h0000_0004 ? array_update_82257 : array_update_82246[4];
  assign array_update_82259[5] = add_81474 == 32'h0000_0005 ? array_update_82257 : array_update_82246[5];
  assign array_update_82259[6] = add_81474 == 32'h0000_0006 ? array_update_82257 : array_update_82246[6];
  assign array_update_82259[7] = add_81474 == 32'h0000_0007 ? array_update_82257 : array_update_82246[7];
  assign array_update_82259[8] = add_81474 == 32'h0000_0008 ? array_update_82257 : array_update_82246[8];
  assign array_update_82259[9] = add_81474 == 32'h0000_0009 ? array_update_82257 : array_update_82246[9];
  assign array_index_82261 = array_update_72021[add_82258 > 32'h0000_0009 ? 4'h9 : add_82258[3:0]];
  assign array_index_82262 = array_update_82259[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_82266 = smul32b_32b_x_32b(array_index_81481[add_82258 > 32'h0000_0009 ? 4'h9 : add_82258[3:0]], array_index_82261[add_82152 > 32'h0000_0009 ? 4'h9 : add_82152[3:0]]);
  assign add_82268 = array_index_82262[add_82152 > 32'h0000_0009 ? 4'h9 : add_82152[3:0]] + smul_82266;
  assign array_update_82270[0] = add_82152 == 32'h0000_0000 ? add_82268 : array_index_82262[0];
  assign array_update_82270[1] = add_82152 == 32'h0000_0001 ? add_82268 : array_index_82262[1];
  assign array_update_82270[2] = add_82152 == 32'h0000_0002 ? add_82268 : array_index_82262[2];
  assign array_update_82270[3] = add_82152 == 32'h0000_0003 ? add_82268 : array_index_82262[3];
  assign array_update_82270[4] = add_82152 == 32'h0000_0004 ? add_82268 : array_index_82262[4];
  assign array_update_82270[5] = add_82152 == 32'h0000_0005 ? add_82268 : array_index_82262[5];
  assign array_update_82270[6] = add_82152 == 32'h0000_0006 ? add_82268 : array_index_82262[6];
  assign array_update_82270[7] = add_82152 == 32'h0000_0007 ? add_82268 : array_index_82262[7];
  assign array_update_82270[8] = add_82152 == 32'h0000_0008 ? add_82268 : array_index_82262[8];
  assign array_update_82270[9] = add_82152 == 32'h0000_0009 ? add_82268 : array_index_82262[9];
  assign add_82271 = add_82258 + 32'h0000_0001;
  assign array_update_82272[0] = add_81474 == 32'h0000_0000 ? array_update_82270 : array_update_82259[0];
  assign array_update_82272[1] = add_81474 == 32'h0000_0001 ? array_update_82270 : array_update_82259[1];
  assign array_update_82272[2] = add_81474 == 32'h0000_0002 ? array_update_82270 : array_update_82259[2];
  assign array_update_82272[3] = add_81474 == 32'h0000_0003 ? array_update_82270 : array_update_82259[3];
  assign array_update_82272[4] = add_81474 == 32'h0000_0004 ? array_update_82270 : array_update_82259[4];
  assign array_update_82272[5] = add_81474 == 32'h0000_0005 ? array_update_82270 : array_update_82259[5];
  assign array_update_82272[6] = add_81474 == 32'h0000_0006 ? array_update_82270 : array_update_82259[6];
  assign array_update_82272[7] = add_81474 == 32'h0000_0007 ? array_update_82270 : array_update_82259[7];
  assign array_update_82272[8] = add_81474 == 32'h0000_0008 ? array_update_82270 : array_update_82259[8];
  assign array_update_82272[9] = add_81474 == 32'h0000_0009 ? array_update_82270 : array_update_82259[9];
  assign array_index_82274 = array_update_72021[add_82271 > 32'h0000_0009 ? 4'h9 : add_82271[3:0]];
  assign array_index_82275 = array_update_82272[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_82279 = smul32b_32b_x_32b(array_index_81481[add_82271 > 32'h0000_0009 ? 4'h9 : add_82271[3:0]], array_index_82274[add_82152 > 32'h0000_0009 ? 4'h9 : add_82152[3:0]]);
  assign add_82281 = array_index_82275[add_82152 > 32'h0000_0009 ? 4'h9 : add_82152[3:0]] + smul_82279;
  assign array_update_82282[0] = add_82152 == 32'h0000_0000 ? add_82281 : array_index_82275[0];
  assign array_update_82282[1] = add_82152 == 32'h0000_0001 ? add_82281 : array_index_82275[1];
  assign array_update_82282[2] = add_82152 == 32'h0000_0002 ? add_82281 : array_index_82275[2];
  assign array_update_82282[3] = add_82152 == 32'h0000_0003 ? add_82281 : array_index_82275[3];
  assign array_update_82282[4] = add_82152 == 32'h0000_0004 ? add_82281 : array_index_82275[4];
  assign array_update_82282[5] = add_82152 == 32'h0000_0005 ? add_82281 : array_index_82275[5];
  assign array_update_82282[6] = add_82152 == 32'h0000_0006 ? add_82281 : array_index_82275[6];
  assign array_update_82282[7] = add_82152 == 32'h0000_0007 ? add_82281 : array_index_82275[7];
  assign array_update_82282[8] = add_82152 == 32'h0000_0008 ? add_82281 : array_index_82275[8];
  assign array_update_82282[9] = add_82152 == 32'h0000_0009 ? add_82281 : array_index_82275[9];
  assign array_update_82283[0] = add_81474 == 32'h0000_0000 ? array_update_82282 : array_update_82272[0];
  assign array_update_82283[1] = add_81474 == 32'h0000_0001 ? array_update_82282 : array_update_82272[1];
  assign array_update_82283[2] = add_81474 == 32'h0000_0002 ? array_update_82282 : array_update_82272[2];
  assign array_update_82283[3] = add_81474 == 32'h0000_0003 ? array_update_82282 : array_update_82272[3];
  assign array_update_82283[4] = add_81474 == 32'h0000_0004 ? array_update_82282 : array_update_82272[4];
  assign array_update_82283[5] = add_81474 == 32'h0000_0005 ? array_update_82282 : array_update_82272[5];
  assign array_update_82283[6] = add_81474 == 32'h0000_0006 ? array_update_82282 : array_update_82272[6];
  assign array_update_82283[7] = add_81474 == 32'h0000_0007 ? array_update_82282 : array_update_82272[7];
  assign array_update_82283[8] = add_81474 == 32'h0000_0008 ? array_update_82282 : array_update_82272[8];
  assign array_update_82283[9] = add_81474 == 32'h0000_0009 ? array_update_82282 : array_update_82272[9];
  assign array_index_82285 = array_update_82283[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign add_82287 = add_82152 + 32'h0000_0001;
  assign array_update_82288[0] = add_82287 == 32'h0000_0000 ? 32'h0000_0000 : array_index_82285[0];
  assign array_update_82288[1] = add_82287 == 32'h0000_0001 ? 32'h0000_0000 : array_index_82285[1];
  assign array_update_82288[2] = add_82287 == 32'h0000_0002 ? 32'h0000_0000 : array_index_82285[2];
  assign array_update_82288[3] = add_82287 == 32'h0000_0003 ? 32'h0000_0000 : array_index_82285[3];
  assign array_update_82288[4] = add_82287 == 32'h0000_0004 ? 32'h0000_0000 : array_index_82285[4];
  assign array_update_82288[5] = add_82287 == 32'h0000_0005 ? 32'h0000_0000 : array_index_82285[5];
  assign array_update_82288[6] = add_82287 == 32'h0000_0006 ? 32'h0000_0000 : array_index_82285[6];
  assign array_update_82288[7] = add_82287 == 32'h0000_0007 ? 32'h0000_0000 : array_index_82285[7];
  assign array_update_82288[8] = add_82287 == 32'h0000_0008 ? 32'h0000_0000 : array_index_82285[8];
  assign array_update_82288[9] = add_82287 == 32'h0000_0009 ? 32'h0000_0000 : array_index_82285[9];
  assign literal_82289 = 32'h0000_0000;
  assign array_update_82290[0] = add_81474 == 32'h0000_0000 ? array_update_82288 : array_update_82283[0];
  assign array_update_82290[1] = add_81474 == 32'h0000_0001 ? array_update_82288 : array_update_82283[1];
  assign array_update_82290[2] = add_81474 == 32'h0000_0002 ? array_update_82288 : array_update_82283[2];
  assign array_update_82290[3] = add_81474 == 32'h0000_0003 ? array_update_82288 : array_update_82283[3];
  assign array_update_82290[4] = add_81474 == 32'h0000_0004 ? array_update_82288 : array_update_82283[4];
  assign array_update_82290[5] = add_81474 == 32'h0000_0005 ? array_update_82288 : array_update_82283[5];
  assign array_update_82290[6] = add_81474 == 32'h0000_0006 ? array_update_82288 : array_update_82283[6];
  assign array_update_82290[7] = add_81474 == 32'h0000_0007 ? array_update_82288 : array_update_82283[7];
  assign array_update_82290[8] = add_81474 == 32'h0000_0008 ? array_update_82288 : array_update_82283[8];
  assign array_update_82290[9] = add_81474 == 32'h0000_0009 ? array_update_82288 : array_update_82283[9];
  assign array_index_82292 = array_update_72021[literal_82289 > 32'h0000_0009 ? 4'h9 : literal_82289[3:0]];
  assign array_index_82293 = array_update_82290[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_82297 = smul32b_32b_x_32b(array_index_81481[literal_82289 > 32'h0000_0009 ? 4'h9 : literal_82289[3:0]], array_index_82292[add_82287 > 32'h0000_0009 ? 4'h9 : add_82287[3:0]]);
  assign add_82299 = array_index_82293[add_82287 > 32'h0000_0009 ? 4'h9 : add_82287[3:0]] + smul_82297;
  assign array_update_82301[0] = add_82287 == 32'h0000_0000 ? add_82299 : array_index_82293[0];
  assign array_update_82301[1] = add_82287 == 32'h0000_0001 ? add_82299 : array_index_82293[1];
  assign array_update_82301[2] = add_82287 == 32'h0000_0002 ? add_82299 : array_index_82293[2];
  assign array_update_82301[3] = add_82287 == 32'h0000_0003 ? add_82299 : array_index_82293[3];
  assign array_update_82301[4] = add_82287 == 32'h0000_0004 ? add_82299 : array_index_82293[4];
  assign array_update_82301[5] = add_82287 == 32'h0000_0005 ? add_82299 : array_index_82293[5];
  assign array_update_82301[6] = add_82287 == 32'h0000_0006 ? add_82299 : array_index_82293[6];
  assign array_update_82301[7] = add_82287 == 32'h0000_0007 ? add_82299 : array_index_82293[7];
  assign array_update_82301[8] = add_82287 == 32'h0000_0008 ? add_82299 : array_index_82293[8];
  assign array_update_82301[9] = add_82287 == 32'h0000_0009 ? add_82299 : array_index_82293[9];
  assign add_82302 = literal_82289 + 32'h0000_0001;
  assign array_update_82303[0] = add_81474 == 32'h0000_0000 ? array_update_82301 : array_update_82290[0];
  assign array_update_82303[1] = add_81474 == 32'h0000_0001 ? array_update_82301 : array_update_82290[1];
  assign array_update_82303[2] = add_81474 == 32'h0000_0002 ? array_update_82301 : array_update_82290[2];
  assign array_update_82303[3] = add_81474 == 32'h0000_0003 ? array_update_82301 : array_update_82290[3];
  assign array_update_82303[4] = add_81474 == 32'h0000_0004 ? array_update_82301 : array_update_82290[4];
  assign array_update_82303[5] = add_81474 == 32'h0000_0005 ? array_update_82301 : array_update_82290[5];
  assign array_update_82303[6] = add_81474 == 32'h0000_0006 ? array_update_82301 : array_update_82290[6];
  assign array_update_82303[7] = add_81474 == 32'h0000_0007 ? array_update_82301 : array_update_82290[7];
  assign array_update_82303[8] = add_81474 == 32'h0000_0008 ? array_update_82301 : array_update_82290[8];
  assign array_update_82303[9] = add_81474 == 32'h0000_0009 ? array_update_82301 : array_update_82290[9];
  assign array_index_82305 = array_update_72021[add_82302 > 32'h0000_0009 ? 4'h9 : add_82302[3:0]];
  assign array_index_82306 = array_update_82303[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_82310 = smul32b_32b_x_32b(array_index_81481[add_82302 > 32'h0000_0009 ? 4'h9 : add_82302[3:0]], array_index_82305[add_82287 > 32'h0000_0009 ? 4'h9 : add_82287[3:0]]);
  assign add_82312 = array_index_82306[add_82287 > 32'h0000_0009 ? 4'h9 : add_82287[3:0]] + smul_82310;
  assign array_update_82314[0] = add_82287 == 32'h0000_0000 ? add_82312 : array_index_82306[0];
  assign array_update_82314[1] = add_82287 == 32'h0000_0001 ? add_82312 : array_index_82306[1];
  assign array_update_82314[2] = add_82287 == 32'h0000_0002 ? add_82312 : array_index_82306[2];
  assign array_update_82314[3] = add_82287 == 32'h0000_0003 ? add_82312 : array_index_82306[3];
  assign array_update_82314[4] = add_82287 == 32'h0000_0004 ? add_82312 : array_index_82306[4];
  assign array_update_82314[5] = add_82287 == 32'h0000_0005 ? add_82312 : array_index_82306[5];
  assign array_update_82314[6] = add_82287 == 32'h0000_0006 ? add_82312 : array_index_82306[6];
  assign array_update_82314[7] = add_82287 == 32'h0000_0007 ? add_82312 : array_index_82306[7];
  assign array_update_82314[8] = add_82287 == 32'h0000_0008 ? add_82312 : array_index_82306[8];
  assign array_update_82314[9] = add_82287 == 32'h0000_0009 ? add_82312 : array_index_82306[9];
  assign add_82315 = add_82302 + 32'h0000_0001;
  assign array_update_82316[0] = add_81474 == 32'h0000_0000 ? array_update_82314 : array_update_82303[0];
  assign array_update_82316[1] = add_81474 == 32'h0000_0001 ? array_update_82314 : array_update_82303[1];
  assign array_update_82316[2] = add_81474 == 32'h0000_0002 ? array_update_82314 : array_update_82303[2];
  assign array_update_82316[3] = add_81474 == 32'h0000_0003 ? array_update_82314 : array_update_82303[3];
  assign array_update_82316[4] = add_81474 == 32'h0000_0004 ? array_update_82314 : array_update_82303[4];
  assign array_update_82316[5] = add_81474 == 32'h0000_0005 ? array_update_82314 : array_update_82303[5];
  assign array_update_82316[6] = add_81474 == 32'h0000_0006 ? array_update_82314 : array_update_82303[6];
  assign array_update_82316[7] = add_81474 == 32'h0000_0007 ? array_update_82314 : array_update_82303[7];
  assign array_update_82316[8] = add_81474 == 32'h0000_0008 ? array_update_82314 : array_update_82303[8];
  assign array_update_82316[9] = add_81474 == 32'h0000_0009 ? array_update_82314 : array_update_82303[9];
  assign array_index_82318 = array_update_72021[add_82315 > 32'h0000_0009 ? 4'h9 : add_82315[3:0]];
  assign array_index_82319 = array_update_82316[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_82323 = smul32b_32b_x_32b(array_index_81481[add_82315 > 32'h0000_0009 ? 4'h9 : add_82315[3:0]], array_index_82318[add_82287 > 32'h0000_0009 ? 4'h9 : add_82287[3:0]]);
  assign add_82325 = array_index_82319[add_82287 > 32'h0000_0009 ? 4'h9 : add_82287[3:0]] + smul_82323;
  assign array_update_82327[0] = add_82287 == 32'h0000_0000 ? add_82325 : array_index_82319[0];
  assign array_update_82327[1] = add_82287 == 32'h0000_0001 ? add_82325 : array_index_82319[1];
  assign array_update_82327[2] = add_82287 == 32'h0000_0002 ? add_82325 : array_index_82319[2];
  assign array_update_82327[3] = add_82287 == 32'h0000_0003 ? add_82325 : array_index_82319[3];
  assign array_update_82327[4] = add_82287 == 32'h0000_0004 ? add_82325 : array_index_82319[4];
  assign array_update_82327[5] = add_82287 == 32'h0000_0005 ? add_82325 : array_index_82319[5];
  assign array_update_82327[6] = add_82287 == 32'h0000_0006 ? add_82325 : array_index_82319[6];
  assign array_update_82327[7] = add_82287 == 32'h0000_0007 ? add_82325 : array_index_82319[7];
  assign array_update_82327[8] = add_82287 == 32'h0000_0008 ? add_82325 : array_index_82319[8];
  assign array_update_82327[9] = add_82287 == 32'h0000_0009 ? add_82325 : array_index_82319[9];
  assign add_82328 = add_82315 + 32'h0000_0001;
  assign array_update_82329[0] = add_81474 == 32'h0000_0000 ? array_update_82327 : array_update_82316[0];
  assign array_update_82329[1] = add_81474 == 32'h0000_0001 ? array_update_82327 : array_update_82316[1];
  assign array_update_82329[2] = add_81474 == 32'h0000_0002 ? array_update_82327 : array_update_82316[2];
  assign array_update_82329[3] = add_81474 == 32'h0000_0003 ? array_update_82327 : array_update_82316[3];
  assign array_update_82329[4] = add_81474 == 32'h0000_0004 ? array_update_82327 : array_update_82316[4];
  assign array_update_82329[5] = add_81474 == 32'h0000_0005 ? array_update_82327 : array_update_82316[5];
  assign array_update_82329[6] = add_81474 == 32'h0000_0006 ? array_update_82327 : array_update_82316[6];
  assign array_update_82329[7] = add_81474 == 32'h0000_0007 ? array_update_82327 : array_update_82316[7];
  assign array_update_82329[8] = add_81474 == 32'h0000_0008 ? array_update_82327 : array_update_82316[8];
  assign array_update_82329[9] = add_81474 == 32'h0000_0009 ? array_update_82327 : array_update_82316[9];
  assign array_index_82331 = array_update_72021[add_82328 > 32'h0000_0009 ? 4'h9 : add_82328[3:0]];
  assign array_index_82332 = array_update_82329[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_82336 = smul32b_32b_x_32b(array_index_81481[add_82328 > 32'h0000_0009 ? 4'h9 : add_82328[3:0]], array_index_82331[add_82287 > 32'h0000_0009 ? 4'h9 : add_82287[3:0]]);
  assign add_82338 = array_index_82332[add_82287 > 32'h0000_0009 ? 4'h9 : add_82287[3:0]] + smul_82336;
  assign array_update_82340[0] = add_82287 == 32'h0000_0000 ? add_82338 : array_index_82332[0];
  assign array_update_82340[1] = add_82287 == 32'h0000_0001 ? add_82338 : array_index_82332[1];
  assign array_update_82340[2] = add_82287 == 32'h0000_0002 ? add_82338 : array_index_82332[2];
  assign array_update_82340[3] = add_82287 == 32'h0000_0003 ? add_82338 : array_index_82332[3];
  assign array_update_82340[4] = add_82287 == 32'h0000_0004 ? add_82338 : array_index_82332[4];
  assign array_update_82340[5] = add_82287 == 32'h0000_0005 ? add_82338 : array_index_82332[5];
  assign array_update_82340[6] = add_82287 == 32'h0000_0006 ? add_82338 : array_index_82332[6];
  assign array_update_82340[7] = add_82287 == 32'h0000_0007 ? add_82338 : array_index_82332[7];
  assign array_update_82340[8] = add_82287 == 32'h0000_0008 ? add_82338 : array_index_82332[8];
  assign array_update_82340[9] = add_82287 == 32'h0000_0009 ? add_82338 : array_index_82332[9];
  assign add_82341 = add_82328 + 32'h0000_0001;
  assign array_update_82342[0] = add_81474 == 32'h0000_0000 ? array_update_82340 : array_update_82329[0];
  assign array_update_82342[1] = add_81474 == 32'h0000_0001 ? array_update_82340 : array_update_82329[1];
  assign array_update_82342[2] = add_81474 == 32'h0000_0002 ? array_update_82340 : array_update_82329[2];
  assign array_update_82342[3] = add_81474 == 32'h0000_0003 ? array_update_82340 : array_update_82329[3];
  assign array_update_82342[4] = add_81474 == 32'h0000_0004 ? array_update_82340 : array_update_82329[4];
  assign array_update_82342[5] = add_81474 == 32'h0000_0005 ? array_update_82340 : array_update_82329[5];
  assign array_update_82342[6] = add_81474 == 32'h0000_0006 ? array_update_82340 : array_update_82329[6];
  assign array_update_82342[7] = add_81474 == 32'h0000_0007 ? array_update_82340 : array_update_82329[7];
  assign array_update_82342[8] = add_81474 == 32'h0000_0008 ? array_update_82340 : array_update_82329[8];
  assign array_update_82342[9] = add_81474 == 32'h0000_0009 ? array_update_82340 : array_update_82329[9];
  assign array_index_82344 = array_update_72021[add_82341 > 32'h0000_0009 ? 4'h9 : add_82341[3:0]];
  assign array_index_82345 = array_update_82342[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_82349 = smul32b_32b_x_32b(array_index_81481[add_82341 > 32'h0000_0009 ? 4'h9 : add_82341[3:0]], array_index_82344[add_82287 > 32'h0000_0009 ? 4'h9 : add_82287[3:0]]);
  assign add_82351 = array_index_82345[add_82287 > 32'h0000_0009 ? 4'h9 : add_82287[3:0]] + smul_82349;
  assign array_update_82353[0] = add_82287 == 32'h0000_0000 ? add_82351 : array_index_82345[0];
  assign array_update_82353[1] = add_82287 == 32'h0000_0001 ? add_82351 : array_index_82345[1];
  assign array_update_82353[2] = add_82287 == 32'h0000_0002 ? add_82351 : array_index_82345[2];
  assign array_update_82353[3] = add_82287 == 32'h0000_0003 ? add_82351 : array_index_82345[3];
  assign array_update_82353[4] = add_82287 == 32'h0000_0004 ? add_82351 : array_index_82345[4];
  assign array_update_82353[5] = add_82287 == 32'h0000_0005 ? add_82351 : array_index_82345[5];
  assign array_update_82353[6] = add_82287 == 32'h0000_0006 ? add_82351 : array_index_82345[6];
  assign array_update_82353[7] = add_82287 == 32'h0000_0007 ? add_82351 : array_index_82345[7];
  assign array_update_82353[8] = add_82287 == 32'h0000_0008 ? add_82351 : array_index_82345[8];
  assign array_update_82353[9] = add_82287 == 32'h0000_0009 ? add_82351 : array_index_82345[9];
  assign add_82354 = add_82341 + 32'h0000_0001;
  assign array_update_82355[0] = add_81474 == 32'h0000_0000 ? array_update_82353 : array_update_82342[0];
  assign array_update_82355[1] = add_81474 == 32'h0000_0001 ? array_update_82353 : array_update_82342[1];
  assign array_update_82355[2] = add_81474 == 32'h0000_0002 ? array_update_82353 : array_update_82342[2];
  assign array_update_82355[3] = add_81474 == 32'h0000_0003 ? array_update_82353 : array_update_82342[3];
  assign array_update_82355[4] = add_81474 == 32'h0000_0004 ? array_update_82353 : array_update_82342[4];
  assign array_update_82355[5] = add_81474 == 32'h0000_0005 ? array_update_82353 : array_update_82342[5];
  assign array_update_82355[6] = add_81474 == 32'h0000_0006 ? array_update_82353 : array_update_82342[6];
  assign array_update_82355[7] = add_81474 == 32'h0000_0007 ? array_update_82353 : array_update_82342[7];
  assign array_update_82355[8] = add_81474 == 32'h0000_0008 ? array_update_82353 : array_update_82342[8];
  assign array_update_82355[9] = add_81474 == 32'h0000_0009 ? array_update_82353 : array_update_82342[9];
  assign array_index_82357 = array_update_72021[add_82354 > 32'h0000_0009 ? 4'h9 : add_82354[3:0]];
  assign array_index_82358 = array_update_82355[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_82362 = smul32b_32b_x_32b(array_index_81481[add_82354 > 32'h0000_0009 ? 4'h9 : add_82354[3:0]], array_index_82357[add_82287 > 32'h0000_0009 ? 4'h9 : add_82287[3:0]]);
  assign add_82364 = array_index_82358[add_82287 > 32'h0000_0009 ? 4'h9 : add_82287[3:0]] + smul_82362;
  assign array_update_82366[0] = add_82287 == 32'h0000_0000 ? add_82364 : array_index_82358[0];
  assign array_update_82366[1] = add_82287 == 32'h0000_0001 ? add_82364 : array_index_82358[1];
  assign array_update_82366[2] = add_82287 == 32'h0000_0002 ? add_82364 : array_index_82358[2];
  assign array_update_82366[3] = add_82287 == 32'h0000_0003 ? add_82364 : array_index_82358[3];
  assign array_update_82366[4] = add_82287 == 32'h0000_0004 ? add_82364 : array_index_82358[4];
  assign array_update_82366[5] = add_82287 == 32'h0000_0005 ? add_82364 : array_index_82358[5];
  assign array_update_82366[6] = add_82287 == 32'h0000_0006 ? add_82364 : array_index_82358[6];
  assign array_update_82366[7] = add_82287 == 32'h0000_0007 ? add_82364 : array_index_82358[7];
  assign array_update_82366[8] = add_82287 == 32'h0000_0008 ? add_82364 : array_index_82358[8];
  assign array_update_82366[9] = add_82287 == 32'h0000_0009 ? add_82364 : array_index_82358[9];
  assign add_82367 = add_82354 + 32'h0000_0001;
  assign array_update_82368[0] = add_81474 == 32'h0000_0000 ? array_update_82366 : array_update_82355[0];
  assign array_update_82368[1] = add_81474 == 32'h0000_0001 ? array_update_82366 : array_update_82355[1];
  assign array_update_82368[2] = add_81474 == 32'h0000_0002 ? array_update_82366 : array_update_82355[2];
  assign array_update_82368[3] = add_81474 == 32'h0000_0003 ? array_update_82366 : array_update_82355[3];
  assign array_update_82368[4] = add_81474 == 32'h0000_0004 ? array_update_82366 : array_update_82355[4];
  assign array_update_82368[5] = add_81474 == 32'h0000_0005 ? array_update_82366 : array_update_82355[5];
  assign array_update_82368[6] = add_81474 == 32'h0000_0006 ? array_update_82366 : array_update_82355[6];
  assign array_update_82368[7] = add_81474 == 32'h0000_0007 ? array_update_82366 : array_update_82355[7];
  assign array_update_82368[8] = add_81474 == 32'h0000_0008 ? array_update_82366 : array_update_82355[8];
  assign array_update_82368[9] = add_81474 == 32'h0000_0009 ? array_update_82366 : array_update_82355[9];
  assign array_index_82370 = array_update_72021[add_82367 > 32'h0000_0009 ? 4'h9 : add_82367[3:0]];
  assign array_index_82371 = array_update_82368[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_82375 = smul32b_32b_x_32b(array_index_81481[add_82367 > 32'h0000_0009 ? 4'h9 : add_82367[3:0]], array_index_82370[add_82287 > 32'h0000_0009 ? 4'h9 : add_82287[3:0]]);
  assign add_82377 = array_index_82371[add_82287 > 32'h0000_0009 ? 4'h9 : add_82287[3:0]] + smul_82375;
  assign array_update_82379[0] = add_82287 == 32'h0000_0000 ? add_82377 : array_index_82371[0];
  assign array_update_82379[1] = add_82287 == 32'h0000_0001 ? add_82377 : array_index_82371[1];
  assign array_update_82379[2] = add_82287 == 32'h0000_0002 ? add_82377 : array_index_82371[2];
  assign array_update_82379[3] = add_82287 == 32'h0000_0003 ? add_82377 : array_index_82371[3];
  assign array_update_82379[4] = add_82287 == 32'h0000_0004 ? add_82377 : array_index_82371[4];
  assign array_update_82379[5] = add_82287 == 32'h0000_0005 ? add_82377 : array_index_82371[5];
  assign array_update_82379[6] = add_82287 == 32'h0000_0006 ? add_82377 : array_index_82371[6];
  assign array_update_82379[7] = add_82287 == 32'h0000_0007 ? add_82377 : array_index_82371[7];
  assign array_update_82379[8] = add_82287 == 32'h0000_0008 ? add_82377 : array_index_82371[8];
  assign array_update_82379[9] = add_82287 == 32'h0000_0009 ? add_82377 : array_index_82371[9];
  assign add_82380 = add_82367 + 32'h0000_0001;
  assign array_update_82381[0] = add_81474 == 32'h0000_0000 ? array_update_82379 : array_update_82368[0];
  assign array_update_82381[1] = add_81474 == 32'h0000_0001 ? array_update_82379 : array_update_82368[1];
  assign array_update_82381[2] = add_81474 == 32'h0000_0002 ? array_update_82379 : array_update_82368[2];
  assign array_update_82381[3] = add_81474 == 32'h0000_0003 ? array_update_82379 : array_update_82368[3];
  assign array_update_82381[4] = add_81474 == 32'h0000_0004 ? array_update_82379 : array_update_82368[4];
  assign array_update_82381[5] = add_81474 == 32'h0000_0005 ? array_update_82379 : array_update_82368[5];
  assign array_update_82381[6] = add_81474 == 32'h0000_0006 ? array_update_82379 : array_update_82368[6];
  assign array_update_82381[7] = add_81474 == 32'h0000_0007 ? array_update_82379 : array_update_82368[7];
  assign array_update_82381[8] = add_81474 == 32'h0000_0008 ? array_update_82379 : array_update_82368[8];
  assign array_update_82381[9] = add_81474 == 32'h0000_0009 ? array_update_82379 : array_update_82368[9];
  assign array_index_82383 = array_update_72021[add_82380 > 32'h0000_0009 ? 4'h9 : add_82380[3:0]];
  assign array_index_82384 = array_update_82381[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_82388 = smul32b_32b_x_32b(array_index_81481[add_82380 > 32'h0000_0009 ? 4'h9 : add_82380[3:0]], array_index_82383[add_82287 > 32'h0000_0009 ? 4'h9 : add_82287[3:0]]);
  assign add_82390 = array_index_82384[add_82287 > 32'h0000_0009 ? 4'h9 : add_82287[3:0]] + smul_82388;
  assign array_update_82392[0] = add_82287 == 32'h0000_0000 ? add_82390 : array_index_82384[0];
  assign array_update_82392[1] = add_82287 == 32'h0000_0001 ? add_82390 : array_index_82384[1];
  assign array_update_82392[2] = add_82287 == 32'h0000_0002 ? add_82390 : array_index_82384[2];
  assign array_update_82392[3] = add_82287 == 32'h0000_0003 ? add_82390 : array_index_82384[3];
  assign array_update_82392[4] = add_82287 == 32'h0000_0004 ? add_82390 : array_index_82384[4];
  assign array_update_82392[5] = add_82287 == 32'h0000_0005 ? add_82390 : array_index_82384[5];
  assign array_update_82392[6] = add_82287 == 32'h0000_0006 ? add_82390 : array_index_82384[6];
  assign array_update_82392[7] = add_82287 == 32'h0000_0007 ? add_82390 : array_index_82384[7];
  assign array_update_82392[8] = add_82287 == 32'h0000_0008 ? add_82390 : array_index_82384[8];
  assign array_update_82392[9] = add_82287 == 32'h0000_0009 ? add_82390 : array_index_82384[9];
  assign add_82393 = add_82380 + 32'h0000_0001;
  assign array_update_82394[0] = add_81474 == 32'h0000_0000 ? array_update_82392 : array_update_82381[0];
  assign array_update_82394[1] = add_81474 == 32'h0000_0001 ? array_update_82392 : array_update_82381[1];
  assign array_update_82394[2] = add_81474 == 32'h0000_0002 ? array_update_82392 : array_update_82381[2];
  assign array_update_82394[3] = add_81474 == 32'h0000_0003 ? array_update_82392 : array_update_82381[3];
  assign array_update_82394[4] = add_81474 == 32'h0000_0004 ? array_update_82392 : array_update_82381[4];
  assign array_update_82394[5] = add_81474 == 32'h0000_0005 ? array_update_82392 : array_update_82381[5];
  assign array_update_82394[6] = add_81474 == 32'h0000_0006 ? array_update_82392 : array_update_82381[6];
  assign array_update_82394[7] = add_81474 == 32'h0000_0007 ? array_update_82392 : array_update_82381[7];
  assign array_update_82394[8] = add_81474 == 32'h0000_0008 ? array_update_82392 : array_update_82381[8];
  assign array_update_82394[9] = add_81474 == 32'h0000_0009 ? array_update_82392 : array_update_82381[9];
  assign array_index_82396 = array_update_72021[add_82393 > 32'h0000_0009 ? 4'h9 : add_82393[3:0]];
  assign array_index_82397 = array_update_82394[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_82401 = smul32b_32b_x_32b(array_index_81481[add_82393 > 32'h0000_0009 ? 4'h9 : add_82393[3:0]], array_index_82396[add_82287 > 32'h0000_0009 ? 4'h9 : add_82287[3:0]]);
  assign add_82403 = array_index_82397[add_82287 > 32'h0000_0009 ? 4'h9 : add_82287[3:0]] + smul_82401;
  assign array_update_82405[0] = add_82287 == 32'h0000_0000 ? add_82403 : array_index_82397[0];
  assign array_update_82405[1] = add_82287 == 32'h0000_0001 ? add_82403 : array_index_82397[1];
  assign array_update_82405[2] = add_82287 == 32'h0000_0002 ? add_82403 : array_index_82397[2];
  assign array_update_82405[3] = add_82287 == 32'h0000_0003 ? add_82403 : array_index_82397[3];
  assign array_update_82405[4] = add_82287 == 32'h0000_0004 ? add_82403 : array_index_82397[4];
  assign array_update_82405[5] = add_82287 == 32'h0000_0005 ? add_82403 : array_index_82397[5];
  assign array_update_82405[6] = add_82287 == 32'h0000_0006 ? add_82403 : array_index_82397[6];
  assign array_update_82405[7] = add_82287 == 32'h0000_0007 ? add_82403 : array_index_82397[7];
  assign array_update_82405[8] = add_82287 == 32'h0000_0008 ? add_82403 : array_index_82397[8];
  assign array_update_82405[9] = add_82287 == 32'h0000_0009 ? add_82403 : array_index_82397[9];
  assign add_82406 = add_82393 + 32'h0000_0001;
  assign array_update_82407[0] = add_81474 == 32'h0000_0000 ? array_update_82405 : array_update_82394[0];
  assign array_update_82407[1] = add_81474 == 32'h0000_0001 ? array_update_82405 : array_update_82394[1];
  assign array_update_82407[2] = add_81474 == 32'h0000_0002 ? array_update_82405 : array_update_82394[2];
  assign array_update_82407[3] = add_81474 == 32'h0000_0003 ? array_update_82405 : array_update_82394[3];
  assign array_update_82407[4] = add_81474 == 32'h0000_0004 ? array_update_82405 : array_update_82394[4];
  assign array_update_82407[5] = add_81474 == 32'h0000_0005 ? array_update_82405 : array_update_82394[5];
  assign array_update_82407[6] = add_81474 == 32'h0000_0006 ? array_update_82405 : array_update_82394[6];
  assign array_update_82407[7] = add_81474 == 32'h0000_0007 ? array_update_82405 : array_update_82394[7];
  assign array_update_82407[8] = add_81474 == 32'h0000_0008 ? array_update_82405 : array_update_82394[8];
  assign array_update_82407[9] = add_81474 == 32'h0000_0009 ? array_update_82405 : array_update_82394[9];
  assign array_index_82409 = array_update_72021[add_82406 > 32'h0000_0009 ? 4'h9 : add_82406[3:0]];
  assign array_index_82410 = array_update_82407[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_82414 = smul32b_32b_x_32b(array_index_81481[add_82406 > 32'h0000_0009 ? 4'h9 : add_82406[3:0]], array_index_82409[add_82287 > 32'h0000_0009 ? 4'h9 : add_82287[3:0]]);
  assign add_82416 = array_index_82410[add_82287 > 32'h0000_0009 ? 4'h9 : add_82287[3:0]] + smul_82414;
  assign array_update_82417[0] = add_82287 == 32'h0000_0000 ? add_82416 : array_index_82410[0];
  assign array_update_82417[1] = add_82287 == 32'h0000_0001 ? add_82416 : array_index_82410[1];
  assign array_update_82417[2] = add_82287 == 32'h0000_0002 ? add_82416 : array_index_82410[2];
  assign array_update_82417[3] = add_82287 == 32'h0000_0003 ? add_82416 : array_index_82410[3];
  assign array_update_82417[4] = add_82287 == 32'h0000_0004 ? add_82416 : array_index_82410[4];
  assign array_update_82417[5] = add_82287 == 32'h0000_0005 ? add_82416 : array_index_82410[5];
  assign array_update_82417[6] = add_82287 == 32'h0000_0006 ? add_82416 : array_index_82410[6];
  assign array_update_82417[7] = add_82287 == 32'h0000_0007 ? add_82416 : array_index_82410[7];
  assign array_update_82417[8] = add_82287 == 32'h0000_0008 ? add_82416 : array_index_82410[8];
  assign array_update_82417[9] = add_82287 == 32'h0000_0009 ? add_82416 : array_index_82410[9];
  assign array_update_82418[0] = add_81474 == 32'h0000_0000 ? array_update_82417 : array_update_82407[0];
  assign array_update_82418[1] = add_81474 == 32'h0000_0001 ? array_update_82417 : array_update_82407[1];
  assign array_update_82418[2] = add_81474 == 32'h0000_0002 ? array_update_82417 : array_update_82407[2];
  assign array_update_82418[3] = add_81474 == 32'h0000_0003 ? array_update_82417 : array_update_82407[3];
  assign array_update_82418[4] = add_81474 == 32'h0000_0004 ? array_update_82417 : array_update_82407[4];
  assign array_update_82418[5] = add_81474 == 32'h0000_0005 ? array_update_82417 : array_update_82407[5];
  assign array_update_82418[6] = add_81474 == 32'h0000_0006 ? array_update_82417 : array_update_82407[6];
  assign array_update_82418[7] = add_81474 == 32'h0000_0007 ? array_update_82417 : array_update_82407[7];
  assign array_update_82418[8] = add_81474 == 32'h0000_0008 ? array_update_82417 : array_update_82407[8];
  assign array_update_82418[9] = add_81474 == 32'h0000_0009 ? array_update_82417 : array_update_82407[9];
  assign array_index_82420 = array_update_82418[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign add_82422 = add_82287 + 32'h0000_0001;
  assign array_update_82423[0] = add_82422 == 32'h0000_0000 ? 32'h0000_0000 : array_index_82420[0];
  assign array_update_82423[1] = add_82422 == 32'h0000_0001 ? 32'h0000_0000 : array_index_82420[1];
  assign array_update_82423[2] = add_82422 == 32'h0000_0002 ? 32'h0000_0000 : array_index_82420[2];
  assign array_update_82423[3] = add_82422 == 32'h0000_0003 ? 32'h0000_0000 : array_index_82420[3];
  assign array_update_82423[4] = add_82422 == 32'h0000_0004 ? 32'h0000_0000 : array_index_82420[4];
  assign array_update_82423[5] = add_82422 == 32'h0000_0005 ? 32'h0000_0000 : array_index_82420[5];
  assign array_update_82423[6] = add_82422 == 32'h0000_0006 ? 32'h0000_0000 : array_index_82420[6];
  assign array_update_82423[7] = add_82422 == 32'h0000_0007 ? 32'h0000_0000 : array_index_82420[7];
  assign array_update_82423[8] = add_82422 == 32'h0000_0008 ? 32'h0000_0000 : array_index_82420[8];
  assign array_update_82423[9] = add_82422 == 32'h0000_0009 ? 32'h0000_0000 : array_index_82420[9];
  assign literal_82424 = 32'h0000_0000;
  assign array_update_82425[0] = add_81474 == 32'h0000_0000 ? array_update_82423 : array_update_82418[0];
  assign array_update_82425[1] = add_81474 == 32'h0000_0001 ? array_update_82423 : array_update_82418[1];
  assign array_update_82425[2] = add_81474 == 32'h0000_0002 ? array_update_82423 : array_update_82418[2];
  assign array_update_82425[3] = add_81474 == 32'h0000_0003 ? array_update_82423 : array_update_82418[3];
  assign array_update_82425[4] = add_81474 == 32'h0000_0004 ? array_update_82423 : array_update_82418[4];
  assign array_update_82425[5] = add_81474 == 32'h0000_0005 ? array_update_82423 : array_update_82418[5];
  assign array_update_82425[6] = add_81474 == 32'h0000_0006 ? array_update_82423 : array_update_82418[6];
  assign array_update_82425[7] = add_81474 == 32'h0000_0007 ? array_update_82423 : array_update_82418[7];
  assign array_update_82425[8] = add_81474 == 32'h0000_0008 ? array_update_82423 : array_update_82418[8];
  assign array_update_82425[9] = add_81474 == 32'h0000_0009 ? array_update_82423 : array_update_82418[9];
  assign array_index_82427 = array_update_72021[literal_82424 > 32'h0000_0009 ? 4'h9 : literal_82424[3:0]];
  assign array_index_82428 = array_update_82425[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_82432 = smul32b_32b_x_32b(array_index_81481[literal_82424 > 32'h0000_0009 ? 4'h9 : literal_82424[3:0]], array_index_82427[add_82422 > 32'h0000_0009 ? 4'h9 : add_82422[3:0]]);
  assign add_82434 = array_index_82428[add_82422 > 32'h0000_0009 ? 4'h9 : add_82422[3:0]] + smul_82432;
  assign array_update_82436[0] = add_82422 == 32'h0000_0000 ? add_82434 : array_index_82428[0];
  assign array_update_82436[1] = add_82422 == 32'h0000_0001 ? add_82434 : array_index_82428[1];
  assign array_update_82436[2] = add_82422 == 32'h0000_0002 ? add_82434 : array_index_82428[2];
  assign array_update_82436[3] = add_82422 == 32'h0000_0003 ? add_82434 : array_index_82428[3];
  assign array_update_82436[4] = add_82422 == 32'h0000_0004 ? add_82434 : array_index_82428[4];
  assign array_update_82436[5] = add_82422 == 32'h0000_0005 ? add_82434 : array_index_82428[5];
  assign array_update_82436[6] = add_82422 == 32'h0000_0006 ? add_82434 : array_index_82428[6];
  assign array_update_82436[7] = add_82422 == 32'h0000_0007 ? add_82434 : array_index_82428[7];
  assign array_update_82436[8] = add_82422 == 32'h0000_0008 ? add_82434 : array_index_82428[8];
  assign array_update_82436[9] = add_82422 == 32'h0000_0009 ? add_82434 : array_index_82428[9];
  assign add_82437 = literal_82424 + 32'h0000_0001;
  assign array_update_82438[0] = add_81474 == 32'h0000_0000 ? array_update_82436 : array_update_82425[0];
  assign array_update_82438[1] = add_81474 == 32'h0000_0001 ? array_update_82436 : array_update_82425[1];
  assign array_update_82438[2] = add_81474 == 32'h0000_0002 ? array_update_82436 : array_update_82425[2];
  assign array_update_82438[3] = add_81474 == 32'h0000_0003 ? array_update_82436 : array_update_82425[3];
  assign array_update_82438[4] = add_81474 == 32'h0000_0004 ? array_update_82436 : array_update_82425[4];
  assign array_update_82438[5] = add_81474 == 32'h0000_0005 ? array_update_82436 : array_update_82425[5];
  assign array_update_82438[6] = add_81474 == 32'h0000_0006 ? array_update_82436 : array_update_82425[6];
  assign array_update_82438[7] = add_81474 == 32'h0000_0007 ? array_update_82436 : array_update_82425[7];
  assign array_update_82438[8] = add_81474 == 32'h0000_0008 ? array_update_82436 : array_update_82425[8];
  assign array_update_82438[9] = add_81474 == 32'h0000_0009 ? array_update_82436 : array_update_82425[9];
  assign array_index_82440 = array_update_72021[add_82437 > 32'h0000_0009 ? 4'h9 : add_82437[3:0]];
  assign array_index_82441 = array_update_82438[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_82445 = smul32b_32b_x_32b(array_index_81481[add_82437 > 32'h0000_0009 ? 4'h9 : add_82437[3:0]], array_index_82440[add_82422 > 32'h0000_0009 ? 4'h9 : add_82422[3:0]]);
  assign add_82447 = array_index_82441[add_82422 > 32'h0000_0009 ? 4'h9 : add_82422[3:0]] + smul_82445;
  assign array_update_82449[0] = add_82422 == 32'h0000_0000 ? add_82447 : array_index_82441[0];
  assign array_update_82449[1] = add_82422 == 32'h0000_0001 ? add_82447 : array_index_82441[1];
  assign array_update_82449[2] = add_82422 == 32'h0000_0002 ? add_82447 : array_index_82441[2];
  assign array_update_82449[3] = add_82422 == 32'h0000_0003 ? add_82447 : array_index_82441[3];
  assign array_update_82449[4] = add_82422 == 32'h0000_0004 ? add_82447 : array_index_82441[4];
  assign array_update_82449[5] = add_82422 == 32'h0000_0005 ? add_82447 : array_index_82441[5];
  assign array_update_82449[6] = add_82422 == 32'h0000_0006 ? add_82447 : array_index_82441[6];
  assign array_update_82449[7] = add_82422 == 32'h0000_0007 ? add_82447 : array_index_82441[7];
  assign array_update_82449[8] = add_82422 == 32'h0000_0008 ? add_82447 : array_index_82441[8];
  assign array_update_82449[9] = add_82422 == 32'h0000_0009 ? add_82447 : array_index_82441[9];
  assign add_82450 = add_82437 + 32'h0000_0001;
  assign array_update_82451[0] = add_81474 == 32'h0000_0000 ? array_update_82449 : array_update_82438[0];
  assign array_update_82451[1] = add_81474 == 32'h0000_0001 ? array_update_82449 : array_update_82438[1];
  assign array_update_82451[2] = add_81474 == 32'h0000_0002 ? array_update_82449 : array_update_82438[2];
  assign array_update_82451[3] = add_81474 == 32'h0000_0003 ? array_update_82449 : array_update_82438[3];
  assign array_update_82451[4] = add_81474 == 32'h0000_0004 ? array_update_82449 : array_update_82438[4];
  assign array_update_82451[5] = add_81474 == 32'h0000_0005 ? array_update_82449 : array_update_82438[5];
  assign array_update_82451[6] = add_81474 == 32'h0000_0006 ? array_update_82449 : array_update_82438[6];
  assign array_update_82451[7] = add_81474 == 32'h0000_0007 ? array_update_82449 : array_update_82438[7];
  assign array_update_82451[8] = add_81474 == 32'h0000_0008 ? array_update_82449 : array_update_82438[8];
  assign array_update_82451[9] = add_81474 == 32'h0000_0009 ? array_update_82449 : array_update_82438[9];
  assign array_index_82453 = array_update_72021[add_82450 > 32'h0000_0009 ? 4'h9 : add_82450[3:0]];
  assign array_index_82454 = array_update_82451[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_82458 = smul32b_32b_x_32b(array_index_81481[add_82450 > 32'h0000_0009 ? 4'h9 : add_82450[3:0]], array_index_82453[add_82422 > 32'h0000_0009 ? 4'h9 : add_82422[3:0]]);
  assign add_82460 = array_index_82454[add_82422 > 32'h0000_0009 ? 4'h9 : add_82422[3:0]] + smul_82458;
  assign array_update_82462[0] = add_82422 == 32'h0000_0000 ? add_82460 : array_index_82454[0];
  assign array_update_82462[1] = add_82422 == 32'h0000_0001 ? add_82460 : array_index_82454[1];
  assign array_update_82462[2] = add_82422 == 32'h0000_0002 ? add_82460 : array_index_82454[2];
  assign array_update_82462[3] = add_82422 == 32'h0000_0003 ? add_82460 : array_index_82454[3];
  assign array_update_82462[4] = add_82422 == 32'h0000_0004 ? add_82460 : array_index_82454[4];
  assign array_update_82462[5] = add_82422 == 32'h0000_0005 ? add_82460 : array_index_82454[5];
  assign array_update_82462[6] = add_82422 == 32'h0000_0006 ? add_82460 : array_index_82454[6];
  assign array_update_82462[7] = add_82422 == 32'h0000_0007 ? add_82460 : array_index_82454[7];
  assign array_update_82462[8] = add_82422 == 32'h0000_0008 ? add_82460 : array_index_82454[8];
  assign array_update_82462[9] = add_82422 == 32'h0000_0009 ? add_82460 : array_index_82454[9];
  assign add_82463 = add_82450 + 32'h0000_0001;
  assign array_update_82464[0] = add_81474 == 32'h0000_0000 ? array_update_82462 : array_update_82451[0];
  assign array_update_82464[1] = add_81474 == 32'h0000_0001 ? array_update_82462 : array_update_82451[1];
  assign array_update_82464[2] = add_81474 == 32'h0000_0002 ? array_update_82462 : array_update_82451[2];
  assign array_update_82464[3] = add_81474 == 32'h0000_0003 ? array_update_82462 : array_update_82451[3];
  assign array_update_82464[4] = add_81474 == 32'h0000_0004 ? array_update_82462 : array_update_82451[4];
  assign array_update_82464[5] = add_81474 == 32'h0000_0005 ? array_update_82462 : array_update_82451[5];
  assign array_update_82464[6] = add_81474 == 32'h0000_0006 ? array_update_82462 : array_update_82451[6];
  assign array_update_82464[7] = add_81474 == 32'h0000_0007 ? array_update_82462 : array_update_82451[7];
  assign array_update_82464[8] = add_81474 == 32'h0000_0008 ? array_update_82462 : array_update_82451[8];
  assign array_update_82464[9] = add_81474 == 32'h0000_0009 ? array_update_82462 : array_update_82451[9];
  assign array_index_82466 = array_update_72021[add_82463 > 32'h0000_0009 ? 4'h9 : add_82463[3:0]];
  assign array_index_82467 = array_update_82464[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_82471 = smul32b_32b_x_32b(array_index_81481[add_82463 > 32'h0000_0009 ? 4'h9 : add_82463[3:0]], array_index_82466[add_82422 > 32'h0000_0009 ? 4'h9 : add_82422[3:0]]);
  assign add_82473 = array_index_82467[add_82422 > 32'h0000_0009 ? 4'h9 : add_82422[3:0]] + smul_82471;
  assign array_update_82475[0] = add_82422 == 32'h0000_0000 ? add_82473 : array_index_82467[0];
  assign array_update_82475[1] = add_82422 == 32'h0000_0001 ? add_82473 : array_index_82467[1];
  assign array_update_82475[2] = add_82422 == 32'h0000_0002 ? add_82473 : array_index_82467[2];
  assign array_update_82475[3] = add_82422 == 32'h0000_0003 ? add_82473 : array_index_82467[3];
  assign array_update_82475[4] = add_82422 == 32'h0000_0004 ? add_82473 : array_index_82467[4];
  assign array_update_82475[5] = add_82422 == 32'h0000_0005 ? add_82473 : array_index_82467[5];
  assign array_update_82475[6] = add_82422 == 32'h0000_0006 ? add_82473 : array_index_82467[6];
  assign array_update_82475[7] = add_82422 == 32'h0000_0007 ? add_82473 : array_index_82467[7];
  assign array_update_82475[8] = add_82422 == 32'h0000_0008 ? add_82473 : array_index_82467[8];
  assign array_update_82475[9] = add_82422 == 32'h0000_0009 ? add_82473 : array_index_82467[9];
  assign add_82476 = add_82463 + 32'h0000_0001;
  assign array_update_82477[0] = add_81474 == 32'h0000_0000 ? array_update_82475 : array_update_82464[0];
  assign array_update_82477[1] = add_81474 == 32'h0000_0001 ? array_update_82475 : array_update_82464[1];
  assign array_update_82477[2] = add_81474 == 32'h0000_0002 ? array_update_82475 : array_update_82464[2];
  assign array_update_82477[3] = add_81474 == 32'h0000_0003 ? array_update_82475 : array_update_82464[3];
  assign array_update_82477[4] = add_81474 == 32'h0000_0004 ? array_update_82475 : array_update_82464[4];
  assign array_update_82477[5] = add_81474 == 32'h0000_0005 ? array_update_82475 : array_update_82464[5];
  assign array_update_82477[6] = add_81474 == 32'h0000_0006 ? array_update_82475 : array_update_82464[6];
  assign array_update_82477[7] = add_81474 == 32'h0000_0007 ? array_update_82475 : array_update_82464[7];
  assign array_update_82477[8] = add_81474 == 32'h0000_0008 ? array_update_82475 : array_update_82464[8];
  assign array_update_82477[9] = add_81474 == 32'h0000_0009 ? array_update_82475 : array_update_82464[9];
  assign array_index_82479 = array_update_72021[add_82476 > 32'h0000_0009 ? 4'h9 : add_82476[3:0]];
  assign array_index_82480 = array_update_82477[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_82484 = smul32b_32b_x_32b(array_index_81481[add_82476 > 32'h0000_0009 ? 4'h9 : add_82476[3:0]], array_index_82479[add_82422 > 32'h0000_0009 ? 4'h9 : add_82422[3:0]]);
  assign add_82486 = array_index_82480[add_82422 > 32'h0000_0009 ? 4'h9 : add_82422[3:0]] + smul_82484;
  assign array_update_82488[0] = add_82422 == 32'h0000_0000 ? add_82486 : array_index_82480[0];
  assign array_update_82488[1] = add_82422 == 32'h0000_0001 ? add_82486 : array_index_82480[1];
  assign array_update_82488[2] = add_82422 == 32'h0000_0002 ? add_82486 : array_index_82480[2];
  assign array_update_82488[3] = add_82422 == 32'h0000_0003 ? add_82486 : array_index_82480[3];
  assign array_update_82488[4] = add_82422 == 32'h0000_0004 ? add_82486 : array_index_82480[4];
  assign array_update_82488[5] = add_82422 == 32'h0000_0005 ? add_82486 : array_index_82480[5];
  assign array_update_82488[6] = add_82422 == 32'h0000_0006 ? add_82486 : array_index_82480[6];
  assign array_update_82488[7] = add_82422 == 32'h0000_0007 ? add_82486 : array_index_82480[7];
  assign array_update_82488[8] = add_82422 == 32'h0000_0008 ? add_82486 : array_index_82480[8];
  assign array_update_82488[9] = add_82422 == 32'h0000_0009 ? add_82486 : array_index_82480[9];
  assign add_82489 = add_82476 + 32'h0000_0001;
  assign array_update_82490[0] = add_81474 == 32'h0000_0000 ? array_update_82488 : array_update_82477[0];
  assign array_update_82490[1] = add_81474 == 32'h0000_0001 ? array_update_82488 : array_update_82477[1];
  assign array_update_82490[2] = add_81474 == 32'h0000_0002 ? array_update_82488 : array_update_82477[2];
  assign array_update_82490[3] = add_81474 == 32'h0000_0003 ? array_update_82488 : array_update_82477[3];
  assign array_update_82490[4] = add_81474 == 32'h0000_0004 ? array_update_82488 : array_update_82477[4];
  assign array_update_82490[5] = add_81474 == 32'h0000_0005 ? array_update_82488 : array_update_82477[5];
  assign array_update_82490[6] = add_81474 == 32'h0000_0006 ? array_update_82488 : array_update_82477[6];
  assign array_update_82490[7] = add_81474 == 32'h0000_0007 ? array_update_82488 : array_update_82477[7];
  assign array_update_82490[8] = add_81474 == 32'h0000_0008 ? array_update_82488 : array_update_82477[8];
  assign array_update_82490[9] = add_81474 == 32'h0000_0009 ? array_update_82488 : array_update_82477[9];
  assign array_index_82492 = array_update_72021[add_82489 > 32'h0000_0009 ? 4'h9 : add_82489[3:0]];
  assign array_index_82493 = array_update_82490[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_82497 = smul32b_32b_x_32b(array_index_81481[add_82489 > 32'h0000_0009 ? 4'h9 : add_82489[3:0]], array_index_82492[add_82422 > 32'h0000_0009 ? 4'h9 : add_82422[3:0]]);
  assign add_82499 = array_index_82493[add_82422 > 32'h0000_0009 ? 4'h9 : add_82422[3:0]] + smul_82497;
  assign array_update_82501[0] = add_82422 == 32'h0000_0000 ? add_82499 : array_index_82493[0];
  assign array_update_82501[1] = add_82422 == 32'h0000_0001 ? add_82499 : array_index_82493[1];
  assign array_update_82501[2] = add_82422 == 32'h0000_0002 ? add_82499 : array_index_82493[2];
  assign array_update_82501[3] = add_82422 == 32'h0000_0003 ? add_82499 : array_index_82493[3];
  assign array_update_82501[4] = add_82422 == 32'h0000_0004 ? add_82499 : array_index_82493[4];
  assign array_update_82501[5] = add_82422 == 32'h0000_0005 ? add_82499 : array_index_82493[5];
  assign array_update_82501[6] = add_82422 == 32'h0000_0006 ? add_82499 : array_index_82493[6];
  assign array_update_82501[7] = add_82422 == 32'h0000_0007 ? add_82499 : array_index_82493[7];
  assign array_update_82501[8] = add_82422 == 32'h0000_0008 ? add_82499 : array_index_82493[8];
  assign array_update_82501[9] = add_82422 == 32'h0000_0009 ? add_82499 : array_index_82493[9];
  assign add_82502 = add_82489 + 32'h0000_0001;
  assign array_update_82503[0] = add_81474 == 32'h0000_0000 ? array_update_82501 : array_update_82490[0];
  assign array_update_82503[1] = add_81474 == 32'h0000_0001 ? array_update_82501 : array_update_82490[1];
  assign array_update_82503[2] = add_81474 == 32'h0000_0002 ? array_update_82501 : array_update_82490[2];
  assign array_update_82503[3] = add_81474 == 32'h0000_0003 ? array_update_82501 : array_update_82490[3];
  assign array_update_82503[4] = add_81474 == 32'h0000_0004 ? array_update_82501 : array_update_82490[4];
  assign array_update_82503[5] = add_81474 == 32'h0000_0005 ? array_update_82501 : array_update_82490[5];
  assign array_update_82503[6] = add_81474 == 32'h0000_0006 ? array_update_82501 : array_update_82490[6];
  assign array_update_82503[7] = add_81474 == 32'h0000_0007 ? array_update_82501 : array_update_82490[7];
  assign array_update_82503[8] = add_81474 == 32'h0000_0008 ? array_update_82501 : array_update_82490[8];
  assign array_update_82503[9] = add_81474 == 32'h0000_0009 ? array_update_82501 : array_update_82490[9];
  assign array_index_82505 = array_update_72021[add_82502 > 32'h0000_0009 ? 4'h9 : add_82502[3:0]];
  assign array_index_82506 = array_update_82503[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_82510 = smul32b_32b_x_32b(array_index_81481[add_82502 > 32'h0000_0009 ? 4'h9 : add_82502[3:0]], array_index_82505[add_82422 > 32'h0000_0009 ? 4'h9 : add_82422[3:0]]);
  assign add_82512 = array_index_82506[add_82422 > 32'h0000_0009 ? 4'h9 : add_82422[3:0]] + smul_82510;
  assign array_update_82514[0] = add_82422 == 32'h0000_0000 ? add_82512 : array_index_82506[0];
  assign array_update_82514[1] = add_82422 == 32'h0000_0001 ? add_82512 : array_index_82506[1];
  assign array_update_82514[2] = add_82422 == 32'h0000_0002 ? add_82512 : array_index_82506[2];
  assign array_update_82514[3] = add_82422 == 32'h0000_0003 ? add_82512 : array_index_82506[3];
  assign array_update_82514[4] = add_82422 == 32'h0000_0004 ? add_82512 : array_index_82506[4];
  assign array_update_82514[5] = add_82422 == 32'h0000_0005 ? add_82512 : array_index_82506[5];
  assign array_update_82514[6] = add_82422 == 32'h0000_0006 ? add_82512 : array_index_82506[6];
  assign array_update_82514[7] = add_82422 == 32'h0000_0007 ? add_82512 : array_index_82506[7];
  assign array_update_82514[8] = add_82422 == 32'h0000_0008 ? add_82512 : array_index_82506[8];
  assign array_update_82514[9] = add_82422 == 32'h0000_0009 ? add_82512 : array_index_82506[9];
  assign add_82515 = add_82502 + 32'h0000_0001;
  assign array_update_82516[0] = add_81474 == 32'h0000_0000 ? array_update_82514 : array_update_82503[0];
  assign array_update_82516[1] = add_81474 == 32'h0000_0001 ? array_update_82514 : array_update_82503[1];
  assign array_update_82516[2] = add_81474 == 32'h0000_0002 ? array_update_82514 : array_update_82503[2];
  assign array_update_82516[3] = add_81474 == 32'h0000_0003 ? array_update_82514 : array_update_82503[3];
  assign array_update_82516[4] = add_81474 == 32'h0000_0004 ? array_update_82514 : array_update_82503[4];
  assign array_update_82516[5] = add_81474 == 32'h0000_0005 ? array_update_82514 : array_update_82503[5];
  assign array_update_82516[6] = add_81474 == 32'h0000_0006 ? array_update_82514 : array_update_82503[6];
  assign array_update_82516[7] = add_81474 == 32'h0000_0007 ? array_update_82514 : array_update_82503[7];
  assign array_update_82516[8] = add_81474 == 32'h0000_0008 ? array_update_82514 : array_update_82503[8];
  assign array_update_82516[9] = add_81474 == 32'h0000_0009 ? array_update_82514 : array_update_82503[9];
  assign array_index_82518 = array_update_72021[add_82515 > 32'h0000_0009 ? 4'h9 : add_82515[3:0]];
  assign array_index_82519 = array_update_82516[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_82523 = smul32b_32b_x_32b(array_index_81481[add_82515 > 32'h0000_0009 ? 4'h9 : add_82515[3:0]], array_index_82518[add_82422 > 32'h0000_0009 ? 4'h9 : add_82422[3:0]]);
  assign add_82525 = array_index_82519[add_82422 > 32'h0000_0009 ? 4'h9 : add_82422[3:0]] + smul_82523;
  assign array_update_82527[0] = add_82422 == 32'h0000_0000 ? add_82525 : array_index_82519[0];
  assign array_update_82527[1] = add_82422 == 32'h0000_0001 ? add_82525 : array_index_82519[1];
  assign array_update_82527[2] = add_82422 == 32'h0000_0002 ? add_82525 : array_index_82519[2];
  assign array_update_82527[3] = add_82422 == 32'h0000_0003 ? add_82525 : array_index_82519[3];
  assign array_update_82527[4] = add_82422 == 32'h0000_0004 ? add_82525 : array_index_82519[4];
  assign array_update_82527[5] = add_82422 == 32'h0000_0005 ? add_82525 : array_index_82519[5];
  assign array_update_82527[6] = add_82422 == 32'h0000_0006 ? add_82525 : array_index_82519[6];
  assign array_update_82527[7] = add_82422 == 32'h0000_0007 ? add_82525 : array_index_82519[7];
  assign array_update_82527[8] = add_82422 == 32'h0000_0008 ? add_82525 : array_index_82519[8];
  assign array_update_82527[9] = add_82422 == 32'h0000_0009 ? add_82525 : array_index_82519[9];
  assign add_82528 = add_82515 + 32'h0000_0001;
  assign array_update_82529[0] = add_81474 == 32'h0000_0000 ? array_update_82527 : array_update_82516[0];
  assign array_update_82529[1] = add_81474 == 32'h0000_0001 ? array_update_82527 : array_update_82516[1];
  assign array_update_82529[2] = add_81474 == 32'h0000_0002 ? array_update_82527 : array_update_82516[2];
  assign array_update_82529[3] = add_81474 == 32'h0000_0003 ? array_update_82527 : array_update_82516[3];
  assign array_update_82529[4] = add_81474 == 32'h0000_0004 ? array_update_82527 : array_update_82516[4];
  assign array_update_82529[5] = add_81474 == 32'h0000_0005 ? array_update_82527 : array_update_82516[5];
  assign array_update_82529[6] = add_81474 == 32'h0000_0006 ? array_update_82527 : array_update_82516[6];
  assign array_update_82529[7] = add_81474 == 32'h0000_0007 ? array_update_82527 : array_update_82516[7];
  assign array_update_82529[8] = add_81474 == 32'h0000_0008 ? array_update_82527 : array_update_82516[8];
  assign array_update_82529[9] = add_81474 == 32'h0000_0009 ? array_update_82527 : array_update_82516[9];
  assign array_index_82531 = array_update_72021[add_82528 > 32'h0000_0009 ? 4'h9 : add_82528[3:0]];
  assign array_index_82532 = array_update_82529[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_82536 = smul32b_32b_x_32b(array_index_81481[add_82528 > 32'h0000_0009 ? 4'h9 : add_82528[3:0]], array_index_82531[add_82422 > 32'h0000_0009 ? 4'h9 : add_82422[3:0]]);
  assign add_82538 = array_index_82532[add_82422 > 32'h0000_0009 ? 4'h9 : add_82422[3:0]] + smul_82536;
  assign array_update_82540[0] = add_82422 == 32'h0000_0000 ? add_82538 : array_index_82532[0];
  assign array_update_82540[1] = add_82422 == 32'h0000_0001 ? add_82538 : array_index_82532[1];
  assign array_update_82540[2] = add_82422 == 32'h0000_0002 ? add_82538 : array_index_82532[2];
  assign array_update_82540[3] = add_82422 == 32'h0000_0003 ? add_82538 : array_index_82532[3];
  assign array_update_82540[4] = add_82422 == 32'h0000_0004 ? add_82538 : array_index_82532[4];
  assign array_update_82540[5] = add_82422 == 32'h0000_0005 ? add_82538 : array_index_82532[5];
  assign array_update_82540[6] = add_82422 == 32'h0000_0006 ? add_82538 : array_index_82532[6];
  assign array_update_82540[7] = add_82422 == 32'h0000_0007 ? add_82538 : array_index_82532[7];
  assign array_update_82540[8] = add_82422 == 32'h0000_0008 ? add_82538 : array_index_82532[8];
  assign array_update_82540[9] = add_82422 == 32'h0000_0009 ? add_82538 : array_index_82532[9];
  assign add_82541 = add_82528 + 32'h0000_0001;
  assign array_update_82542[0] = add_81474 == 32'h0000_0000 ? array_update_82540 : array_update_82529[0];
  assign array_update_82542[1] = add_81474 == 32'h0000_0001 ? array_update_82540 : array_update_82529[1];
  assign array_update_82542[2] = add_81474 == 32'h0000_0002 ? array_update_82540 : array_update_82529[2];
  assign array_update_82542[3] = add_81474 == 32'h0000_0003 ? array_update_82540 : array_update_82529[3];
  assign array_update_82542[4] = add_81474 == 32'h0000_0004 ? array_update_82540 : array_update_82529[4];
  assign array_update_82542[5] = add_81474 == 32'h0000_0005 ? array_update_82540 : array_update_82529[5];
  assign array_update_82542[6] = add_81474 == 32'h0000_0006 ? array_update_82540 : array_update_82529[6];
  assign array_update_82542[7] = add_81474 == 32'h0000_0007 ? array_update_82540 : array_update_82529[7];
  assign array_update_82542[8] = add_81474 == 32'h0000_0008 ? array_update_82540 : array_update_82529[8];
  assign array_update_82542[9] = add_81474 == 32'h0000_0009 ? array_update_82540 : array_update_82529[9];
  assign array_index_82544 = array_update_72021[add_82541 > 32'h0000_0009 ? 4'h9 : add_82541[3:0]];
  assign array_index_82545 = array_update_82542[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_82549 = smul32b_32b_x_32b(array_index_81481[add_82541 > 32'h0000_0009 ? 4'h9 : add_82541[3:0]], array_index_82544[add_82422 > 32'h0000_0009 ? 4'h9 : add_82422[3:0]]);
  assign add_82551 = array_index_82545[add_82422 > 32'h0000_0009 ? 4'h9 : add_82422[3:0]] + smul_82549;
  assign array_update_82552[0] = add_82422 == 32'h0000_0000 ? add_82551 : array_index_82545[0];
  assign array_update_82552[1] = add_82422 == 32'h0000_0001 ? add_82551 : array_index_82545[1];
  assign array_update_82552[2] = add_82422 == 32'h0000_0002 ? add_82551 : array_index_82545[2];
  assign array_update_82552[3] = add_82422 == 32'h0000_0003 ? add_82551 : array_index_82545[3];
  assign array_update_82552[4] = add_82422 == 32'h0000_0004 ? add_82551 : array_index_82545[4];
  assign array_update_82552[5] = add_82422 == 32'h0000_0005 ? add_82551 : array_index_82545[5];
  assign array_update_82552[6] = add_82422 == 32'h0000_0006 ? add_82551 : array_index_82545[6];
  assign array_update_82552[7] = add_82422 == 32'h0000_0007 ? add_82551 : array_index_82545[7];
  assign array_update_82552[8] = add_82422 == 32'h0000_0008 ? add_82551 : array_index_82545[8];
  assign array_update_82552[9] = add_82422 == 32'h0000_0009 ? add_82551 : array_index_82545[9];
  assign array_update_82553[0] = add_81474 == 32'h0000_0000 ? array_update_82552 : array_update_82542[0];
  assign array_update_82553[1] = add_81474 == 32'h0000_0001 ? array_update_82552 : array_update_82542[1];
  assign array_update_82553[2] = add_81474 == 32'h0000_0002 ? array_update_82552 : array_update_82542[2];
  assign array_update_82553[3] = add_81474 == 32'h0000_0003 ? array_update_82552 : array_update_82542[3];
  assign array_update_82553[4] = add_81474 == 32'h0000_0004 ? array_update_82552 : array_update_82542[4];
  assign array_update_82553[5] = add_81474 == 32'h0000_0005 ? array_update_82552 : array_update_82542[5];
  assign array_update_82553[6] = add_81474 == 32'h0000_0006 ? array_update_82552 : array_update_82542[6];
  assign array_update_82553[7] = add_81474 == 32'h0000_0007 ? array_update_82552 : array_update_82542[7];
  assign array_update_82553[8] = add_81474 == 32'h0000_0008 ? array_update_82552 : array_update_82542[8];
  assign array_update_82553[9] = add_81474 == 32'h0000_0009 ? array_update_82552 : array_update_82542[9];
  assign array_index_82555 = array_update_82553[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign add_82557 = add_82422 + 32'h0000_0001;
  assign array_update_82558[0] = add_82557 == 32'h0000_0000 ? 32'h0000_0000 : array_index_82555[0];
  assign array_update_82558[1] = add_82557 == 32'h0000_0001 ? 32'h0000_0000 : array_index_82555[1];
  assign array_update_82558[2] = add_82557 == 32'h0000_0002 ? 32'h0000_0000 : array_index_82555[2];
  assign array_update_82558[3] = add_82557 == 32'h0000_0003 ? 32'h0000_0000 : array_index_82555[3];
  assign array_update_82558[4] = add_82557 == 32'h0000_0004 ? 32'h0000_0000 : array_index_82555[4];
  assign array_update_82558[5] = add_82557 == 32'h0000_0005 ? 32'h0000_0000 : array_index_82555[5];
  assign array_update_82558[6] = add_82557 == 32'h0000_0006 ? 32'h0000_0000 : array_index_82555[6];
  assign array_update_82558[7] = add_82557 == 32'h0000_0007 ? 32'h0000_0000 : array_index_82555[7];
  assign array_update_82558[8] = add_82557 == 32'h0000_0008 ? 32'h0000_0000 : array_index_82555[8];
  assign array_update_82558[9] = add_82557 == 32'h0000_0009 ? 32'h0000_0000 : array_index_82555[9];
  assign literal_82559 = 32'h0000_0000;
  assign array_update_82560[0] = add_81474 == 32'h0000_0000 ? array_update_82558 : array_update_82553[0];
  assign array_update_82560[1] = add_81474 == 32'h0000_0001 ? array_update_82558 : array_update_82553[1];
  assign array_update_82560[2] = add_81474 == 32'h0000_0002 ? array_update_82558 : array_update_82553[2];
  assign array_update_82560[3] = add_81474 == 32'h0000_0003 ? array_update_82558 : array_update_82553[3];
  assign array_update_82560[4] = add_81474 == 32'h0000_0004 ? array_update_82558 : array_update_82553[4];
  assign array_update_82560[5] = add_81474 == 32'h0000_0005 ? array_update_82558 : array_update_82553[5];
  assign array_update_82560[6] = add_81474 == 32'h0000_0006 ? array_update_82558 : array_update_82553[6];
  assign array_update_82560[7] = add_81474 == 32'h0000_0007 ? array_update_82558 : array_update_82553[7];
  assign array_update_82560[8] = add_81474 == 32'h0000_0008 ? array_update_82558 : array_update_82553[8];
  assign array_update_82560[9] = add_81474 == 32'h0000_0009 ? array_update_82558 : array_update_82553[9];
  assign array_index_82562 = array_update_72021[literal_82559 > 32'h0000_0009 ? 4'h9 : literal_82559[3:0]];
  assign array_index_82563 = array_update_82560[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_82567 = smul32b_32b_x_32b(array_index_81481[literal_82559 > 32'h0000_0009 ? 4'h9 : literal_82559[3:0]], array_index_82562[add_82557 > 32'h0000_0009 ? 4'h9 : add_82557[3:0]]);
  assign add_82569 = array_index_82563[add_82557 > 32'h0000_0009 ? 4'h9 : add_82557[3:0]] + smul_82567;
  assign array_update_82571[0] = add_82557 == 32'h0000_0000 ? add_82569 : array_index_82563[0];
  assign array_update_82571[1] = add_82557 == 32'h0000_0001 ? add_82569 : array_index_82563[1];
  assign array_update_82571[2] = add_82557 == 32'h0000_0002 ? add_82569 : array_index_82563[2];
  assign array_update_82571[3] = add_82557 == 32'h0000_0003 ? add_82569 : array_index_82563[3];
  assign array_update_82571[4] = add_82557 == 32'h0000_0004 ? add_82569 : array_index_82563[4];
  assign array_update_82571[5] = add_82557 == 32'h0000_0005 ? add_82569 : array_index_82563[5];
  assign array_update_82571[6] = add_82557 == 32'h0000_0006 ? add_82569 : array_index_82563[6];
  assign array_update_82571[7] = add_82557 == 32'h0000_0007 ? add_82569 : array_index_82563[7];
  assign array_update_82571[8] = add_82557 == 32'h0000_0008 ? add_82569 : array_index_82563[8];
  assign array_update_82571[9] = add_82557 == 32'h0000_0009 ? add_82569 : array_index_82563[9];
  assign add_82572 = literal_82559 + 32'h0000_0001;
  assign array_update_82573[0] = add_81474 == 32'h0000_0000 ? array_update_82571 : array_update_82560[0];
  assign array_update_82573[1] = add_81474 == 32'h0000_0001 ? array_update_82571 : array_update_82560[1];
  assign array_update_82573[2] = add_81474 == 32'h0000_0002 ? array_update_82571 : array_update_82560[2];
  assign array_update_82573[3] = add_81474 == 32'h0000_0003 ? array_update_82571 : array_update_82560[3];
  assign array_update_82573[4] = add_81474 == 32'h0000_0004 ? array_update_82571 : array_update_82560[4];
  assign array_update_82573[5] = add_81474 == 32'h0000_0005 ? array_update_82571 : array_update_82560[5];
  assign array_update_82573[6] = add_81474 == 32'h0000_0006 ? array_update_82571 : array_update_82560[6];
  assign array_update_82573[7] = add_81474 == 32'h0000_0007 ? array_update_82571 : array_update_82560[7];
  assign array_update_82573[8] = add_81474 == 32'h0000_0008 ? array_update_82571 : array_update_82560[8];
  assign array_update_82573[9] = add_81474 == 32'h0000_0009 ? array_update_82571 : array_update_82560[9];
  assign array_index_82575 = array_update_72021[add_82572 > 32'h0000_0009 ? 4'h9 : add_82572[3:0]];
  assign array_index_82576 = array_update_82573[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_82580 = smul32b_32b_x_32b(array_index_81481[add_82572 > 32'h0000_0009 ? 4'h9 : add_82572[3:0]], array_index_82575[add_82557 > 32'h0000_0009 ? 4'h9 : add_82557[3:0]]);
  assign add_82582 = array_index_82576[add_82557 > 32'h0000_0009 ? 4'h9 : add_82557[3:0]] + smul_82580;
  assign array_update_82584[0] = add_82557 == 32'h0000_0000 ? add_82582 : array_index_82576[0];
  assign array_update_82584[1] = add_82557 == 32'h0000_0001 ? add_82582 : array_index_82576[1];
  assign array_update_82584[2] = add_82557 == 32'h0000_0002 ? add_82582 : array_index_82576[2];
  assign array_update_82584[3] = add_82557 == 32'h0000_0003 ? add_82582 : array_index_82576[3];
  assign array_update_82584[4] = add_82557 == 32'h0000_0004 ? add_82582 : array_index_82576[4];
  assign array_update_82584[5] = add_82557 == 32'h0000_0005 ? add_82582 : array_index_82576[5];
  assign array_update_82584[6] = add_82557 == 32'h0000_0006 ? add_82582 : array_index_82576[6];
  assign array_update_82584[7] = add_82557 == 32'h0000_0007 ? add_82582 : array_index_82576[7];
  assign array_update_82584[8] = add_82557 == 32'h0000_0008 ? add_82582 : array_index_82576[8];
  assign array_update_82584[9] = add_82557 == 32'h0000_0009 ? add_82582 : array_index_82576[9];
  assign add_82585 = add_82572 + 32'h0000_0001;
  assign array_update_82586[0] = add_81474 == 32'h0000_0000 ? array_update_82584 : array_update_82573[0];
  assign array_update_82586[1] = add_81474 == 32'h0000_0001 ? array_update_82584 : array_update_82573[1];
  assign array_update_82586[2] = add_81474 == 32'h0000_0002 ? array_update_82584 : array_update_82573[2];
  assign array_update_82586[3] = add_81474 == 32'h0000_0003 ? array_update_82584 : array_update_82573[3];
  assign array_update_82586[4] = add_81474 == 32'h0000_0004 ? array_update_82584 : array_update_82573[4];
  assign array_update_82586[5] = add_81474 == 32'h0000_0005 ? array_update_82584 : array_update_82573[5];
  assign array_update_82586[6] = add_81474 == 32'h0000_0006 ? array_update_82584 : array_update_82573[6];
  assign array_update_82586[7] = add_81474 == 32'h0000_0007 ? array_update_82584 : array_update_82573[7];
  assign array_update_82586[8] = add_81474 == 32'h0000_0008 ? array_update_82584 : array_update_82573[8];
  assign array_update_82586[9] = add_81474 == 32'h0000_0009 ? array_update_82584 : array_update_82573[9];
  assign array_index_82588 = array_update_72021[add_82585 > 32'h0000_0009 ? 4'h9 : add_82585[3:0]];
  assign array_index_82589 = array_update_82586[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_82593 = smul32b_32b_x_32b(array_index_81481[add_82585 > 32'h0000_0009 ? 4'h9 : add_82585[3:0]], array_index_82588[add_82557 > 32'h0000_0009 ? 4'h9 : add_82557[3:0]]);
  assign add_82595 = array_index_82589[add_82557 > 32'h0000_0009 ? 4'h9 : add_82557[3:0]] + smul_82593;
  assign array_update_82597[0] = add_82557 == 32'h0000_0000 ? add_82595 : array_index_82589[0];
  assign array_update_82597[1] = add_82557 == 32'h0000_0001 ? add_82595 : array_index_82589[1];
  assign array_update_82597[2] = add_82557 == 32'h0000_0002 ? add_82595 : array_index_82589[2];
  assign array_update_82597[3] = add_82557 == 32'h0000_0003 ? add_82595 : array_index_82589[3];
  assign array_update_82597[4] = add_82557 == 32'h0000_0004 ? add_82595 : array_index_82589[4];
  assign array_update_82597[5] = add_82557 == 32'h0000_0005 ? add_82595 : array_index_82589[5];
  assign array_update_82597[6] = add_82557 == 32'h0000_0006 ? add_82595 : array_index_82589[6];
  assign array_update_82597[7] = add_82557 == 32'h0000_0007 ? add_82595 : array_index_82589[7];
  assign array_update_82597[8] = add_82557 == 32'h0000_0008 ? add_82595 : array_index_82589[8];
  assign array_update_82597[9] = add_82557 == 32'h0000_0009 ? add_82595 : array_index_82589[9];
  assign add_82598 = add_82585 + 32'h0000_0001;
  assign array_update_82599[0] = add_81474 == 32'h0000_0000 ? array_update_82597 : array_update_82586[0];
  assign array_update_82599[1] = add_81474 == 32'h0000_0001 ? array_update_82597 : array_update_82586[1];
  assign array_update_82599[2] = add_81474 == 32'h0000_0002 ? array_update_82597 : array_update_82586[2];
  assign array_update_82599[3] = add_81474 == 32'h0000_0003 ? array_update_82597 : array_update_82586[3];
  assign array_update_82599[4] = add_81474 == 32'h0000_0004 ? array_update_82597 : array_update_82586[4];
  assign array_update_82599[5] = add_81474 == 32'h0000_0005 ? array_update_82597 : array_update_82586[5];
  assign array_update_82599[6] = add_81474 == 32'h0000_0006 ? array_update_82597 : array_update_82586[6];
  assign array_update_82599[7] = add_81474 == 32'h0000_0007 ? array_update_82597 : array_update_82586[7];
  assign array_update_82599[8] = add_81474 == 32'h0000_0008 ? array_update_82597 : array_update_82586[8];
  assign array_update_82599[9] = add_81474 == 32'h0000_0009 ? array_update_82597 : array_update_82586[9];
  assign array_index_82601 = array_update_72021[add_82598 > 32'h0000_0009 ? 4'h9 : add_82598[3:0]];
  assign array_index_82602 = array_update_82599[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_82606 = smul32b_32b_x_32b(array_index_81481[add_82598 > 32'h0000_0009 ? 4'h9 : add_82598[3:0]], array_index_82601[add_82557 > 32'h0000_0009 ? 4'h9 : add_82557[3:0]]);
  assign add_82608 = array_index_82602[add_82557 > 32'h0000_0009 ? 4'h9 : add_82557[3:0]] + smul_82606;
  assign array_update_82610[0] = add_82557 == 32'h0000_0000 ? add_82608 : array_index_82602[0];
  assign array_update_82610[1] = add_82557 == 32'h0000_0001 ? add_82608 : array_index_82602[1];
  assign array_update_82610[2] = add_82557 == 32'h0000_0002 ? add_82608 : array_index_82602[2];
  assign array_update_82610[3] = add_82557 == 32'h0000_0003 ? add_82608 : array_index_82602[3];
  assign array_update_82610[4] = add_82557 == 32'h0000_0004 ? add_82608 : array_index_82602[4];
  assign array_update_82610[5] = add_82557 == 32'h0000_0005 ? add_82608 : array_index_82602[5];
  assign array_update_82610[6] = add_82557 == 32'h0000_0006 ? add_82608 : array_index_82602[6];
  assign array_update_82610[7] = add_82557 == 32'h0000_0007 ? add_82608 : array_index_82602[7];
  assign array_update_82610[8] = add_82557 == 32'h0000_0008 ? add_82608 : array_index_82602[8];
  assign array_update_82610[9] = add_82557 == 32'h0000_0009 ? add_82608 : array_index_82602[9];
  assign add_82611 = add_82598 + 32'h0000_0001;
  assign array_update_82612[0] = add_81474 == 32'h0000_0000 ? array_update_82610 : array_update_82599[0];
  assign array_update_82612[1] = add_81474 == 32'h0000_0001 ? array_update_82610 : array_update_82599[1];
  assign array_update_82612[2] = add_81474 == 32'h0000_0002 ? array_update_82610 : array_update_82599[2];
  assign array_update_82612[3] = add_81474 == 32'h0000_0003 ? array_update_82610 : array_update_82599[3];
  assign array_update_82612[4] = add_81474 == 32'h0000_0004 ? array_update_82610 : array_update_82599[4];
  assign array_update_82612[5] = add_81474 == 32'h0000_0005 ? array_update_82610 : array_update_82599[5];
  assign array_update_82612[6] = add_81474 == 32'h0000_0006 ? array_update_82610 : array_update_82599[6];
  assign array_update_82612[7] = add_81474 == 32'h0000_0007 ? array_update_82610 : array_update_82599[7];
  assign array_update_82612[8] = add_81474 == 32'h0000_0008 ? array_update_82610 : array_update_82599[8];
  assign array_update_82612[9] = add_81474 == 32'h0000_0009 ? array_update_82610 : array_update_82599[9];
  assign array_index_82614 = array_update_72021[add_82611 > 32'h0000_0009 ? 4'h9 : add_82611[3:0]];
  assign array_index_82615 = array_update_82612[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_82619 = smul32b_32b_x_32b(array_index_81481[add_82611 > 32'h0000_0009 ? 4'h9 : add_82611[3:0]], array_index_82614[add_82557 > 32'h0000_0009 ? 4'h9 : add_82557[3:0]]);
  assign add_82621 = array_index_82615[add_82557 > 32'h0000_0009 ? 4'h9 : add_82557[3:0]] + smul_82619;
  assign array_update_82623[0] = add_82557 == 32'h0000_0000 ? add_82621 : array_index_82615[0];
  assign array_update_82623[1] = add_82557 == 32'h0000_0001 ? add_82621 : array_index_82615[1];
  assign array_update_82623[2] = add_82557 == 32'h0000_0002 ? add_82621 : array_index_82615[2];
  assign array_update_82623[3] = add_82557 == 32'h0000_0003 ? add_82621 : array_index_82615[3];
  assign array_update_82623[4] = add_82557 == 32'h0000_0004 ? add_82621 : array_index_82615[4];
  assign array_update_82623[5] = add_82557 == 32'h0000_0005 ? add_82621 : array_index_82615[5];
  assign array_update_82623[6] = add_82557 == 32'h0000_0006 ? add_82621 : array_index_82615[6];
  assign array_update_82623[7] = add_82557 == 32'h0000_0007 ? add_82621 : array_index_82615[7];
  assign array_update_82623[8] = add_82557 == 32'h0000_0008 ? add_82621 : array_index_82615[8];
  assign array_update_82623[9] = add_82557 == 32'h0000_0009 ? add_82621 : array_index_82615[9];
  assign add_82624 = add_82611 + 32'h0000_0001;
  assign array_update_82625[0] = add_81474 == 32'h0000_0000 ? array_update_82623 : array_update_82612[0];
  assign array_update_82625[1] = add_81474 == 32'h0000_0001 ? array_update_82623 : array_update_82612[1];
  assign array_update_82625[2] = add_81474 == 32'h0000_0002 ? array_update_82623 : array_update_82612[2];
  assign array_update_82625[3] = add_81474 == 32'h0000_0003 ? array_update_82623 : array_update_82612[3];
  assign array_update_82625[4] = add_81474 == 32'h0000_0004 ? array_update_82623 : array_update_82612[4];
  assign array_update_82625[5] = add_81474 == 32'h0000_0005 ? array_update_82623 : array_update_82612[5];
  assign array_update_82625[6] = add_81474 == 32'h0000_0006 ? array_update_82623 : array_update_82612[6];
  assign array_update_82625[7] = add_81474 == 32'h0000_0007 ? array_update_82623 : array_update_82612[7];
  assign array_update_82625[8] = add_81474 == 32'h0000_0008 ? array_update_82623 : array_update_82612[8];
  assign array_update_82625[9] = add_81474 == 32'h0000_0009 ? array_update_82623 : array_update_82612[9];
  assign array_index_82627 = array_update_72021[add_82624 > 32'h0000_0009 ? 4'h9 : add_82624[3:0]];
  assign array_index_82628 = array_update_82625[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_82632 = smul32b_32b_x_32b(array_index_81481[add_82624 > 32'h0000_0009 ? 4'h9 : add_82624[3:0]], array_index_82627[add_82557 > 32'h0000_0009 ? 4'h9 : add_82557[3:0]]);
  assign add_82634 = array_index_82628[add_82557 > 32'h0000_0009 ? 4'h9 : add_82557[3:0]] + smul_82632;
  assign array_update_82636[0] = add_82557 == 32'h0000_0000 ? add_82634 : array_index_82628[0];
  assign array_update_82636[1] = add_82557 == 32'h0000_0001 ? add_82634 : array_index_82628[1];
  assign array_update_82636[2] = add_82557 == 32'h0000_0002 ? add_82634 : array_index_82628[2];
  assign array_update_82636[3] = add_82557 == 32'h0000_0003 ? add_82634 : array_index_82628[3];
  assign array_update_82636[4] = add_82557 == 32'h0000_0004 ? add_82634 : array_index_82628[4];
  assign array_update_82636[5] = add_82557 == 32'h0000_0005 ? add_82634 : array_index_82628[5];
  assign array_update_82636[6] = add_82557 == 32'h0000_0006 ? add_82634 : array_index_82628[6];
  assign array_update_82636[7] = add_82557 == 32'h0000_0007 ? add_82634 : array_index_82628[7];
  assign array_update_82636[8] = add_82557 == 32'h0000_0008 ? add_82634 : array_index_82628[8];
  assign array_update_82636[9] = add_82557 == 32'h0000_0009 ? add_82634 : array_index_82628[9];
  assign add_82637 = add_82624 + 32'h0000_0001;
  assign array_update_82638[0] = add_81474 == 32'h0000_0000 ? array_update_82636 : array_update_82625[0];
  assign array_update_82638[1] = add_81474 == 32'h0000_0001 ? array_update_82636 : array_update_82625[1];
  assign array_update_82638[2] = add_81474 == 32'h0000_0002 ? array_update_82636 : array_update_82625[2];
  assign array_update_82638[3] = add_81474 == 32'h0000_0003 ? array_update_82636 : array_update_82625[3];
  assign array_update_82638[4] = add_81474 == 32'h0000_0004 ? array_update_82636 : array_update_82625[4];
  assign array_update_82638[5] = add_81474 == 32'h0000_0005 ? array_update_82636 : array_update_82625[5];
  assign array_update_82638[6] = add_81474 == 32'h0000_0006 ? array_update_82636 : array_update_82625[6];
  assign array_update_82638[7] = add_81474 == 32'h0000_0007 ? array_update_82636 : array_update_82625[7];
  assign array_update_82638[8] = add_81474 == 32'h0000_0008 ? array_update_82636 : array_update_82625[8];
  assign array_update_82638[9] = add_81474 == 32'h0000_0009 ? array_update_82636 : array_update_82625[9];
  assign array_index_82640 = array_update_72021[add_82637 > 32'h0000_0009 ? 4'h9 : add_82637[3:0]];
  assign array_index_82641 = array_update_82638[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_82645 = smul32b_32b_x_32b(array_index_81481[add_82637 > 32'h0000_0009 ? 4'h9 : add_82637[3:0]], array_index_82640[add_82557 > 32'h0000_0009 ? 4'h9 : add_82557[3:0]]);
  assign add_82647 = array_index_82641[add_82557 > 32'h0000_0009 ? 4'h9 : add_82557[3:0]] + smul_82645;
  assign array_update_82649[0] = add_82557 == 32'h0000_0000 ? add_82647 : array_index_82641[0];
  assign array_update_82649[1] = add_82557 == 32'h0000_0001 ? add_82647 : array_index_82641[1];
  assign array_update_82649[2] = add_82557 == 32'h0000_0002 ? add_82647 : array_index_82641[2];
  assign array_update_82649[3] = add_82557 == 32'h0000_0003 ? add_82647 : array_index_82641[3];
  assign array_update_82649[4] = add_82557 == 32'h0000_0004 ? add_82647 : array_index_82641[4];
  assign array_update_82649[5] = add_82557 == 32'h0000_0005 ? add_82647 : array_index_82641[5];
  assign array_update_82649[6] = add_82557 == 32'h0000_0006 ? add_82647 : array_index_82641[6];
  assign array_update_82649[7] = add_82557 == 32'h0000_0007 ? add_82647 : array_index_82641[7];
  assign array_update_82649[8] = add_82557 == 32'h0000_0008 ? add_82647 : array_index_82641[8];
  assign array_update_82649[9] = add_82557 == 32'h0000_0009 ? add_82647 : array_index_82641[9];
  assign add_82650 = add_82637 + 32'h0000_0001;
  assign array_update_82651[0] = add_81474 == 32'h0000_0000 ? array_update_82649 : array_update_82638[0];
  assign array_update_82651[1] = add_81474 == 32'h0000_0001 ? array_update_82649 : array_update_82638[1];
  assign array_update_82651[2] = add_81474 == 32'h0000_0002 ? array_update_82649 : array_update_82638[2];
  assign array_update_82651[3] = add_81474 == 32'h0000_0003 ? array_update_82649 : array_update_82638[3];
  assign array_update_82651[4] = add_81474 == 32'h0000_0004 ? array_update_82649 : array_update_82638[4];
  assign array_update_82651[5] = add_81474 == 32'h0000_0005 ? array_update_82649 : array_update_82638[5];
  assign array_update_82651[6] = add_81474 == 32'h0000_0006 ? array_update_82649 : array_update_82638[6];
  assign array_update_82651[7] = add_81474 == 32'h0000_0007 ? array_update_82649 : array_update_82638[7];
  assign array_update_82651[8] = add_81474 == 32'h0000_0008 ? array_update_82649 : array_update_82638[8];
  assign array_update_82651[9] = add_81474 == 32'h0000_0009 ? array_update_82649 : array_update_82638[9];
  assign array_index_82653 = array_update_72021[add_82650 > 32'h0000_0009 ? 4'h9 : add_82650[3:0]];
  assign array_index_82654 = array_update_82651[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_82658 = smul32b_32b_x_32b(array_index_81481[add_82650 > 32'h0000_0009 ? 4'h9 : add_82650[3:0]], array_index_82653[add_82557 > 32'h0000_0009 ? 4'h9 : add_82557[3:0]]);
  assign add_82660 = array_index_82654[add_82557 > 32'h0000_0009 ? 4'h9 : add_82557[3:0]] + smul_82658;
  assign array_update_82662[0] = add_82557 == 32'h0000_0000 ? add_82660 : array_index_82654[0];
  assign array_update_82662[1] = add_82557 == 32'h0000_0001 ? add_82660 : array_index_82654[1];
  assign array_update_82662[2] = add_82557 == 32'h0000_0002 ? add_82660 : array_index_82654[2];
  assign array_update_82662[3] = add_82557 == 32'h0000_0003 ? add_82660 : array_index_82654[3];
  assign array_update_82662[4] = add_82557 == 32'h0000_0004 ? add_82660 : array_index_82654[4];
  assign array_update_82662[5] = add_82557 == 32'h0000_0005 ? add_82660 : array_index_82654[5];
  assign array_update_82662[6] = add_82557 == 32'h0000_0006 ? add_82660 : array_index_82654[6];
  assign array_update_82662[7] = add_82557 == 32'h0000_0007 ? add_82660 : array_index_82654[7];
  assign array_update_82662[8] = add_82557 == 32'h0000_0008 ? add_82660 : array_index_82654[8];
  assign array_update_82662[9] = add_82557 == 32'h0000_0009 ? add_82660 : array_index_82654[9];
  assign add_82663 = add_82650 + 32'h0000_0001;
  assign array_update_82664[0] = add_81474 == 32'h0000_0000 ? array_update_82662 : array_update_82651[0];
  assign array_update_82664[1] = add_81474 == 32'h0000_0001 ? array_update_82662 : array_update_82651[1];
  assign array_update_82664[2] = add_81474 == 32'h0000_0002 ? array_update_82662 : array_update_82651[2];
  assign array_update_82664[3] = add_81474 == 32'h0000_0003 ? array_update_82662 : array_update_82651[3];
  assign array_update_82664[4] = add_81474 == 32'h0000_0004 ? array_update_82662 : array_update_82651[4];
  assign array_update_82664[5] = add_81474 == 32'h0000_0005 ? array_update_82662 : array_update_82651[5];
  assign array_update_82664[6] = add_81474 == 32'h0000_0006 ? array_update_82662 : array_update_82651[6];
  assign array_update_82664[7] = add_81474 == 32'h0000_0007 ? array_update_82662 : array_update_82651[7];
  assign array_update_82664[8] = add_81474 == 32'h0000_0008 ? array_update_82662 : array_update_82651[8];
  assign array_update_82664[9] = add_81474 == 32'h0000_0009 ? array_update_82662 : array_update_82651[9];
  assign array_index_82666 = array_update_72021[add_82663 > 32'h0000_0009 ? 4'h9 : add_82663[3:0]];
  assign array_index_82667 = array_update_82664[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_82671 = smul32b_32b_x_32b(array_index_81481[add_82663 > 32'h0000_0009 ? 4'h9 : add_82663[3:0]], array_index_82666[add_82557 > 32'h0000_0009 ? 4'h9 : add_82557[3:0]]);
  assign add_82673 = array_index_82667[add_82557 > 32'h0000_0009 ? 4'h9 : add_82557[3:0]] + smul_82671;
  assign array_update_82675[0] = add_82557 == 32'h0000_0000 ? add_82673 : array_index_82667[0];
  assign array_update_82675[1] = add_82557 == 32'h0000_0001 ? add_82673 : array_index_82667[1];
  assign array_update_82675[2] = add_82557 == 32'h0000_0002 ? add_82673 : array_index_82667[2];
  assign array_update_82675[3] = add_82557 == 32'h0000_0003 ? add_82673 : array_index_82667[3];
  assign array_update_82675[4] = add_82557 == 32'h0000_0004 ? add_82673 : array_index_82667[4];
  assign array_update_82675[5] = add_82557 == 32'h0000_0005 ? add_82673 : array_index_82667[5];
  assign array_update_82675[6] = add_82557 == 32'h0000_0006 ? add_82673 : array_index_82667[6];
  assign array_update_82675[7] = add_82557 == 32'h0000_0007 ? add_82673 : array_index_82667[7];
  assign array_update_82675[8] = add_82557 == 32'h0000_0008 ? add_82673 : array_index_82667[8];
  assign array_update_82675[9] = add_82557 == 32'h0000_0009 ? add_82673 : array_index_82667[9];
  assign add_82676 = add_82663 + 32'h0000_0001;
  assign array_update_82677[0] = add_81474 == 32'h0000_0000 ? array_update_82675 : array_update_82664[0];
  assign array_update_82677[1] = add_81474 == 32'h0000_0001 ? array_update_82675 : array_update_82664[1];
  assign array_update_82677[2] = add_81474 == 32'h0000_0002 ? array_update_82675 : array_update_82664[2];
  assign array_update_82677[3] = add_81474 == 32'h0000_0003 ? array_update_82675 : array_update_82664[3];
  assign array_update_82677[4] = add_81474 == 32'h0000_0004 ? array_update_82675 : array_update_82664[4];
  assign array_update_82677[5] = add_81474 == 32'h0000_0005 ? array_update_82675 : array_update_82664[5];
  assign array_update_82677[6] = add_81474 == 32'h0000_0006 ? array_update_82675 : array_update_82664[6];
  assign array_update_82677[7] = add_81474 == 32'h0000_0007 ? array_update_82675 : array_update_82664[7];
  assign array_update_82677[8] = add_81474 == 32'h0000_0008 ? array_update_82675 : array_update_82664[8];
  assign array_update_82677[9] = add_81474 == 32'h0000_0009 ? array_update_82675 : array_update_82664[9];
  assign array_index_82679 = array_update_72021[add_82676 > 32'h0000_0009 ? 4'h9 : add_82676[3:0]];
  assign array_index_82680 = array_update_82677[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_82684 = smul32b_32b_x_32b(array_index_81481[add_82676 > 32'h0000_0009 ? 4'h9 : add_82676[3:0]], array_index_82679[add_82557 > 32'h0000_0009 ? 4'h9 : add_82557[3:0]]);
  assign add_82686 = array_index_82680[add_82557 > 32'h0000_0009 ? 4'h9 : add_82557[3:0]] + smul_82684;
  assign array_update_82687[0] = add_82557 == 32'h0000_0000 ? add_82686 : array_index_82680[0];
  assign array_update_82687[1] = add_82557 == 32'h0000_0001 ? add_82686 : array_index_82680[1];
  assign array_update_82687[2] = add_82557 == 32'h0000_0002 ? add_82686 : array_index_82680[2];
  assign array_update_82687[3] = add_82557 == 32'h0000_0003 ? add_82686 : array_index_82680[3];
  assign array_update_82687[4] = add_82557 == 32'h0000_0004 ? add_82686 : array_index_82680[4];
  assign array_update_82687[5] = add_82557 == 32'h0000_0005 ? add_82686 : array_index_82680[5];
  assign array_update_82687[6] = add_82557 == 32'h0000_0006 ? add_82686 : array_index_82680[6];
  assign array_update_82687[7] = add_82557 == 32'h0000_0007 ? add_82686 : array_index_82680[7];
  assign array_update_82687[8] = add_82557 == 32'h0000_0008 ? add_82686 : array_index_82680[8];
  assign array_update_82687[9] = add_82557 == 32'h0000_0009 ? add_82686 : array_index_82680[9];
  assign array_update_82688[0] = add_81474 == 32'h0000_0000 ? array_update_82687 : array_update_82677[0];
  assign array_update_82688[1] = add_81474 == 32'h0000_0001 ? array_update_82687 : array_update_82677[1];
  assign array_update_82688[2] = add_81474 == 32'h0000_0002 ? array_update_82687 : array_update_82677[2];
  assign array_update_82688[3] = add_81474 == 32'h0000_0003 ? array_update_82687 : array_update_82677[3];
  assign array_update_82688[4] = add_81474 == 32'h0000_0004 ? array_update_82687 : array_update_82677[4];
  assign array_update_82688[5] = add_81474 == 32'h0000_0005 ? array_update_82687 : array_update_82677[5];
  assign array_update_82688[6] = add_81474 == 32'h0000_0006 ? array_update_82687 : array_update_82677[6];
  assign array_update_82688[7] = add_81474 == 32'h0000_0007 ? array_update_82687 : array_update_82677[7];
  assign array_update_82688[8] = add_81474 == 32'h0000_0008 ? array_update_82687 : array_update_82677[8];
  assign array_update_82688[9] = add_81474 == 32'h0000_0009 ? array_update_82687 : array_update_82677[9];
  assign array_index_82690 = array_update_82688[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign add_82692 = add_82557 + 32'h0000_0001;
  assign array_update_82693[0] = add_82692 == 32'h0000_0000 ? 32'h0000_0000 : array_index_82690[0];
  assign array_update_82693[1] = add_82692 == 32'h0000_0001 ? 32'h0000_0000 : array_index_82690[1];
  assign array_update_82693[2] = add_82692 == 32'h0000_0002 ? 32'h0000_0000 : array_index_82690[2];
  assign array_update_82693[3] = add_82692 == 32'h0000_0003 ? 32'h0000_0000 : array_index_82690[3];
  assign array_update_82693[4] = add_82692 == 32'h0000_0004 ? 32'h0000_0000 : array_index_82690[4];
  assign array_update_82693[5] = add_82692 == 32'h0000_0005 ? 32'h0000_0000 : array_index_82690[5];
  assign array_update_82693[6] = add_82692 == 32'h0000_0006 ? 32'h0000_0000 : array_index_82690[6];
  assign array_update_82693[7] = add_82692 == 32'h0000_0007 ? 32'h0000_0000 : array_index_82690[7];
  assign array_update_82693[8] = add_82692 == 32'h0000_0008 ? 32'h0000_0000 : array_index_82690[8];
  assign array_update_82693[9] = add_82692 == 32'h0000_0009 ? 32'h0000_0000 : array_index_82690[9];
  assign literal_82694 = 32'h0000_0000;
  assign array_update_82695[0] = add_81474 == 32'h0000_0000 ? array_update_82693 : array_update_82688[0];
  assign array_update_82695[1] = add_81474 == 32'h0000_0001 ? array_update_82693 : array_update_82688[1];
  assign array_update_82695[2] = add_81474 == 32'h0000_0002 ? array_update_82693 : array_update_82688[2];
  assign array_update_82695[3] = add_81474 == 32'h0000_0003 ? array_update_82693 : array_update_82688[3];
  assign array_update_82695[4] = add_81474 == 32'h0000_0004 ? array_update_82693 : array_update_82688[4];
  assign array_update_82695[5] = add_81474 == 32'h0000_0005 ? array_update_82693 : array_update_82688[5];
  assign array_update_82695[6] = add_81474 == 32'h0000_0006 ? array_update_82693 : array_update_82688[6];
  assign array_update_82695[7] = add_81474 == 32'h0000_0007 ? array_update_82693 : array_update_82688[7];
  assign array_update_82695[8] = add_81474 == 32'h0000_0008 ? array_update_82693 : array_update_82688[8];
  assign array_update_82695[9] = add_81474 == 32'h0000_0009 ? array_update_82693 : array_update_82688[9];
  assign array_index_82697 = array_update_72021[literal_82694 > 32'h0000_0009 ? 4'h9 : literal_82694[3:0]];
  assign array_index_82698 = array_update_82695[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_82702 = smul32b_32b_x_32b(array_index_81481[literal_82694 > 32'h0000_0009 ? 4'h9 : literal_82694[3:0]], array_index_82697[add_82692 > 32'h0000_0009 ? 4'h9 : add_82692[3:0]]);
  assign add_82704 = array_index_82698[add_82692 > 32'h0000_0009 ? 4'h9 : add_82692[3:0]] + smul_82702;
  assign array_update_82706[0] = add_82692 == 32'h0000_0000 ? add_82704 : array_index_82698[0];
  assign array_update_82706[1] = add_82692 == 32'h0000_0001 ? add_82704 : array_index_82698[1];
  assign array_update_82706[2] = add_82692 == 32'h0000_0002 ? add_82704 : array_index_82698[2];
  assign array_update_82706[3] = add_82692 == 32'h0000_0003 ? add_82704 : array_index_82698[3];
  assign array_update_82706[4] = add_82692 == 32'h0000_0004 ? add_82704 : array_index_82698[4];
  assign array_update_82706[5] = add_82692 == 32'h0000_0005 ? add_82704 : array_index_82698[5];
  assign array_update_82706[6] = add_82692 == 32'h0000_0006 ? add_82704 : array_index_82698[6];
  assign array_update_82706[7] = add_82692 == 32'h0000_0007 ? add_82704 : array_index_82698[7];
  assign array_update_82706[8] = add_82692 == 32'h0000_0008 ? add_82704 : array_index_82698[8];
  assign array_update_82706[9] = add_82692 == 32'h0000_0009 ? add_82704 : array_index_82698[9];
  assign add_82707 = literal_82694 + 32'h0000_0001;
  assign array_update_82708[0] = add_81474 == 32'h0000_0000 ? array_update_82706 : array_update_82695[0];
  assign array_update_82708[1] = add_81474 == 32'h0000_0001 ? array_update_82706 : array_update_82695[1];
  assign array_update_82708[2] = add_81474 == 32'h0000_0002 ? array_update_82706 : array_update_82695[2];
  assign array_update_82708[3] = add_81474 == 32'h0000_0003 ? array_update_82706 : array_update_82695[3];
  assign array_update_82708[4] = add_81474 == 32'h0000_0004 ? array_update_82706 : array_update_82695[4];
  assign array_update_82708[5] = add_81474 == 32'h0000_0005 ? array_update_82706 : array_update_82695[5];
  assign array_update_82708[6] = add_81474 == 32'h0000_0006 ? array_update_82706 : array_update_82695[6];
  assign array_update_82708[7] = add_81474 == 32'h0000_0007 ? array_update_82706 : array_update_82695[7];
  assign array_update_82708[8] = add_81474 == 32'h0000_0008 ? array_update_82706 : array_update_82695[8];
  assign array_update_82708[9] = add_81474 == 32'h0000_0009 ? array_update_82706 : array_update_82695[9];
  assign array_index_82710 = array_update_72021[add_82707 > 32'h0000_0009 ? 4'h9 : add_82707[3:0]];
  assign array_index_82711 = array_update_82708[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_82715 = smul32b_32b_x_32b(array_index_81481[add_82707 > 32'h0000_0009 ? 4'h9 : add_82707[3:0]], array_index_82710[add_82692 > 32'h0000_0009 ? 4'h9 : add_82692[3:0]]);
  assign add_82717 = array_index_82711[add_82692 > 32'h0000_0009 ? 4'h9 : add_82692[3:0]] + smul_82715;
  assign array_update_82719[0] = add_82692 == 32'h0000_0000 ? add_82717 : array_index_82711[0];
  assign array_update_82719[1] = add_82692 == 32'h0000_0001 ? add_82717 : array_index_82711[1];
  assign array_update_82719[2] = add_82692 == 32'h0000_0002 ? add_82717 : array_index_82711[2];
  assign array_update_82719[3] = add_82692 == 32'h0000_0003 ? add_82717 : array_index_82711[3];
  assign array_update_82719[4] = add_82692 == 32'h0000_0004 ? add_82717 : array_index_82711[4];
  assign array_update_82719[5] = add_82692 == 32'h0000_0005 ? add_82717 : array_index_82711[5];
  assign array_update_82719[6] = add_82692 == 32'h0000_0006 ? add_82717 : array_index_82711[6];
  assign array_update_82719[7] = add_82692 == 32'h0000_0007 ? add_82717 : array_index_82711[7];
  assign array_update_82719[8] = add_82692 == 32'h0000_0008 ? add_82717 : array_index_82711[8];
  assign array_update_82719[9] = add_82692 == 32'h0000_0009 ? add_82717 : array_index_82711[9];
  assign add_82720 = add_82707 + 32'h0000_0001;
  assign array_update_82721[0] = add_81474 == 32'h0000_0000 ? array_update_82719 : array_update_82708[0];
  assign array_update_82721[1] = add_81474 == 32'h0000_0001 ? array_update_82719 : array_update_82708[1];
  assign array_update_82721[2] = add_81474 == 32'h0000_0002 ? array_update_82719 : array_update_82708[2];
  assign array_update_82721[3] = add_81474 == 32'h0000_0003 ? array_update_82719 : array_update_82708[3];
  assign array_update_82721[4] = add_81474 == 32'h0000_0004 ? array_update_82719 : array_update_82708[4];
  assign array_update_82721[5] = add_81474 == 32'h0000_0005 ? array_update_82719 : array_update_82708[5];
  assign array_update_82721[6] = add_81474 == 32'h0000_0006 ? array_update_82719 : array_update_82708[6];
  assign array_update_82721[7] = add_81474 == 32'h0000_0007 ? array_update_82719 : array_update_82708[7];
  assign array_update_82721[8] = add_81474 == 32'h0000_0008 ? array_update_82719 : array_update_82708[8];
  assign array_update_82721[9] = add_81474 == 32'h0000_0009 ? array_update_82719 : array_update_82708[9];
  assign array_index_82723 = array_update_72021[add_82720 > 32'h0000_0009 ? 4'h9 : add_82720[3:0]];
  assign array_index_82724 = array_update_82721[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_82728 = smul32b_32b_x_32b(array_index_81481[add_82720 > 32'h0000_0009 ? 4'h9 : add_82720[3:0]], array_index_82723[add_82692 > 32'h0000_0009 ? 4'h9 : add_82692[3:0]]);
  assign add_82730 = array_index_82724[add_82692 > 32'h0000_0009 ? 4'h9 : add_82692[3:0]] + smul_82728;
  assign array_update_82732[0] = add_82692 == 32'h0000_0000 ? add_82730 : array_index_82724[0];
  assign array_update_82732[1] = add_82692 == 32'h0000_0001 ? add_82730 : array_index_82724[1];
  assign array_update_82732[2] = add_82692 == 32'h0000_0002 ? add_82730 : array_index_82724[2];
  assign array_update_82732[3] = add_82692 == 32'h0000_0003 ? add_82730 : array_index_82724[3];
  assign array_update_82732[4] = add_82692 == 32'h0000_0004 ? add_82730 : array_index_82724[4];
  assign array_update_82732[5] = add_82692 == 32'h0000_0005 ? add_82730 : array_index_82724[5];
  assign array_update_82732[6] = add_82692 == 32'h0000_0006 ? add_82730 : array_index_82724[6];
  assign array_update_82732[7] = add_82692 == 32'h0000_0007 ? add_82730 : array_index_82724[7];
  assign array_update_82732[8] = add_82692 == 32'h0000_0008 ? add_82730 : array_index_82724[8];
  assign array_update_82732[9] = add_82692 == 32'h0000_0009 ? add_82730 : array_index_82724[9];
  assign add_82733 = add_82720 + 32'h0000_0001;
  assign array_update_82734[0] = add_81474 == 32'h0000_0000 ? array_update_82732 : array_update_82721[0];
  assign array_update_82734[1] = add_81474 == 32'h0000_0001 ? array_update_82732 : array_update_82721[1];
  assign array_update_82734[2] = add_81474 == 32'h0000_0002 ? array_update_82732 : array_update_82721[2];
  assign array_update_82734[3] = add_81474 == 32'h0000_0003 ? array_update_82732 : array_update_82721[3];
  assign array_update_82734[4] = add_81474 == 32'h0000_0004 ? array_update_82732 : array_update_82721[4];
  assign array_update_82734[5] = add_81474 == 32'h0000_0005 ? array_update_82732 : array_update_82721[5];
  assign array_update_82734[6] = add_81474 == 32'h0000_0006 ? array_update_82732 : array_update_82721[6];
  assign array_update_82734[7] = add_81474 == 32'h0000_0007 ? array_update_82732 : array_update_82721[7];
  assign array_update_82734[8] = add_81474 == 32'h0000_0008 ? array_update_82732 : array_update_82721[8];
  assign array_update_82734[9] = add_81474 == 32'h0000_0009 ? array_update_82732 : array_update_82721[9];
  assign array_index_82736 = array_update_72021[add_82733 > 32'h0000_0009 ? 4'h9 : add_82733[3:0]];
  assign array_index_82737 = array_update_82734[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_82741 = smul32b_32b_x_32b(array_index_81481[add_82733 > 32'h0000_0009 ? 4'h9 : add_82733[3:0]], array_index_82736[add_82692 > 32'h0000_0009 ? 4'h9 : add_82692[3:0]]);
  assign add_82743 = array_index_82737[add_82692 > 32'h0000_0009 ? 4'h9 : add_82692[3:0]] + smul_82741;
  assign array_update_82745[0] = add_82692 == 32'h0000_0000 ? add_82743 : array_index_82737[0];
  assign array_update_82745[1] = add_82692 == 32'h0000_0001 ? add_82743 : array_index_82737[1];
  assign array_update_82745[2] = add_82692 == 32'h0000_0002 ? add_82743 : array_index_82737[2];
  assign array_update_82745[3] = add_82692 == 32'h0000_0003 ? add_82743 : array_index_82737[3];
  assign array_update_82745[4] = add_82692 == 32'h0000_0004 ? add_82743 : array_index_82737[4];
  assign array_update_82745[5] = add_82692 == 32'h0000_0005 ? add_82743 : array_index_82737[5];
  assign array_update_82745[6] = add_82692 == 32'h0000_0006 ? add_82743 : array_index_82737[6];
  assign array_update_82745[7] = add_82692 == 32'h0000_0007 ? add_82743 : array_index_82737[7];
  assign array_update_82745[8] = add_82692 == 32'h0000_0008 ? add_82743 : array_index_82737[8];
  assign array_update_82745[9] = add_82692 == 32'h0000_0009 ? add_82743 : array_index_82737[9];
  assign add_82746 = add_82733 + 32'h0000_0001;
  assign array_update_82747[0] = add_81474 == 32'h0000_0000 ? array_update_82745 : array_update_82734[0];
  assign array_update_82747[1] = add_81474 == 32'h0000_0001 ? array_update_82745 : array_update_82734[1];
  assign array_update_82747[2] = add_81474 == 32'h0000_0002 ? array_update_82745 : array_update_82734[2];
  assign array_update_82747[3] = add_81474 == 32'h0000_0003 ? array_update_82745 : array_update_82734[3];
  assign array_update_82747[4] = add_81474 == 32'h0000_0004 ? array_update_82745 : array_update_82734[4];
  assign array_update_82747[5] = add_81474 == 32'h0000_0005 ? array_update_82745 : array_update_82734[5];
  assign array_update_82747[6] = add_81474 == 32'h0000_0006 ? array_update_82745 : array_update_82734[6];
  assign array_update_82747[7] = add_81474 == 32'h0000_0007 ? array_update_82745 : array_update_82734[7];
  assign array_update_82747[8] = add_81474 == 32'h0000_0008 ? array_update_82745 : array_update_82734[8];
  assign array_update_82747[9] = add_81474 == 32'h0000_0009 ? array_update_82745 : array_update_82734[9];
  assign array_index_82749 = array_update_72021[add_82746 > 32'h0000_0009 ? 4'h9 : add_82746[3:0]];
  assign array_index_82750 = array_update_82747[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_82754 = smul32b_32b_x_32b(array_index_81481[add_82746 > 32'h0000_0009 ? 4'h9 : add_82746[3:0]], array_index_82749[add_82692 > 32'h0000_0009 ? 4'h9 : add_82692[3:0]]);
  assign add_82756 = array_index_82750[add_82692 > 32'h0000_0009 ? 4'h9 : add_82692[3:0]] + smul_82754;
  assign array_update_82758[0] = add_82692 == 32'h0000_0000 ? add_82756 : array_index_82750[0];
  assign array_update_82758[1] = add_82692 == 32'h0000_0001 ? add_82756 : array_index_82750[1];
  assign array_update_82758[2] = add_82692 == 32'h0000_0002 ? add_82756 : array_index_82750[2];
  assign array_update_82758[3] = add_82692 == 32'h0000_0003 ? add_82756 : array_index_82750[3];
  assign array_update_82758[4] = add_82692 == 32'h0000_0004 ? add_82756 : array_index_82750[4];
  assign array_update_82758[5] = add_82692 == 32'h0000_0005 ? add_82756 : array_index_82750[5];
  assign array_update_82758[6] = add_82692 == 32'h0000_0006 ? add_82756 : array_index_82750[6];
  assign array_update_82758[7] = add_82692 == 32'h0000_0007 ? add_82756 : array_index_82750[7];
  assign array_update_82758[8] = add_82692 == 32'h0000_0008 ? add_82756 : array_index_82750[8];
  assign array_update_82758[9] = add_82692 == 32'h0000_0009 ? add_82756 : array_index_82750[9];
  assign add_82759 = add_82746 + 32'h0000_0001;
  assign array_update_82760[0] = add_81474 == 32'h0000_0000 ? array_update_82758 : array_update_82747[0];
  assign array_update_82760[1] = add_81474 == 32'h0000_0001 ? array_update_82758 : array_update_82747[1];
  assign array_update_82760[2] = add_81474 == 32'h0000_0002 ? array_update_82758 : array_update_82747[2];
  assign array_update_82760[3] = add_81474 == 32'h0000_0003 ? array_update_82758 : array_update_82747[3];
  assign array_update_82760[4] = add_81474 == 32'h0000_0004 ? array_update_82758 : array_update_82747[4];
  assign array_update_82760[5] = add_81474 == 32'h0000_0005 ? array_update_82758 : array_update_82747[5];
  assign array_update_82760[6] = add_81474 == 32'h0000_0006 ? array_update_82758 : array_update_82747[6];
  assign array_update_82760[7] = add_81474 == 32'h0000_0007 ? array_update_82758 : array_update_82747[7];
  assign array_update_82760[8] = add_81474 == 32'h0000_0008 ? array_update_82758 : array_update_82747[8];
  assign array_update_82760[9] = add_81474 == 32'h0000_0009 ? array_update_82758 : array_update_82747[9];
  assign array_index_82762 = array_update_72021[add_82759 > 32'h0000_0009 ? 4'h9 : add_82759[3:0]];
  assign array_index_82763 = array_update_82760[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_82767 = smul32b_32b_x_32b(array_index_81481[add_82759 > 32'h0000_0009 ? 4'h9 : add_82759[3:0]], array_index_82762[add_82692 > 32'h0000_0009 ? 4'h9 : add_82692[3:0]]);
  assign add_82769 = array_index_82763[add_82692 > 32'h0000_0009 ? 4'h9 : add_82692[3:0]] + smul_82767;
  assign array_update_82771[0] = add_82692 == 32'h0000_0000 ? add_82769 : array_index_82763[0];
  assign array_update_82771[1] = add_82692 == 32'h0000_0001 ? add_82769 : array_index_82763[1];
  assign array_update_82771[2] = add_82692 == 32'h0000_0002 ? add_82769 : array_index_82763[2];
  assign array_update_82771[3] = add_82692 == 32'h0000_0003 ? add_82769 : array_index_82763[3];
  assign array_update_82771[4] = add_82692 == 32'h0000_0004 ? add_82769 : array_index_82763[4];
  assign array_update_82771[5] = add_82692 == 32'h0000_0005 ? add_82769 : array_index_82763[5];
  assign array_update_82771[6] = add_82692 == 32'h0000_0006 ? add_82769 : array_index_82763[6];
  assign array_update_82771[7] = add_82692 == 32'h0000_0007 ? add_82769 : array_index_82763[7];
  assign array_update_82771[8] = add_82692 == 32'h0000_0008 ? add_82769 : array_index_82763[8];
  assign array_update_82771[9] = add_82692 == 32'h0000_0009 ? add_82769 : array_index_82763[9];
  assign add_82772 = add_82759 + 32'h0000_0001;
  assign array_update_82773[0] = add_81474 == 32'h0000_0000 ? array_update_82771 : array_update_82760[0];
  assign array_update_82773[1] = add_81474 == 32'h0000_0001 ? array_update_82771 : array_update_82760[1];
  assign array_update_82773[2] = add_81474 == 32'h0000_0002 ? array_update_82771 : array_update_82760[2];
  assign array_update_82773[3] = add_81474 == 32'h0000_0003 ? array_update_82771 : array_update_82760[3];
  assign array_update_82773[4] = add_81474 == 32'h0000_0004 ? array_update_82771 : array_update_82760[4];
  assign array_update_82773[5] = add_81474 == 32'h0000_0005 ? array_update_82771 : array_update_82760[5];
  assign array_update_82773[6] = add_81474 == 32'h0000_0006 ? array_update_82771 : array_update_82760[6];
  assign array_update_82773[7] = add_81474 == 32'h0000_0007 ? array_update_82771 : array_update_82760[7];
  assign array_update_82773[8] = add_81474 == 32'h0000_0008 ? array_update_82771 : array_update_82760[8];
  assign array_update_82773[9] = add_81474 == 32'h0000_0009 ? array_update_82771 : array_update_82760[9];
  assign array_index_82775 = array_update_72021[add_82772 > 32'h0000_0009 ? 4'h9 : add_82772[3:0]];
  assign array_index_82776 = array_update_82773[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_82780 = smul32b_32b_x_32b(array_index_81481[add_82772 > 32'h0000_0009 ? 4'h9 : add_82772[3:0]], array_index_82775[add_82692 > 32'h0000_0009 ? 4'h9 : add_82692[3:0]]);
  assign add_82782 = array_index_82776[add_82692 > 32'h0000_0009 ? 4'h9 : add_82692[3:0]] + smul_82780;
  assign array_update_82784[0] = add_82692 == 32'h0000_0000 ? add_82782 : array_index_82776[0];
  assign array_update_82784[1] = add_82692 == 32'h0000_0001 ? add_82782 : array_index_82776[1];
  assign array_update_82784[2] = add_82692 == 32'h0000_0002 ? add_82782 : array_index_82776[2];
  assign array_update_82784[3] = add_82692 == 32'h0000_0003 ? add_82782 : array_index_82776[3];
  assign array_update_82784[4] = add_82692 == 32'h0000_0004 ? add_82782 : array_index_82776[4];
  assign array_update_82784[5] = add_82692 == 32'h0000_0005 ? add_82782 : array_index_82776[5];
  assign array_update_82784[6] = add_82692 == 32'h0000_0006 ? add_82782 : array_index_82776[6];
  assign array_update_82784[7] = add_82692 == 32'h0000_0007 ? add_82782 : array_index_82776[7];
  assign array_update_82784[8] = add_82692 == 32'h0000_0008 ? add_82782 : array_index_82776[8];
  assign array_update_82784[9] = add_82692 == 32'h0000_0009 ? add_82782 : array_index_82776[9];
  assign add_82785 = add_82772 + 32'h0000_0001;
  assign array_update_82786[0] = add_81474 == 32'h0000_0000 ? array_update_82784 : array_update_82773[0];
  assign array_update_82786[1] = add_81474 == 32'h0000_0001 ? array_update_82784 : array_update_82773[1];
  assign array_update_82786[2] = add_81474 == 32'h0000_0002 ? array_update_82784 : array_update_82773[2];
  assign array_update_82786[3] = add_81474 == 32'h0000_0003 ? array_update_82784 : array_update_82773[3];
  assign array_update_82786[4] = add_81474 == 32'h0000_0004 ? array_update_82784 : array_update_82773[4];
  assign array_update_82786[5] = add_81474 == 32'h0000_0005 ? array_update_82784 : array_update_82773[5];
  assign array_update_82786[6] = add_81474 == 32'h0000_0006 ? array_update_82784 : array_update_82773[6];
  assign array_update_82786[7] = add_81474 == 32'h0000_0007 ? array_update_82784 : array_update_82773[7];
  assign array_update_82786[8] = add_81474 == 32'h0000_0008 ? array_update_82784 : array_update_82773[8];
  assign array_update_82786[9] = add_81474 == 32'h0000_0009 ? array_update_82784 : array_update_82773[9];
  assign array_index_82788 = array_update_72021[add_82785 > 32'h0000_0009 ? 4'h9 : add_82785[3:0]];
  assign array_index_82789 = array_update_82786[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_82793 = smul32b_32b_x_32b(array_index_81481[add_82785 > 32'h0000_0009 ? 4'h9 : add_82785[3:0]], array_index_82788[add_82692 > 32'h0000_0009 ? 4'h9 : add_82692[3:0]]);
  assign add_82795 = array_index_82789[add_82692 > 32'h0000_0009 ? 4'h9 : add_82692[3:0]] + smul_82793;
  assign array_update_82797[0] = add_82692 == 32'h0000_0000 ? add_82795 : array_index_82789[0];
  assign array_update_82797[1] = add_82692 == 32'h0000_0001 ? add_82795 : array_index_82789[1];
  assign array_update_82797[2] = add_82692 == 32'h0000_0002 ? add_82795 : array_index_82789[2];
  assign array_update_82797[3] = add_82692 == 32'h0000_0003 ? add_82795 : array_index_82789[3];
  assign array_update_82797[4] = add_82692 == 32'h0000_0004 ? add_82795 : array_index_82789[4];
  assign array_update_82797[5] = add_82692 == 32'h0000_0005 ? add_82795 : array_index_82789[5];
  assign array_update_82797[6] = add_82692 == 32'h0000_0006 ? add_82795 : array_index_82789[6];
  assign array_update_82797[7] = add_82692 == 32'h0000_0007 ? add_82795 : array_index_82789[7];
  assign array_update_82797[8] = add_82692 == 32'h0000_0008 ? add_82795 : array_index_82789[8];
  assign array_update_82797[9] = add_82692 == 32'h0000_0009 ? add_82795 : array_index_82789[9];
  assign add_82798 = add_82785 + 32'h0000_0001;
  assign array_update_82799[0] = add_81474 == 32'h0000_0000 ? array_update_82797 : array_update_82786[0];
  assign array_update_82799[1] = add_81474 == 32'h0000_0001 ? array_update_82797 : array_update_82786[1];
  assign array_update_82799[2] = add_81474 == 32'h0000_0002 ? array_update_82797 : array_update_82786[2];
  assign array_update_82799[3] = add_81474 == 32'h0000_0003 ? array_update_82797 : array_update_82786[3];
  assign array_update_82799[4] = add_81474 == 32'h0000_0004 ? array_update_82797 : array_update_82786[4];
  assign array_update_82799[5] = add_81474 == 32'h0000_0005 ? array_update_82797 : array_update_82786[5];
  assign array_update_82799[6] = add_81474 == 32'h0000_0006 ? array_update_82797 : array_update_82786[6];
  assign array_update_82799[7] = add_81474 == 32'h0000_0007 ? array_update_82797 : array_update_82786[7];
  assign array_update_82799[8] = add_81474 == 32'h0000_0008 ? array_update_82797 : array_update_82786[8];
  assign array_update_82799[9] = add_81474 == 32'h0000_0009 ? array_update_82797 : array_update_82786[9];
  assign array_index_82801 = array_update_72021[add_82798 > 32'h0000_0009 ? 4'h9 : add_82798[3:0]];
  assign array_index_82802 = array_update_82799[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_82806 = smul32b_32b_x_32b(array_index_81481[add_82798 > 32'h0000_0009 ? 4'h9 : add_82798[3:0]], array_index_82801[add_82692 > 32'h0000_0009 ? 4'h9 : add_82692[3:0]]);
  assign add_82808 = array_index_82802[add_82692 > 32'h0000_0009 ? 4'h9 : add_82692[3:0]] + smul_82806;
  assign array_update_82810[0] = add_82692 == 32'h0000_0000 ? add_82808 : array_index_82802[0];
  assign array_update_82810[1] = add_82692 == 32'h0000_0001 ? add_82808 : array_index_82802[1];
  assign array_update_82810[2] = add_82692 == 32'h0000_0002 ? add_82808 : array_index_82802[2];
  assign array_update_82810[3] = add_82692 == 32'h0000_0003 ? add_82808 : array_index_82802[3];
  assign array_update_82810[4] = add_82692 == 32'h0000_0004 ? add_82808 : array_index_82802[4];
  assign array_update_82810[5] = add_82692 == 32'h0000_0005 ? add_82808 : array_index_82802[5];
  assign array_update_82810[6] = add_82692 == 32'h0000_0006 ? add_82808 : array_index_82802[6];
  assign array_update_82810[7] = add_82692 == 32'h0000_0007 ? add_82808 : array_index_82802[7];
  assign array_update_82810[8] = add_82692 == 32'h0000_0008 ? add_82808 : array_index_82802[8];
  assign array_update_82810[9] = add_82692 == 32'h0000_0009 ? add_82808 : array_index_82802[9];
  assign add_82811 = add_82798 + 32'h0000_0001;
  assign array_update_82812[0] = add_81474 == 32'h0000_0000 ? array_update_82810 : array_update_82799[0];
  assign array_update_82812[1] = add_81474 == 32'h0000_0001 ? array_update_82810 : array_update_82799[1];
  assign array_update_82812[2] = add_81474 == 32'h0000_0002 ? array_update_82810 : array_update_82799[2];
  assign array_update_82812[3] = add_81474 == 32'h0000_0003 ? array_update_82810 : array_update_82799[3];
  assign array_update_82812[4] = add_81474 == 32'h0000_0004 ? array_update_82810 : array_update_82799[4];
  assign array_update_82812[5] = add_81474 == 32'h0000_0005 ? array_update_82810 : array_update_82799[5];
  assign array_update_82812[6] = add_81474 == 32'h0000_0006 ? array_update_82810 : array_update_82799[6];
  assign array_update_82812[7] = add_81474 == 32'h0000_0007 ? array_update_82810 : array_update_82799[7];
  assign array_update_82812[8] = add_81474 == 32'h0000_0008 ? array_update_82810 : array_update_82799[8];
  assign array_update_82812[9] = add_81474 == 32'h0000_0009 ? array_update_82810 : array_update_82799[9];
  assign array_index_82814 = array_update_72021[add_82811 > 32'h0000_0009 ? 4'h9 : add_82811[3:0]];
  assign array_index_82815 = array_update_82812[add_81474 > 32'h0000_0009 ? 4'h9 : add_81474[3:0]];
  assign smul_82819 = smul32b_32b_x_32b(array_index_81481[add_82811 > 32'h0000_0009 ? 4'h9 : add_82811[3:0]], array_index_82814[add_82692 > 32'h0000_0009 ? 4'h9 : add_82692[3:0]]);
  assign add_82821 = array_index_82815[add_82692 > 32'h0000_0009 ? 4'h9 : add_82692[3:0]] + smul_82819;
  assign array_update_82822[0] = add_82692 == 32'h0000_0000 ? add_82821 : array_index_82815[0];
  assign array_update_82822[1] = add_82692 == 32'h0000_0001 ? add_82821 : array_index_82815[1];
  assign array_update_82822[2] = add_82692 == 32'h0000_0002 ? add_82821 : array_index_82815[2];
  assign array_update_82822[3] = add_82692 == 32'h0000_0003 ? add_82821 : array_index_82815[3];
  assign array_update_82822[4] = add_82692 == 32'h0000_0004 ? add_82821 : array_index_82815[4];
  assign array_update_82822[5] = add_82692 == 32'h0000_0005 ? add_82821 : array_index_82815[5];
  assign array_update_82822[6] = add_82692 == 32'h0000_0006 ? add_82821 : array_index_82815[6];
  assign array_update_82822[7] = add_82692 == 32'h0000_0007 ? add_82821 : array_index_82815[7];
  assign array_update_82822[8] = add_82692 == 32'h0000_0008 ? add_82821 : array_index_82815[8];
  assign array_update_82822[9] = add_82692 == 32'h0000_0009 ? add_82821 : array_index_82815[9];
  assign array_update_82824[0] = add_81474 == 32'h0000_0000 ? array_update_82822 : array_update_82812[0];
  assign array_update_82824[1] = add_81474 == 32'h0000_0001 ? array_update_82822 : array_update_82812[1];
  assign array_update_82824[2] = add_81474 == 32'h0000_0002 ? array_update_82822 : array_update_82812[2];
  assign array_update_82824[3] = add_81474 == 32'h0000_0003 ? array_update_82822 : array_update_82812[3];
  assign array_update_82824[4] = add_81474 == 32'h0000_0004 ? array_update_82822 : array_update_82812[4];
  assign array_update_82824[5] = add_81474 == 32'h0000_0005 ? array_update_82822 : array_update_82812[5];
  assign array_update_82824[6] = add_81474 == 32'h0000_0006 ? array_update_82822 : array_update_82812[6];
  assign array_update_82824[7] = add_81474 == 32'h0000_0007 ? array_update_82822 : array_update_82812[7];
  assign array_update_82824[8] = add_81474 == 32'h0000_0008 ? array_update_82822 : array_update_82812[8];
  assign array_update_82824[9] = add_81474 == 32'h0000_0009 ? array_update_82822 : array_update_82812[9];
  assign add_82825 = add_81474 + 32'h0000_0001;
  assign array_index_82826 = array_update_82824[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign literal_82828 = 32'h0000_0000;
  assign array_update_82829[0] = literal_82828 == 32'h0000_0000 ? 32'h0000_0000 : array_index_82826[0];
  assign array_update_82829[1] = literal_82828 == 32'h0000_0001 ? 32'h0000_0000 : array_index_82826[1];
  assign array_update_82829[2] = literal_82828 == 32'h0000_0002 ? 32'h0000_0000 : array_index_82826[2];
  assign array_update_82829[3] = literal_82828 == 32'h0000_0003 ? 32'h0000_0000 : array_index_82826[3];
  assign array_update_82829[4] = literal_82828 == 32'h0000_0004 ? 32'h0000_0000 : array_index_82826[4];
  assign array_update_82829[5] = literal_82828 == 32'h0000_0005 ? 32'h0000_0000 : array_index_82826[5];
  assign array_update_82829[6] = literal_82828 == 32'h0000_0006 ? 32'h0000_0000 : array_index_82826[6];
  assign array_update_82829[7] = literal_82828 == 32'h0000_0007 ? 32'h0000_0000 : array_index_82826[7];
  assign array_update_82829[8] = literal_82828 == 32'h0000_0008 ? 32'h0000_0000 : array_index_82826[8];
  assign array_update_82829[9] = literal_82828 == 32'h0000_0009 ? 32'h0000_0000 : array_index_82826[9];
  assign literal_82830 = 32'h0000_0000;
  assign array_update_82831[0] = add_82825 == 32'h0000_0000 ? array_update_82829 : array_update_82824[0];
  assign array_update_82831[1] = add_82825 == 32'h0000_0001 ? array_update_82829 : array_update_82824[1];
  assign array_update_82831[2] = add_82825 == 32'h0000_0002 ? array_update_82829 : array_update_82824[2];
  assign array_update_82831[3] = add_82825 == 32'h0000_0003 ? array_update_82829 : array_update_82824[3];
  assign array_update_82831[4] = add_82825 == 32'h0000_0004 ? array_update_82829 : array_update_82824[4];
  assign array_update_82831[5] = add_82825 == 32'h0000_0005 ? array_update_82829 : array_update_82824[5];
  assign array_update_82831[6] = add_82825 == 32'h0000_0006 ? array_update_82829 : array_update_82824[6];
  assign array_update_82831[7] = add_82825 == 32'h0000_0007 ? array_update_82829 : array_update_82824[7];
  assign array_update_82831[8] = add_82825 == 32'h0000_0008 ? array_update_82829 : array_update_82824[8];
  assign array_update_82831[9] = add_82825 == 32'h0000_0009 ? array_update_82829 : array_update_82824[9];
  assign array_index_82832 = array_update_72020[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign array_index_82833 = array_update_72021[literal_82830 > 32'h0000_0009 ? 4'h9 : literal_82830[3:0]];
  assign array_index_82834 = array_update_82831[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_82838 = smul32b_32b_x_32b(array_index_82832[literal_82830 > 32'h0000_0009 ? 4'h9 : literal_82830[3:0]], array_index_82833[literal_82828 > 32'h0000_0009 ? 4'h9 : literal_82828[3:0]]);
  assign add_82840 = array_index_82834[literal_82828 > 32'h0000_0009 ? 4'h9 : literal_82828[3:0]] + smul_82838;
  assign array_update_82842[0] = literal_82828 == 32'h0000_0000 ? add_82840 : array_index_82834[0];
  assign array_update_82842[1] = literal_82828 == 32'h0000_0001 ? add_82840 : array_index_82834[1];
  assign array_update_82842[2] = literal_82828 == 32'h0000_0002 ? add_82840 : array_index_82834[2];
  assign array_update_82842[3] = literal_82828 == 32'h0000_0003 ? add_82840 : array_index_82834[3];
  assign array_update_82842[4] = literal_82828 == 32'h0000_0004 ? add_82840 : array_index_82834[4];
  assign array_update_82842[5] = literal_82828 == 32'h0000_0005 ? add_82840 : array_index_82834[5];
  assign array_update_82842[6] = literal_82828 == 32'h0000_0006 ? add_82840 : array_index_82834[6];
  assign array_update_82842[7] = literal_82828 == 32'h0000_0007 ? add_82840 : array_index_82834[7];
  assign array_update_82842[8] = literal_82828 == 32'h0000_0008 ? add_82840 : array_index_82834[8];
  assign array_update_82842[9] = literal_82828 == 32'h0000_0009 ? add_82840 : array_index_82834[9];
  assign add_82843 = literal_82830 + 32'h0000_0001;
  assign array_update_82844[0] = add_82825 == 32'h0000_0000 ? array_update_82842 : array_update_82831[0];
  assign array_update_82844[1] = add_82825 == 32'h0000_0001 ? array_update_82842 : array_update_82831[1];
  assign array_update_82844[2] = add_82825 == 32'h0000_0002 ? array_update_82842 : array_update_82831[2];
  assign array_update_82844[3] = add_82825 == 32'h0000_0003 ? array_update_82842 : array_update_82831[3];
  assign array_update_82844[4] = add_82825 == 32'h0000_0004 ? array_update_82842 : array_update_82831[4];
  assign array_update_82844[5] = add_82825 == 32'h0000_0005 ? array_update_82842 : array_update_82831[5];
  assign array_update_82844[6] = add_82825 == 32'h0000_0006 ? array_update_82842 : array_update_82831[6];
  assign array_update_82844[7] = add_82825 == 32'h0000_0007 ? array_update_82842 : array_update_82831[7];
  assign array_update_82844[8] = add_82825 == 32'h0000_0008 ? array_update_82842 : array_update_82831[8];
  assign array_update_82844[9] = add_82825 == 32'h0000_0009 ? array_update_82842 : array_update_82831[9];
  assign array_index_82846 = array_update_72021[add_82843 > 32'h0000_0009 ? 4'h9 : add_82843[3:0]];
  assign array_index_82847 = array_update_82844[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_82851 = smul32b_32b_x_32b(array_index_82832[add_82843 > 32'h0000_0009 ? 4'h9 : add_82843[3:0]], array_index_82846[literal_82828 > 32'h0000_0009 ? 4'h9 : literal_82828[3:0]]);
  assign add_82853 = array_index_82847[literal_82828 > 32'h0000_0009 ? 4'h9 : literal_82828[3:0]] + smul_82851;
  assign array_update_82855[0] = literal_82828 == 32'h0000_0000 ? add_82853 : array_index_82847[0];
  assign array_update_82855[1] = literal_82828 == 32'h0000_0001 ? add_82853 : array_index_82847[1];
  assign array_update_82855[2] = literal_82828 == 32'h0000_0002 ? add_82853 : array_index_82847[2];
  assign array_update_82855[3] = literal_82828 == 32'h0000_0003 ? add_82853 : array_index_82847[3];
  assign array_update_82855[4] = literal_82828 == 32'h0000_0004 ? add_82853 : array_index_82847[4];
  assign array_update_82855[5] = literal_82828 == 32'h0000_0005 ? add_82853 : array_index_82847[5];
  assign array_update_82855[6] = literal_82828 == 32'h0000_0006 ? add_82853 : array_index_82847[6];
  assign array_update_82855[7] = literal_82828 == 32'h0000_0007 ? add_82853 : array_index_82847[7];
  assign array_update_82855[8] = literal_82828 == 32'h0000_0008 ? add_82853 : array_index_82847[8];
  assign array_update_82855[9] = literal_82828 == 32'h0000_0009 ? add_82853 : array_index_82847[9];
  assign add_82856 = add_82843 + 32'h0000_0001;
  assign array_update_82857[0] = add_82825 == 32'h0000_0000 ? array_update_82855 : array_update_82844[0];
  assign array_update_82857[1] = add_82825 == 32'h0000_0001 ? array_update_82855 : array_update_82844[1];
  assign array_update_82857[2] = add_82825 == 32'h0000_0002 ? array_update_82855 : array_update_82844[2];
  assign array_update_82857[3] = add_82825 == 32'h0000_0003 ? array_update_82855 : array_update_82844[3];
  assign array_update_82857[4] = add_82825 == 32'h0000_0004 ? array_update_82855 : array_update_82844[4];
  assign array_update_82857[5] = add_82825 == 32'h0000_0005 ? array_update_82855 : array_update_82844[5];
  assign array_update_82857[6] = add_82825 == 32'h0000_0006 ? array_update_82855 : array_update_82844[6];
  assign array_update_82857[7] = add_82825 == 32'h0000_0007 ? array_update_82855 : array_update_82844[7];
  assign array_update_82857[8] = add_82825 == 32'h0000_0008 ? array_update_82855 : array_update_82844[8];
  assign array_update_82857[9] = add_82825 == 32'h0000_0009 ? array_update_82855 : array_update_82844[9];
  assign array_index_82859 = array_update_72021[add_82856 > 32'h0000_0009 ? 4'h9 : add_82856[3:0]];
  assign array_index_82860 = array_update_82857[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_82864 = smul32b_32b_x_32b(array_index_82832[add_82856 > 32'h0000_0009 ? 4'h9 : add_82856[3:0]], array_index_82859[literal_82828 > 32'h0000_0009 ? 4'h9 : literal_82828[3:0]]);
  assign add_82866 = array_index_82860[literal_82828 > 32'h0000_0009 ? 4'h9 : literal_82828[3:0]] + smul_82864;
  assign array_update_82868[0] = literal_82828 == 32'h0000_0000 ? add_82866 : array_index_82860[0];
  assign array_update_82868[1] = literal_82828 == 32'h0000_0001 ? add_82866 : array_index_82860[1];
  assign array_update_82868[2] = literal_82828 == 32'h0000_0002 ? add_82866 : array_index_82860[2];
  assign array_update_82868[3] = literal_82828 == 32'h0000_0003 ? add_82866 : array_index_82860[3];
  assign array_update_82868[4] = literal_82828 == 32'h0000_0004 ? add_82866 : array_index_82860[4];
  assign array_update_82868[5] = literal_82828 == 32'h0000_0005 ? add_82866 : array_index_82860[5];
  assign array_update_82868[6] = literal_82828 == 32'h0000_0006 ? add_82866 : array_index_82860[6];
  assign array_update_82868[7] = literal_82828 == 32'h0000_0007 ? add_82866 : array_index_82860[7];
  assign array_update_82868[8] = literal_82828 == 32'h0000_0008 ? add_82866 : array_index_82860[8];
  assign array_update_82868[9] = literal_82828 == 32'h0000_0009 ? add_82866 : array_index_82860[9];
  assign add_82869 = add_82856 + 32'h0000_0001;
  assign array_update_82870[0] = add_82825 == 32'h0000_0000 ? array_update_82868 : array_update_82857[0];
  assign array_update_82870[1] = add_82825 == 32'h0000_0001 ? array_update_82868 : array_update_82857[1];
  assign array_update_82870[2] = add_82825 == 32'h0000_0002 ? array_update_82868 : array_update_82857[2];
  assign array_update_82870[3] = add_82825 == 32'h0000_0003 ? array_update_82868 : array_update_82857[3];
  assign array_update_82870[4] = add_82825 == 32'h0000_0004 ? array_update_82868 : array_update_82857[4];
  assign array_update_82870[5] = add_82825 == 32'h0000_0005 ? array_update_82868 : array_update_82857[5];
  assign array_update_82870[6] = add_82825 == 32'h0000_0006 ? array_update_82868 : array_update_82857[6];
  assign array_update_82870[7] = add_82825 == 32'h0000_0007 ? array_update_82868 : array_update_82857[7];
  assign array_update_82870[8] = add_82825 == 32'h0000_0008 ? array_update_82868 : array_update_82857[8];
  assign array_update_82870[9] = add_82825 == 32'h0000_0009 ? array_update_82868 : array_update_82857[9];
  assign array_index_82872 = array_update_72021[add_82869 > 32'h0000_0009 ? 4'h9 : add_82869[3:0]];
  assign array_index_82873 = array_update_82870[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_82877 = smul32b_32b_x_32b(array_index_82832[add_82869 > 32'h0000_0009 ? 4'h9 : add_82869[3:0]], array_index_82872[literal_82828 > 32'h0000_0009 ? 4'h9 : literal_82828[3:0]]);
  assign add_82879 = array_index_82873[literal_82828 > 32'h0000_0009 ? 4'h9 : literal_82828[3:0]] + smul_82877;
  assign array_update_82881[0] = literal_82828 == 32'h0000_0000 ? add_82879 : array_index_82873[0];
  assign array_update_82881[1] = literal_82828 == 32'h0000_0001 ? add_82879 : array_index_82873[1];
  assign array_update_82881[2] = literal_82828 == 32'h0000_0002 ? add_82879 : array_index_82873[2];
  assign array_update_82881[3] = literal_82828 == 32'h0000_0003 ? add_82879 : array_index_82873[3];
  assign array_update_82881[4] = literal_82828 == 32'h0000_0004 ? add_82879 : array_index_82873[4];
  assign array_update_82881[5] = literal_82828 == 32'h0000_0005 ? add_82879 : array_index_82873[5];
  assign array_update_82881[6] = literal_82828 == 32'h0000_0006 ? add_82879 : array_index_82873[6];
  assign array_update_82881[7] = literal_82828 == 32'h0000_0007 ? add_82879 : array_index_82873[7];
  assign array_update_82881[8] = literal_82828 == 32'h0000_0008 ? add_82879 : array_index_82873[8];
  assign array_update_82881[9] = literal_82828 == 32'h0000_0009 ? add_82879 : array_index_82873[9];
  assign add_82882 = add_82869 + 32'h0000_0001;
  assign array_update_82883[0] = add_82825 == 32'h0000_0000 ? array_update_82881 : array_update_82870[0];
  assign array_update_82883[1] = add_82825 == 32'h0000_0001 ? array_update_82881 : array_update_82870[1];
  assign array_update_82883[2] = add_82825 == 32'h0000_0002 ? array_update_82881 : array_update_82870[2];
  assign array_update_82883[3] = add_82825 == 32'h0000_0003 ? array_update_82881 : array_update_82870[3];
  assign array_update_82883[4] = add_82825 == 32'h0000_0004 ? array_update_82881 : array_update_82870[4];
  assign array_update_82883[5] = add_82825 == 32'h0000_0005 ? array_update_82881 : array_update_82870[5];
  assign array_update_82883[6] = add_82825 == 32'h0000_0006 ? array_update_82881 : array_update_82870[6];
  assign array_update_82883[7] = add_82825 == 32'h0000_0007 ? array_update_82881 : array_update_82870[7];
  assign array_update_82883[8] = add_82825 == 32'h0000_0008 ? array_update_82881 : array_update_82870[8];
  assign array_update_82883[9] = add_82825 == 32'h0000_0009 ? array_update_82881 : array_update_82870[9];
  assign array_index_82885 = array_update_72021[add_82882 > 32'h0000_0009 ? 4'h9 : add_82882[3:0]];
  assign array_index_82886 = array_update_82883[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_82890 = smul32b_32b_x_32b(array_index_82832[add_82882 > 32'h0000_0009 ? 4'h9 : add_82882[3:0]], array_index_82885[literal_82828 > 32'h0000_0009 ? 4'h9 : literal_82828[3:0]]);
  assign add_82892 = array_index_82886[literal_82828 > 32'h0000_0009 ? 4'h9 : literal_82828[3:0]] + smul_82890;
  assign array_update_82894[0] = literal_82828 == 32'h0000_0000 ? add_82892 : array_index_82886[0];
  assign array_update_82894[1] = literal_82828 == 32'h0000_0001 ? add_82892 : array_index_82886[1];
  assign array_update_82894[2] = literal_82828 == 32'h0000_0002 ? add_82892 : array_index_82886[2];
  assign array_update_82894[3] = literal_82828 == 32'h0000_0003 ? add_82892 : array_index_82886[3];
  assign array_update_82894[4] = literal_82828 == 32'h0000_0004 ? add_82892 : array_index_82886[4];
  assign array_update_82894[5] = literal_82828 == 32'h0000_0005 ? add_82892 : array_index_82886[5];
  assign array_update_82894[6] = literal_82828 == 32'h0000_0006 ? add_82892 : array_index_82886[6];
  assign array_update_82894[7] = literal_82828 == 32'h0000_0007 ? add_82892 : array_index_82886[7];
  assign array_update_82894[8] = literal_82828 == 32'h0000_0008 ? add_82892 : array_index_82886[8];
  assign array_update_82894[9] = literal_82828 == 32'h0000_0009 ? add_82892 : array_index_82886[9];
  assign add_82895 = add_82882 + 32'h0000_0001;
  assign array_update_82896[0] = add_82825 == 32'h0000_0000 ? array_update_82894 : array_update_82883[0];
  assign array_update_82896[1] = add_82825 == 32'h0000_0001 ? array_update_82894 : array_update_82883[1];
  assign array_update_82896[2] = add_82825 == 32'h0000_0002 ? array_update_82894 : array_update_82883[2];
  assign array_update_82896[3] = add_82825 == 32'h0000_0003 ? array_update_82894 : array_update_82883[3];
  assign array_update_82896[4] = add_82825 == 32'h0000_0004 ? array_update_82894 : array_update_82883[4];
  assign array_update_82896[5] = add_82825 == 32'h0000_0005 ? array_update_82894 : array_update_82883[5];
  assign array_update_82896[6] = add_82825 == 32'h0000_0006 ? array_update_82894 : array_update_82883[6];
  assign array_update_82896[7] = add_82825 == 32'h0000_0007 ? array_update_82894 : array_update_82883[7];
  assign array_update_82896[8] = add_82825 == 32'h0000_0008 ? array_update_82894 : array_update_82883[8];
  assign array_update_82896[9] = add_82825 == 32'h0000_0009 ? array_update_82894 : array_update_82883[9];
  assign array_index_82898 = array_update_72021[add_82895 > 32'h0000_0009 ? 4'h9 : add_82895[3:0]];
  assign array_index_82899 = array_update_82896[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_82903 = smul32b_32b_x_32b(array_index_82832[add_82895 > 32'h0000_0009 ? 4'h9 : add_82895[3:0]], array_index_82898[literal_82828 > 32'h0000_0009 ? 4'h9 : literal_82828[3:0]]);
  assign add_82905 = array_index_82899[literal_82828 > 32'h0000_0009 ? 4'h9 : literal_82828[3:0]] + smul_82903;
  assign array_update_82907[0] = literal_82828 == 32'h0000_0000 ? add_82905 : array_index_82899[0];
  assign array_update_82907[1] = literal_82828 == 32'h0000_0001 ? add_82905 : array_index_82899[1];
  assign array_update_82907[2] = literal_82828 == 32'h0000_0002 ? add_82905 : array_index_82899[2];
  assign array_update_82907[3] = literal_82828 == 32'h0000_0003 ? add_82905 : array_index_82899[3];
  assign array_update_82907[4] = literal_82828 == 32'h0000_0004 ? add_82905 : array_index_82899[4];
  assign array_update_82907[5] = literal_82828 == 32'h0000_0005 ? add_82905 : array_index_82899[5];
  assign array_update_82907[6] = literal_82828 == 32'h0000_0006 ? add_82905 : array_index_82899[6];
  assign array_update_82907[7] = literal_82828 == 32'h0000_0007 ? add_82905 : array_index_82899[7];
  assign array_update_82907[8] = literal_82828 == 32'h0000_0008 ? add_82905 : array_index_82899[8];
  assign array_update_82907[9] = literal_82828 == 32'h0000_0009 ? add_82905 : array_index_82899[9];
  assign add_82908 = add_82895 + 32'h0000_0001;
  assign array_update_82909[0] = add_82825 == 32'h0000_0000 ? array_update_82907 : array_update_82896[0];
  assign array_update_82909[1] = add_82825 == 32'h0000_0001 ? array_update_82907 : array_update_82896[1];
  assign array_update_82909[2] = add_82825 == 32'h0000_0002 ? array_update_82907 : array_update_82896[2];
  assign array_update_82909[3] = add_82825 == 32'h0000_0003 ? array_update_82907 : array_update_82896[3];
  assign array_update_82909[4] = add_82825 == 32'h0000_0004 ? array_update_82907 : array_update_82896[4];
  assign array_update_82909[5] = add_82825 == 32'h0000_0005 ? array_update_82907 : array_update_82896[5];
  assign array_update_82909[6] = add_82825 == 32'h0000_0006 ? array_update_82907 : array_update_82896[6];
  assign array_update_82909[7] = add_82825 == 32'h0000_0007 ? array_update_82907 : array_update_82896[7];
  assign array_update_82909[8] = add_82825 == 32'h0000_0008 ? array_update_82907 : array_update_82896[8];
  assign array_update_82909[9] = add_82825 == 32'h0000_0009 ? array_update_82907 : array_update_82896[9];
  assign array_index_82911 = array_update_72021[add_82908 > 32'h0000_0009 ? 4'h9 : add_82908[3:0]];
  assign array_index_82912 = array_update_82909[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_82916 = smul32b_32b_x_32b(array_index_82832[add_82908 > 32'h0000_0009 ? 4'h9 : add_82908[3:0]], array_index_82911[literal_82828 > 32'h0000_0009 ? 4'h9 : literal_82828[3:0]]);
  assign add_82918 = array_index_82912[literal_82828 > 32'h0000_0009 ? 4'h9 : literal_82828[3:0]] + smul_82916;
  assign array_update_82920[0] = literal_82828 == 32'h0000_0000 ? add_82918 : array_index_82912[0];
  assign array_update_82920[1] = literal_82828 == 32'h0000_0001 ? add_82918 : array_index_82912[1];
  assign array_update_82920[2] = literal_82828 == 32'h0000_0002 ? add_82918 : array_index_82912[2];
  assign array_update_82920[3] = literal_82828 == 32'h0000_0003 ? add_82918 : array_index_82912[3];
  assign array_update_82920[4] = literal_82828 == 32'h0000_0004 ? add_82918 : array_index_82912[4];
  assign array_update_82920[5] = literal_82828 == 32'h0000_0005 ? add_82918 : array_index_82912[5];
  assign array_update_82920[6] = literal_82828 == 32'h0000_0006 ? add_82918 : array_index_82912[6];
  assign array_update_82920[7] = literal_82828 == 32'h0000_0007 ? add_82918 : array_index_82912[7];
  assign array_update_82920[8] = literal_82828 == 32'h0000_0008 ? add_82918 : array_index_82912[8];
  assign array_update_82920[9] = literal_82828 == 32'h0000_0009 ? add_82918 : array_index_82912[9];
  assign add_82921 = add_82908 + 32'h0000_0001;
  assign array_update_82922[0] = add_82825 == 32'h0000_0000 ? array_update_82920 : array_update_82909[0];
  assign array_update_82922[1] = add_82825 == 32'h0000_0001 ? array_update_82920 : array_update_82909[1];
  assign array_update_82922[2] = add_82825 == 32'h0000_0002 ? array_update_82920 : array_update_82909[2];
  assign array_update_82922[3] = add_82825 == 32'h0000_0003 ? array_update_82920 : array_update_82909[3];
  assign array_update_82922[4] = add_82825 == 32'h0000_0004 ? array_update_82920 : array_update_82909[4];
  assign array_update_82922[5] = add_82825 == 32'h0000_0005 ? array_update_82920 : array_update_82909[5];
  assign array_update_82922[6] = add_82825 == 32'h0000_0006 ? array_update_82920 : array_update_82909[6];
  assign array_update_82922[7] = add_82825 == 32'h0000_0007 ? array_update_82920 : array_update_82909[7];
  assign array_update_82922[8] = add_82825 == 32'h0000_0008 ? array_update_82920 : array_update_82909[8];
  assign array_update_82922[9] = add_82825 == 32'h0000_0009 ? array_update_82920 : array_update_82909[9];
  assign array_index_82924 = array_update_72021[add_82921 > 32'h0000_0009 ? 4'h9 : add_82921[3:0]];
  assign array_index_82925 = array_update_82922[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_82929 = smul32b_32b_x_32b(array_index_82832[add_82921 > 32'h0000_0009 ? 4'h9 : add_82921[3:0]], array_index_82924[literal_82828 > 32'h0000_0009 ? 4'h9 : literal_82828[3:0]]);
  assign add_82931 = array_index_82925[literal_82828 > 32'h0000_0009 ? 4'h9 : literal_82828[3:0]] + smul_82929;
  assign array_update_82933[0] = literal_82828 == 32'h0000_0000 ? add_82931 : array_index_82925[0];
  assign array_update_82933[1] = literal_82828 == 32'h0000_0001 ? add_82931 : array_index_82925[1];
  assign array_update_82933[2] = literal_82828 == 32'h0000_0002 ? add_82931 : array_index_82925[2];
  assign array_update_82933[3] = literal_82828 == 32'h0000_0003 ? add_82931 : array_index_82925[3];
  assign array_update_82933[4] = literal_82828 == 32'h0000_0004 ? add_82931 : array_index_82925[4];
  assign array_update_82933[5] = literal_82828 == 32'h0000_0005 ? add_82931 : array_index_82925[5];
  assign array_update_82933[6] = literal_82828 == 32'h0000_0006 ? add_82931 : array_index_82925[6];
  assign array_update_82933[7] = literal_82828 == 32'h0000_0007 ? add_82931 : array_index_82925[7];
  assign array_update_82933[8] = literal_82828 == 32'h0000_0008 ? add_82931 : array_index_82925[8];
  assign array_update_82933[9] = literal_82828 == 32'h0000_0009 ? add_82931 : array_index_82925[9];
  assign add_82934 = add_82921 + 32'h0000_0001;
  assign array_update_82935[0] = add_82825 == 32'h0000_0000 ? array_update_82933 : array_update_82922[0];
  assign array_update_82935[1] = add_82825 == 32'h0000_0001 ? array_update_82933 : array_update_82922[1];
  assign array_update_82935[2] = add_82825 == 32'h0000_0002 ? array_update_82933 : array_update_82922[2];
  assign array_update_82935[3] = add_82825 == 32'h0000_0003 ? array_update_82933 : array_update_82922[3];
  assign array_update_82935[4] = add_82825 == 32'h0000_0004 ? array_update_82933 : array_update_82922[4];
  assign array_update_82935[5] = add_82825 == 32'h0000_0005 ? array_update_82933 : array_update_82922[5];
  assign array_update_82935[6] = add_82825 == 32'h0000_0006 ? array_update_82933 : array_update_82922[6];
  assign array_update_82935[7] = add_82825 == 32'h0000_0007 ? array_update_82933 : array_update_82922[7];
  assign array_update_82935[8] = add_82825 == 32'h0000_0008 ? array_update_82933 : array_update_82922[8];
  assign array_update_82935[9] = add_82825 == 32'h0000_0009 ? array_update_82933 : array_update_82922[9];
  assign array_index_82937 = array_update_72021[add_82934 > 32'h0000_0009 ? 4'h9 : add_82934[3:0]];
  assign array_index_82938 = array_update_82935[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_82942 = smul32b_32b_x_32b(array_index_82832[add_82934 > 32'h0000_0009 ? 4'h9 : add_82934[3:0]], array_index_82937[literal_82828 > 32'h0000_0009 ? 4'h9 : literal_82828[3:0]]);
  assign add_82944 = array_index_82938[literal_82828 > 32'h0000_0009 ? 4'h9 : literal_82828[3:0]] + smul_82942;
  assign array_update_82946[0] = literal_82828 == 32'h0000_0000 ? add_82944 : array_index_82938[0];
  assign array_update_82946[1] = literal_82828 == 32'h0000_0001 ? add_82944 : array_index_82938[1];
  assign array_update_82946[2] = literal_82828 == 32'h0000_0002 ? add_82944 : array_index_82938[2];
  assign array_update_82946[3] = literal_82828 == 32'h0000_0003 ? add_82944 : array_index_82938[3];
  assign array_update_82946[4] = literal_82828 == 32'h0000_0004 ? add_82944 : array_index_82938[4];
  assign array_update_82946[5] = literal_82828 == 32'h0000_0005 ? add_82944 : array_index_82938[5];
  assign array_update_82946[6] = literal_82828 == 32'h0000_0006 ? add_82944 : array_index_82938[6];
  assign array_update_82946[7] = literal_82828 == 32'h0000_0007 ? add_82944 : array_index_82938[7];
  assign array_update_82946[8] = literal_82828 == 32'h0000_0008 ? add_82944 : array_index_82938[8];
  assign array_update_82946[9] = literal_82828 == 32'h0000_0009 ? add_82944 : array_index_82938[9];
  assign add_82947 = add_82934 + 32'h0000_0001;
  assign array_update_82948[0] = add_82825 == 32'h0000_0000 ? array_update_82946 : array_update_82935[0];
  assign array_update_82948[1] = add_82825 == 32'h0000_0001 ? array_update_82946 : array_update_82935[1];
  assign array_update_82948[2] = add_82825 == 32'h0000_0002 ? array_update_82946 : array_update_82935[2];
  assign array_update_82948[3] = add_82825 == 32'h0000_0003 ? array_update_82946 : array_update_82935[3];
  assign array_update_82948[4] = add_82825 == 32'h0000_0004 ? array_update_82946 : array_update_82935[4];
  assign array_update_82948[5] = add_82825 == 32'h0000_0005 ? array_update_82946 : array_update_82935[5];
  assign array_update_82948[6] = add_82825 == 32'h0000_0006 ? array_update_82946 : array_update_82935[6];
  assign array_update_82948[7] = add_82825 == 32'h0000_0007 ? array_update_82946 : array_update_82935[7];
  assign array_update_82948[8] = add_82825 == 32'h0000_0008 ? array_update_82946 : array_update_82935[8];
  assign array_update_82948[9] = add_82825 == 32'h0000_0009 ? array_update_82946 : array_update_82935[9];
  assign array_index_82950 = array_update_72021[add_82947 > 32'h0000_0009 ? 4'h9 : add_82947[3:0]];
  assign array_index_82951 = array_update_82948[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_82955 = smul32b_32b_x_32b(array_index_82832[add_82947 > 32'h0000_0009 ? 4'h9 : add_82947[3:0]], array_index_82950[literal_82828 > 32'h0000_0009 ? 4'h9 : literal_82828[3:0]]);
  assign add_82957 = array_index_82951[literal_82828 > 32'h0000_0009 ? 4'h9 : literal_82828[3:0]] + smul_82955;
  assign array_update_82958[0] = literal_82828 == 32'h0000_0000 ? add_82957 : array_index_82951[0];
  assign array_update_82958[1] = literal_82828 == 32'h0000_0001 ? add_82957 : array_index_82951[1];
  assign array_update_82958[2] = literal_82828 == 32'h0000_0002 ? add_82957 : array_index_82951[2];
  assign array_update_82958[3] = literal_82828 == 32'h0000_0003 ? add_82957 : array_index_82951[3];
  assign array_update_82958[4] = literal_82828 == 32'h0000_0004 ? add_82957 : array_index_82951[4];
  assign array_update_82958[5] = literal_82828 == 32'h0000_0005 ? add_82957 : array_index_82951[5];
  assign array_update_82958[6] = literal_82828 == 32'h0000_0006 ? add_82957 : array_index_82951[6];
  assign array_update_82958[7] = literal_82828 == 32'h0000_0007 ? add_82957 : array_index_82951[7];
  assign array_update_82958[8] = literal_82828 == 32'h0000_0008 ? add_82957 : array_index_82951[8];
  assign array_update_82958[9] = literal_82828 == 32'h0000_0009 ? add_82957 : array_index_82951[9];
  assign array_update_82959[0] = add_82825 == 32'h0000_0000 ? array_update_82958 : array_update_82948[0];
  assign array_update_82959[1] = add_82825 == 32'h0000_0001 ? array_update_82958 : array_update_82948[1];
  assign array_update_82959[2] = add_82825 == 32'h0000_0002 ? array_update_82958 : array_update_82948[2];
  assign array_update_82959[3] = add_82825 == 32'h0000_0003 ? array_update_82958 : array_update_82948[3];
  assign array_update_82959[4] = add_82825 == 32'h0000_0004 ? array_update_82958 : array_update_82948[4];
  assign array_update_82959[5] = add_82825 == 32'h0000_0005 ? array_update_82958 : array_update_82948[5];
  assign array_update_82959[6] = add_82825 == 32'h0000_0006 ? array_update_82958 : array_update_82948[6];
  assign array_update_82959[7] = add_82825 == 32'h0000_0007 ? array_update_82958 : array_update_82948[7];
  assign array_update_82959[8] = add_82825 == 32'h0000_0008 ? array_update_82958 : array_update_82948[8];
  assign array_update_82959[9] = add_82825 == 32'h0000_0009 ? array_update_82958 : array_update_82948[9];
  assign array_index_82961 = array_update_82959[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign add_82963 = literal_82828 + 32'h0000_0001;
  assign array_update_82964[0] = add_82963 == 32'h0000_0000 ? 32'h0000_0000 : array_index_82961[0];
  assign array_update_82964[1] = add_82963 == 32'h0000_0001 ? 32'h0000_0000 : array_index_82961[1];
  assign array_update_82964[2] = add_82963 == 32'h0000_0002 ? 32'h0000_0000 : array_index_82961[2];
  assign array_update_82964[3] = add_82963 == 32'h0000_0003 ? 32'h0000_0000 : array_index_82961[3];
  assign array_update_82964[4] = add_82963 == 32'h0000_0004 ? 32'h0000_0000 : array_index_82961[4];
  assign array_update_82964[5] = add_82963 == 32'h0000_0005 ? 32'h0000_0000 : array_index_82961[5];
  assign array_update_82964[6] = add_82963 == 32'h0000_0006 ? 32'h0000_0000 : array_index_82961[6];
  assign array_update_82964[7] = add_82963 == 32'h0000_0007 ? 32'h0000_0000 : array_index_82961[7];
  assign array_update_82964[8] = add_82963 == 32'h0000_0008 ? 32'h0000_0000 : array_index_82961[8];
  assign array_update_82964[9] = add_82963 == 32'h0000_0009 ? 32'h0000_0000 : array_index_82961[9];
  assign literal_82965 = 32'h0000_0000;
  assign array_update_82966[0] = add_82825 == 32'h0000_0000 ? array_update_82964 : array_update_82959[0];
  assign array_update_82966[1] = add_82825 == 32'h0000_0001 ? array_update_82964 : array_update_82959[1];
  assign array_update_82966[2] = add_82825 == 32'h0000_0002 ? array_update_82964 : array_update_82959[2];
  assign array_update_82966[3] = add_82825 == 32'h0000_0003 ? array_update_82964 : array_update_82959[3];
  assign array_update_82966[4] = add_82825 == 32'h0000_0004 ? array_update_82964 : array_update_82959[4];
  assign array_update_82966[5] = add_82825 == 32'h0000_0005 ? array_update_82964 : array_update_82959[5];
  assign array_update_82966[6] = add_82825 == 32'h0000_0006 ? array_update_82964 : array_update_82959[6];
  assign array_update_82966[7] = add_82825 == 32'h0000_0007 ? array_update_82964 : array_update_82959[7];
  assign array_update_82966[8] = add_82825 == 32'h0000_0008 ? array_update_82964 : array_update_82959[8];
  assign array_update_82966[9] = add_82825 == 32'h0000_0009 ? array_update_82964 : array_update_82959[9];
  assign array_index_82968 = array_update_72021[literal_82965 > 32'h0000_0009 ? 4'h9 : literal_82965[3:0]];
  assign array_index_82969 = array_update_82966[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_82973 = smul32b_32b_x_32b(array_index_82832[literal_82965 > 32'h0000_0009 ? 4'h9 : literal_82965[3:0]], array_index_82968[add_82963 > 32'h0000_0009 ? 4'h9 : add_82963[3:0]]);
  assign add_82975 = array_index_82969[add_82963 > 32'h0000_0009 ? 4'h9 : add_82963[3:0]] + smul_82973;
  assign array_update_82977[0] = add_82963 == 32'h0000_0000 ? add_82975 : array_index_82969[0];
  assign array_update_82977[1] = add_82963 == 32'h0000_0001 ? add_82975 : array_index_82969[1];
  assign array_update_82977[2] = add_82963 == 32'h0000_0002 ? add_82975 : array_index_82969[2];
  assign array_update_82977[3] = add_82963 == 32'h0000_0003 ? add_82975 : array_index_82969[3];
  assign array_update_82977[4] = add_82963 == 32'h0000_0004 ? add_82975 : array_index_82969[4];
  assign array_update_82977[5] = add_82963 == 32'h0000_0005 ? add_82975 : array_index_82969[5];
  assign array_update_82977[6] = add_82963 == 32'h0000_0006 ? add_82975 : array_index_82969[6];
  assign array_update_82977[7] = add_82963 == 32'h0000_0007 ? add_82975 : array_index_82969[7];
  assign array_update_82977[8] = add_82963 == 32'h0000_0008 ? add_82975 : array_index_82969[8];
  assign array_update_82977[9] = add_82963 == 32'h0000_0009 ? add_82975 : array_index_82969[9];
  assign add_82978 = literal_82965 + 32'h0000_0001;
  assign array_update_82979[0] = add_82825 == 32'h0000_0000 ? array_update_82977 : array_update_82966[0];
  assign array_update_82979[1] = add_82825 == 32'h0000_0001 ? array_update_82977 : array_update_82966[1];
  assign array_update_82979[2] = add_82825 == 32'h0000_0002 ? array_update_82977 : array_update_82966[2];
  assign array_update_82979[3] = add_82825 == 32'h0000_0003 ? array_update_82977 : array_update_82966[3];
  assign array_update_82979[4] = add_82825 == 32'h0000_0004 ? array_update_82977 : array_update_82966[4];
  assign array_update_82979[5] = add_82825 == 32'h0000_0005 ? array_update_82977 : array_update_82966[5];
  assign array_update_82979[6] = add_82825 == 32'h0000_0006 ? array_update_82977 : array_update_82966[6];
  assign array_update_82979[7] = add_82825 == 32'h0000_0007 ? array_update_82977 : array_update_82966[7];
  assign array_update_82979[8] = add_82825 == 32'h0000_0008 ? array_update_82977 : array_update_82966[8];
  assign array_update_82979[9] = add_82825 == 32'h0000_0009 ? array_update_82977 : array_update_82966[9];
  assign array_index_82981 = array_update_72021[add_82978 > 32'h0000_0009 ? 4'h9 : add_82978[3:0]];
  assign array_index_82982 = array_update_82979[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_82986 = smul32b_32b_x_32b(array_index_82832[add_82978 > 32'h0000_0009 ? 4'h9 : add_82978[3:0]], array_index_82981[add_82963 > 32'h0000_0009 ? 4'h9 : add_82963[3:0]]);
  assign add_82988 = array_index_82982[add_82963 > 32'h0000_0009 ? 4'h9 : add_82963[3:0]] + smul_82986;
  assign array_update_82990[0] = add_82963 == 32'h0000_0000 ? add_82988 : array_index_82982[0];
  assign array_update_82990[1] = add_82963 == 32'h0000_0001 ? add_82988 : array_index_82982[1];
  assign array_update_82990[2] = add_82963 == 32'h0000_0002 ? add_82988 : array_index_82982[2];
  assign array_update_82990[3] = add_82963 == 32'h0000_0003 ? add_82988 : array_index_82982[3];
  assign array_update_82990[4] = add_82963 == 32'h0000_0004 ? add_82988 : array_index_82982[4];
  assign array_update_82990[5] = add_82963 == 32'h0000_0005 ? add_82988 : array_index_82982[5];
  assign array_update_82990[6] = add_82963 == 32'h0000_0006 ? add_82988 : array_index_82982[6];
  assign array_update_82990[7] = add_82963 == 32'h0000_0007 ? add_82988 : array_index_82982[7];
  assign array_update_82990[8] = add_82963 == 32'h0000_0008 ? add_82988 : array_index_82982[8];
  assign array_update_82990[9] = add_82963 == 32'h0000_0009 ? add_82988 : array_index_82982[9];
  assign add_82991 = add_82978 + 32'h0000_0001;
  assign array_update_82992[0] = add_82825 == 32'h0000_0000 ? array_update_82990 : array_update_82979[0];
  assign array_update_82992[1] = add_82825 == 32'h0000_0001 ? array_update_82990 : array_update_82979[1];
  assign array_update_82992[2] = add_82825 == 32'h0000_0002 ? array_update_82990 : array_update_82979[2];
  assign array_update_82992[3] = add_82825 == 32'h0000_0003 ? array_update_82990 : array_update_82979[3];
  assign array_update_82992[4] = add_82825 == 32'h0000_0004 ? array_update_82990 : array_update_82979[4];
  assign array_update_82992[5] = add_82825 == 32'h0000_0005 ? array_update_82990 : array_update_82979[5];
  assign array_update_82992[6] = add_82825 == 32'h0000_0006 ? array_update_82990 : array_update_82979[6];
  assign array_update_82992[7] = add_82825 == 32'h0000_0007 ? array_update_82990 : array_update_82979[7];
  assign array_update_82992[8] = add_82825 == 32'h0000_0008 ? array_update_82990 : array_update_82979[8];
  assign array_update_82992[9] = add_82825 == 32'h0000_0009 ? array_update_82990 : array_update_82979[9];
  assign array_index_82994 = array_update_72021[add_82991 > 32'h0000_0009 ? 4'h9 : add_82991[3:0]];
  assign array_index_82995 = array_update_82992[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_82999 = smul32b_32b_x_32b(array_index_82832[add_82991 > 32'h0000_0009 ? 4'h9 : add_82991[3:0]], array_index_82994[add_82963 > 32'h0000_0009 ? 4'h9 : add_82963[3:0]]);
  assign add_83001 = array_index_82995[add_82963 > 32'h0000_0009 ? 4'h9 : add_82963[3:0]] + smul_82999;
  assign array_update_83003[0] = add_82963 == 32'h0000_0000 ? add_83001 : array_index_82995[0];
  assign array_update_83003[1] = add_82963 == 32'h0000_0001 ? add_83001 : array_index_82995[1];
  assign array_update_83003[2] = add_82963 == 32'h0000_0002 ? add_83001 : array_index_82995[2];
  assign array_update_83003[3] = add_82963 == 32'h0000_0003 ? add_83001 : array_index_82995[3];
  assign array_update_83003[4] = add_82963 == 32'h0000_0004 ? add_83001 : array_index_82995[4];
  assign array_update_83003[5] = add_82963 == 32'h0000_0005 ? add_83001 : array_index_82995[5];
  assign array_update_83003[6] = add_82963 == 32'h0000_0006 ? add_83001 : array_index_82995[6];
  assign array_update_83003[7] = add_82963 == 32'h0000_0007 ? add_83001 : array_index_82995[7];
  assign array_update_83003[8] = add_82963 == 32'h0000_0008 ? add_83001 : array_index_82995[8];
  assign array_update_83003[9] = add_82963 == 32'h0000_0009 ? add_83001 : array_index_82995[9];
  assign add_83004 = add_82991 + 32'h0000_0001;
  assign array_update_83005[0] = add_82825 == 32'h0000_0000 ? array_update_83003 : array_update_82992[0];
  assign array_update_83005[1] = add_82825 == 32'h0000_0001 ? array_update_83003 : array_update_82992[1];
  assign array_update_83005[2] = add_82825 == 32'h0000_0002 ? array_update_83003 : array_update_82992[2];
  assign array_update_83005[3] = add_82825 == 32'h0000_0003 ? array_update_83003 : array_update_82992[3];
  assign array_update_83005[4] = add_82825 == 32'h0000_0004 ? array_update_83003 : array_update_82992[4];
  assign array_update_83005[5] = add_82825 == 32'h0000_0005 ? array_update_83003 : array_update_82992[5];
  assign array_update_83005[6] = add_82825 == 32'h0000_0006 ? array_update_83003 : array_update_82992[6];
  assign array_update_83005[7] = add_82825 == 32'h0000_0007 ? array_update_83003 : array_update_82992[7];
  assign array_update_83005[8] = add_82825 == 32'h0000_0008 ? array_update_83003 : array_update_82992[8];
  assign array_update_83005[9] = add_82825 == 32'h0000_0009 ? array_update_83003 : array_update_82992[9];
  assign array_index_83007 = array_update_72021[add_83004 > 32'h0000_0009 ? 4'h9 : add_83004[3:0]];
  assign array_index_83008 = array_update_83005[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_83012 = smul32b_32b_x_32b(array_index_82832[add_83004 > 32'h0000_0009 ? 4'h9 : add_83004[3:0]], array_index_83007[add_82963 > 32'h0000_0009 ? 4'h9 : add_82963[3:0]]);
  assign add_83014 = array_index_83008[add_82963 > 32'h0000_0009 ? 4'h9 : add_82963[3:0]] + smul_83012;
  assign array_update_83016[0] = add_82963 == 32'h0000_0000 ? add_83014 : array_index_83008[0];
  assign array_update_83016[1] = add_82963 == 32'h0000_0001 ? add_83014 : array_index_83008[1];
  assign array_update_83016[2] = add_82963 == 32'h0000_0002 ? add_83014 : array_index_83008[2];
  assign array_update_83016[3] = add_82963 == 32'h0000_0003 ? add_83014 : array_index_83008[3];
  assign array_update_83016[4] = add_82963 == 32'h0000_0004 ? add_83014 : array_index_83008[4];
  assign array_update_83016[5] = add_82963 == 32'h0000_0005 ? add_83014 : array_index_83008[5];
  assign array_update_83016[6] = add_82963 == 32'h0000_0006 ? add_83014 : array_index_83008[6];
  assign array_update_83016[7] = add_82963 == 32'h0000_0007 ? add_83014 : array_index_83008[7];
  assign array_update_83016[8] = add_82963 == 32'h0000_0008 ? add_83014 : array_index_83008[8];
  assign array_update_83016[9] = add_82963 == 32'h0000_0009 ? add_83014 : array_index_83008[9];
  assign add_83017 = add_83004 + 32'h0000_0001;
  assign array_update_83018[0] = add_82825 == 32'h0000_0000 ? array_update_83016 : array_update_83005[0];
  assign array_update_83018[1] = add_82825 == 32'h0000_0001 ? array_update_83016 : array_update_83005[1];
  assign array_update_83018[2] = add_82825 == 32'h0000_0002 ? array_update_83016 : array_update_83005[2];
  assign array_update_83018[3] = add_82825 == 32'h0000_0003 ? array_update_83016 : array_update_83005[3];
  assign array_update_83018[4] = add_82825 == 32'h0000_0004 ? array_update_83016 : array_update_83005[4];
  assign array_update_83018[5] = add_82825 == 32'h0000_0005 ? array_update_83016 : array_update_83005[5];
  assign array_update_83018[6] = add_82825 == 32'h0000_0006 ? array_update_83016 : array_update_83005[6];
  assign array_update_83018[7] = add_82825 == 32'h0000_0007 ? array_update_83016 : array_update_83005[7];
  assign array_update_83018[8] = add_82825 == 32'h0000_0008 ? array_update_83016 : array_update_83005[8];
  assign array_update_83018[9] = add_82825 == 32'h0000_0009 ? array_update_83016 : array_update_83005[9];
  assign array_index_83020 = array_update_72021[add_83017 > 32'h0000_0009 ? 4'h9 : add_83017[3:0]];
  assign array_index_83021 = array_update_83018[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_83025 = smul32b_32b_x_32b(array_index_82832[add_83017 > 32'h0000_0009 ? 4'h9 : add_83017[3:0]], array_index_83020[add_82963 > 32'h0000_0009 ? 4'h9 : add_82963[3:0]]);
  assign add_83027 = array_index_83021[add_82963 > 32'h0000_0009 ? 4'h9 : add_82963[3:0]] + smul_83025;
  assign array_update_83029[0] = add_82963 == 32'h0000_0000 ? add_83027 : array_index_83021[0];
  assign array_update_83029[1] = add_82963 == 32'h0000_0001 ? add_83027 : array_index_83021[1];
  assign array_update_83029[2] = add_82963 == 32'h0000_0002 ? add_83027 : array_index_83021[2];
  assign array_update_83029[3] = add_82963 == 32'h0000_0003 ? add_83027 : array_index_83021[3];
  assign array_update_83029[4] = add_82963 == 32'h0000_0004 ? add_83027 : array_index_83021[4];
  assign array_update_83029[5] = add_82963 == 32'h0000_0005 ? add_83027 : array_index_83021[5];
  assign array_update_83029[6] = add_82963 == 32'h0000_0006 ? add_83027 : array_index_83021[6];
  assign array_update_83029[7] = add_82963 == 32'h0000_0007 ? add_83027 : array_index_83021[7];
  assign array_update_83029[8] = add_82963 == 32'h0000_0008 ? add_83027 : array_index_83021[8];
  assign array_update_83029[9] = add_82963 == 32'h0000_0009 ? add_83027 : array_index_83021[9];
  assign add_83030 = add_83017 + 32'h0000_0001;
  assign array_update_83031[0] = add_82825 == 32'h0000_0000 ? array_update_83029 : array_update_83018[0];
  assign array_update_83031[1] = add_82825 == 32'h0000_0001 ? array_update_83029 : array_update_83018[1];
  assign array_update_83031[2] = add_82825 == 32'h0000_0002 ? array_update_83029 : array_update_83018[2];
  assign array_update_83031[3] = add_82825 == 32'h0000_0003 ? array_update_83029 : array_update_83018[3];
  assign array_update_83031[4] = add_82825 == 32'h0000_0004 ? array_update_83029 : array_update_83018[4];
  assign array_update_83031[5] = add_82825 == 32'h0000_0005 ? array_update_83029 : array_update_83018[5];
  assign array_update_83031[6] = add_82825 == 32'h0000_0006 ? array_update_83029 : array_update_83018[6];
  assign array_update_83031[7] = add_82825 == 32'h0000_0007 ? array_update_83029 : array_update_83018[7];
  assign array_update_83031[8] = add_82825 == 32'h0000_0008 ? array_update_83029 : array_update_83018[8];
  assign array_update_83031[9] = add_82825 == 32'h0000_0009 ? array_update_83029 : array_update_83018[9];
  assign array_index_83033 = array_update_72021[add_83030 > 32'h0000_0009 ? 4'h9 : add_83030[3:0]];
  assign array_index_83034 = array_update_83031[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_83038 = smul32b_32b_x_32b(array_index_82832[add_83030 > 32'h0000_0009 ? 4'h9 : add_83030[3:0]], array_index_83033[add_82963 > 32'h0000_0009 ? 4'h9 : add_82963[3:0]]);
  assign add_83040 = array_index_83034[add_82963 > 32'h0000_0009 ? 4'h9 : add_82963[3:0]] + smul_83038;
  assign array_update_83042[0] = add_82963 == 32'h0000_0000 ? add_83040 : array_index_83034[0];
  assign array_update_83042[1] = add_82963 == 32'h0000_0001 ? add_83040 : array_index_83034[1];
  assign array_update_83042[2] = add_82963 == 32'h0000_0002 ? add_83040 : array_index_83034[2];
  assign array_update_83042[3] = add_82963 == 32'h0000_0003 ? add_83040 : array_index_83034[3];
  assign array_update_83042[4] = add_82963 == 32'h0000_0004 ? add_83040 : array_index_83034[4];
  assign array_update_83042[5] = add_82963 == 32'h0000_0005 ? add_83040 : array_index_83034[5];
  assign array_update_83042[6] = add_82963 == 32'h0000_0006 ? add_83040 : array_index_83034[6];
  assign array_update_83042[7] = add_82963 == 32'h0000_0007 ? add_83040 : array_index_83034[7];
  assign array_update_83042[8] = add_82963 == 32'h0000_0008 ? add_83040 : array_index_83034[8];
  assign array_update_83042[9] = add_82963 == 32'h0000_0009 ? add_83040 : array_index_83034[9];
  assign add_83043 = add_83030 + 32'h0000_0001;
  assign array_update_83044[0] = add_82825 == 32'h0000_0000 ? array_update_83042 : array_update_83031[0];
  assign array_update_83044[1] = add_82825 == 32'h0000_0001 ? array_update_83042 : array_update_83031[1];
  assign array_update_83044[2] = add_82825 == 32'h0000_0002 ? array_update_83042 : array_update_83031[2];
  assign array_update_83044[3] = add_82825 == 32'h0000_0003 ? array_update_83042 : array_update_83031[3];
  assign array_update_83044[4] = add_82825 == 32'h0000_0004 ? array_update_83042 : array_update_83031[4];
  assign array_update_83044[5] = add_82825 == 32'h0000_0005 ? array_update_83042 : array_update_83031[5];
  assign array_update_83044[6] = add_82825 == 32'h0000_0006 ? array_update_83042 : array_update_83031[6];
  assign array_update_83044[7] = add_82825 == 32'h0000_0007 ? array_update_83042 : array_update_83031[7];
  assign array_update_83044[8] = add_82825 == 32'h0000_0008 ? array_update_83042 : array_update_83031[8];
  assign array_update_83044[9] = add_82825 == 32'h0000_0009 ? array_update_83042 : array_update_83031[9];
  assign array_index_83046 = array_update_72021[add_83043 > 32'h0000_0009 ? 4'h9 : add_83043[3:0]];
  assign array_index_83047 = array_update_83044[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_83051 = smul32b_32b_x_32b(array_index_82832[add_83043 > 32'h0000_0009 ? 4'h9 : add_83043[3:0]], array_index_83046[add_82963 > 32'h0000_0009 ? 4'h9 : add_82963[3:0]]);
  assign add_83053 = array_index_83047[add_82963 > 32'h0000_0009 ? 4'h9 : add_82963[3:0]] + smul_83051;
  assign array_update_83055[0] = add_82963 == 32'h0000_0000 ? add_83053 : array_index_83047[0];
  assign array_update_83055[1] = add_82963 == 32'h0000_0001 ? add_83053 : array_index_83047[1];
  assign array_update_83055[2] = add_82963 == 32'h0000_0002 ? add_83053 : array_index_83047[2];
  assign array_update_83055[3] = add_82963 == 32'h0000_0003 ? add_83053 : array_index_83047[3];
  assign array_update_83055[4] = add_82963 == 32'h0000_0004 ? add_83053 : array_index_83047[4];
  assign array_update_83055[5] = add_82963 == 32'h0000_0005 ? add_83053 : array_index_83047[5];
  assign array_update_83055[6] = add_82963 == 32'h0000_0006 ? add_83053 : array_index_83047[6];
  assign array_update_83055[7] = add_82963 == 32'h0000_0007 ? add_83053 : array_index_83047[7];
  assign array_update_83055[8] = add_82963 == 32'h0000_0008 ? add_83053 : array_index_83047[8];
  assign array_update_83055[9] = add_82963 == 32'h0000_0009 ? add_83053 : array_index_83047[9];
  assign add_83056 = add_83043 + 32'h0000_0001;
  assign array_update_83057[0] = add_82825 == 32'h0000_0000 ? array_update_83055 : array_update_83044[0];
  assign array_update_83057[1] = add_82825 == 32'h0000_0001 ? array_update_83055 : array_update_83044[1];
  assign array_update_83057[2] = add_82825 == 32'h0000_0002 ? array_update_83055 : array_update_83044[2];
  assign array_update_83057[3] = add_82825 == 32'h0000_0003 ? array_update_83055 : array_update_83044[3];
  assign array_update_83057[4] = add_82825 == 32'h0000_0004 ? array_update_83055 : array_update_83044[4];
  assign array_update_83057[5] = add_82825 == 32'h0000_0005 ? array_update_83055 : array_update_83044[5];
  assign array_update_83057[6] = add_82825 == 32'h0000_0006 ? array_update_83055 : array_update_83044[6];
  assign array_update_83057[7] = add_82825 == 32'h0000_0007 ? array_update_83055 : array_update_83044[7];
  assign array_update_83057[8] = add_82825 == 32'h0000_0008 ? array_update_83055 : array_update_83044[8];
  assign array_update_83057[9] = add_82825 == 32'h0000_0009 ? array_update_83055 : array_update_83044[9];
  assign array_index_83059 = array_update_72021[add_83056 > 32'h0000_0009 ? 4'h9 : add_83056[3:0]];
  assign array_index_83060 = array_update_83057[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_83064 = smul32b_32b_x_32b(array_index_82832[add_83056 > 32'h0000_0009 ? 4'h9 : add_83056[3:0]], array_index_83059[add_82963 > 32'h0000_0009 ? 4'h9 : add_82963[3:0]]);
  assign add_83066 = array_index_83060[add_82963 > 32'h0000_0009 ? 4'h9 : add_82963[3:0]] + smul_83064;
  assign array_update_83068[0] = add_82963 == 32'h0000_0000 ? add_83066 : array_index_83060[0];
  assign array_update_83068[1] = add_82963 == 32'h0000_0001 ? add_83066 : array_index_83060[1];
  assign array_update_83068[2] = add_82963 == 32'h0000_0002 ? add_83066 : array_index_83060[2];
  assign array_update_83068[3] = add_82963 == 32'h0000_0003 ? add_83066 : array_index_83060[3];
  assign array_update_83068[4] = add_82963 == 32'h0000_0004 ? add_83066 : array_index_83060[4];
  assign array_update_83068[5] = add_82963 == 32'h0000_0005 ? add_83066 : array_index_83060[5];
  assign array_update_83068[6] = add_82963 == 32'h0000_0006 ? add_83066 : array_index_83060[6];
  assign array_update_83068[7] = add_82963 == 32'h0000_0007 ? add_83066 : array_index_83060[7];
  assign array_update_83068[8] = add_82963 == 32'h0000_0008 ? add_83066 : array_index_83060[8];
  assign array_update_83068[9] = add_82963 == 32'h0000_0009 ? add_83066 : array_index_83060[9];
  assign add_83069 = add_83056 + 32'h0000_0001;
  assign array_update_83070[0] = add_82825 == 32'h0000_0000 ? array_update_83068 : array_update_83057[0];
  assign array_update_83070[1] = add_82825 == 32'h0000_0001 ? array_update_83068 : array_update_83057[1];
  assign array_update_83070[2] = add_82825 == 32'h0000_0002 ? array_update_83068 : array_update_83057[2];
  assign array_update_83070[3] = add_82825 == 32'h0000_0003 ? array_update_83068 : array_update_83057[3];
  assign array_update_83070[4] = add_82825 == 32'h0000_0004 ? array_update_83068 : array_update_83057[4];
  assign array_update_83070[5] = add_82825 == 32'h0000_0005 ? array_update_83068 : array_update_83057[5];
  assign array_update_83070[6] = add_82825 == 32'h0000_0006 ? array_update_83068 : array_update_83057[6];
  assign array_update_83070[7] = add_82825 == 32'h0000_0007 ? array_update_83068 : array_update_83057[7];
  assign array_update_83070[8] = add_82825 == 32'h0000_0008 ? array_update_83068 : array_update_83057[8];
  assign array_update_83070[9] = add_82825 == 32'h0000_0009 ? array_update_83068 : array_update_83057[9];
  assign array_index_83072 = array_update_72021[add_83069 > 32'h0000_0009 ? 4'h9 : add_83069[3:0]];
  assign array_index_83073 = array_update_83070[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_83077 = smul32b_32b_x_32b(array_index_82832[add_83069 > 32'h0000_0009 ? 4'h9 : add_83069[3:0]], array_index_83072[add_82963 > 32'h0000_0009 ? 4'h9 : add_82963[3:0]]);
  assign add_83079 = array_index_83073[add_82963 > 32'h0000_0009 ? 4'h9 : add_82963[3:0]] + smul_83077;
  assign array_update_83081[0] = add_82963 == 32'h0000_0000 ? add_83079 : array_index_83073[0];
  assign array_update_83081[1] = add_82963 == 32'h0000_0001 ? add_83079 : array_index_83073[1];
  assign array_update_83081[2] = add_82963 == 32'h0000_0002 ? add_83079 : array_index_83073[2];
  assign array_update_83081[3] = add_82963 == 32'h0000_0003 ? add_83079 : array_index_83073[3];
  assign array_update_83081[4] = add_82963 == 32'h0000_0004 ? add_83079 : array_index_83073[4];
  assign array_update_83081[5] = add_82963 == 32'h0000_0005 ? add_83079 : array_index_83073[5];
  assign array_update_83081[6] = add_82963 == 32'h0000_0006 ? add_83079 : array_index_83073[6];
  assign array_update_83081[7] = add_82963 == 32'h0000_0007 ? add_83079 : array_index_83073[7];
  assign array_update_83081[8] = add_82963 == 32'h0000_0008 ? add_83079 : array_index_83073[8];
  assign array_update_83081[9] = add_82963 == 32'h0000_0009 ? add_83079 : array_index_83073[9];
  assign add_83082 = add_83069 + 32'h0000_0001;
  assign array_update_83083[0] = add_82825 == 32'h0000_0000 ? array_update_83081 : array_update_83070[0];
  assign array_update_83083[1] = add_82825 == 32'h0000_0001 ? array_update_83081 : array_update_83070[1];
  assign array_update_83083[2] = add_82825 == 32'h0000_0002 ? array_update_83081 : array_update_83070[2];
  assign array_update_83083[3] = add_82825 == 32'h0000_0003 ? array_update_83081 : array_update_83070[3];
  assign array_update_83083[4] = add_82825 == 32'h0000_0004 ? array_update_83081 : array_update_83070[4];
  assign array_update_83083[5] = add_82825 == 32'h0000_0005 ? array_update_83081 : array_update_83070[5];
  assign array_update_83083[6] = add_82825 == 32'h0000_0006 ? array_update_83081 : array_update_83070[6];
  assign array_update_83083[7] = add_82825 == 32'h0000_0007 ? array_update_83081 : array_update_83070[7];
  assign array_update_83083[8] = add_82825 == 32'h0000_0008 ? array_update_83081 : array_update_83070[8];
  assign array_update_83083[9] = add_82825 == 32'h0000_0009 ? array_update_83081 : array_update_83070[9];
  assign array_index_83085 = array_update_72021[add_83082 > 32'h0000_0009 ? 4'h9 : add_83082[3:0]];
  assign array_index_83086 = array_update_83083[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_83090 = smul32b_32b_x_32b(array_index_82832[add_83082 > 32'h0000_0009 ? 4'h9 : add_83082[3:0]], array_index_83085[add_82963 > 32'h0000_0009 ? 4'h9 : add_82963[3:0]]);
  assign add_83092 = array_index_83086[add_82963 > 32'h0000_0009 ? 4'h9 : add_82963[3:0]] + smul_83090;
  assign array_update_83093[0] = add_82963 == 32'h0000_0000 ? add_83092 : array_index_83086[0];
  assign array_update_83093[1] = add_82963 == 32'h0000_0001 ? add_83092 : array_index_83086[1];
  assign array_update_83093[2] = add_82963 == 32'h0000_0002 ? add_83092 : array_index_83086[2];
  assign array_update_83093[3] = add_82963 == 32'h0000_0003 ? add_83092 : array_index_83086[3];
  assign array_update_83093[4] = add_82963 == 32'h0000_0004 ? add_83092 : array_index_83086[4];
  assign array_update_83093[5] = add_82963 == 32'h0000_0005 ? add_83092 : array_index_83086[5];
  assign array_update_83093[6] = add_82963 == 32'h0000_0006 ? add_83092 : array_index_83086[6];
  assign array_update_83093[7] = add_82963 == 32'h0000_0007 ? add_83092 : array_index_83086[7];
  assign array_update_83093[8] = add_82963 == 32'h0000_0008 ? add_83092 : array_index_83086[8];
  assign array_update_83093[9] = add_82963 == 32'h0000_0009 ? add_83092 : array_index_83086[9];
  assign array_update_83094[0] = add_82825 == 32'h0000_0000 ? array_update_83093 : array_update_83083[0];
  assign array_update_83094[1] = add_82825 == 32'h0000_0001 ? array_update_83093 : array_update_83083[1];
  assign array_update_83094[2] = add_82825 == 32'h0000_0002 ? array_update_83093 : array_update_83083[2];
  assign array_update_83094[3] = add_82825 == 32'h0000_0003 ? array_update_83093 : array_update_83083[3];
  assign array_update_83094[4] = add_82825 == 32'h0000_0004 ? array_update_83093 : array_update_83083[4];
  assign array_update_83094[5] = add_82825 == 32'h0000_0005 ? array_update_83093 : array_update_83083[5];
  assign array_update_83094[6] = add_82825 == 32'h0000_0006 ? array_update_83093 : array_update_83083[6];
  assign array_update_83094[7] = add_82825 == 32'h0000_0007 ? array_update_83093 : array_update_83083[7];
  assign array_update_83094[8] = add_82825 == 32'h0000_0008 ? array_update_83093 : array_update_83083[8];
  assign array_update_83094[9] = add_82825 == 32'h0000_0009 ? array_update_83093 : array_update_83083[9];
  assign array_index_83096 = array_update_83094[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign add_83098 = add_82963 + 32'h0000_0001;
  assign array_update_83099[0] = add_83098 == 32'h0000_0000 ? 32'h0000_0000 : array_index_83096[0];
  assign array_update_83099[1] = add_83098 == 32'h0000_0001 ? 32'h0000_0000 : array_index_83096[1];
  assign array_update_83099[2] = add_83098 == 32'h0000_0002 ? 32'h0000_0000 : array_index_83096[2];
  assign array_update_83099[3] = add_83098 == 32'h0000_0003 ? 32'h0000_0000 : array_index_83096[3];
  assign array_update_83099[4] = add_83098 == 32'h0000_0004 ? 32'h0000_0000 : array_index_83096[4];
  assign array_update_83099[5] = add_83098 == 32'h0000_0005 ? 32'h0000_0000 : array_index_83096[5];
  assign array_update_83099[6] = add_83098 == 32'h0000_0006 ? 32'h0000_0000 : array_index_83096[6];
  assign array_update_83099[7] = add_83098 == 32'h0000_0007 ? 32'h0000_0000 : array_index_83096[7];
  assign array_update_83099[8] = add_83098 == 32'h0000_0008 ? 32'h0000_0000 : array_index_83096[8];
  assign array_update_83099[9] = add_83098 == 32'h0000_0009 ? 32'h0000_0000 : array_index_83096[9];
  assign literal_83100 = 32'h0000_0000;
  assign array_update_83101[0] = add_82825 == 32'h0000_0000 ? array_update_83099 : array_update_83094[0];
  assign array_update_83101[1] = add_82825 == 32'h0000_0001 ? array_update_83099 : array_update_83094[1];
  assign array_update_83101[2] = add_82825 == 32'h0000_0002 ? array_update_83099 : array_update_83094[2];
  assign array_update_83101[3] = add_82825 == 32'h0000_0003 ? array_update_83099 : array_update_83094[3];
  assign array_update_83101[4] = add_82825 == 32'h0000_0004 ? array_update_83099 : array_update_83094[4];
  assign array_update_83101[5] = add_82825 == 32'h0000_0005 ? array_update_83099 : array_update_83094[5];
  assign array_update_83101[6] = add_82825 == 32'h0000_0006 ? array_update_83099 : array_update_83094[6];
  assign array_update_83101[7] = add_82825 == 32'h0000_0007 ? array_update_83099 : array_update_83094[7];
  assign array_update_83101[8] = add_82825 == 32'h0000_0008 ? array_update_83099 : array_update_83094[8];
  assign array_update_83101[9] = add_82825 == 32'h0000_0009 ? array_update_83099 : array_update_83094[9];
  assign array_index_83103 = array_update_72021[literal_83100 > 32'h0000_0009 ? 4'h9 : literal_83100[3:0]];
  assign array_index_83104 = array_update_83101[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_83108 = smul32b_32b_x_32b(array_index_82832[literal_83100 > 32'h0000_0009 ? 4'h9 : literal_83100[3:0]], array_index_83103[add_83098 > 32'h0000_0009 ? 4'h9 : add_83098[3:0]]);
  assign add_83110 = array_index_83104[add_83098 > 32'h0000_0009 ? 4'h9 : add_83098[3:0]] + smul_83108;
  assign array_update_83112[0] = add_83098 == 32'h0000_0000 ? add_83110 : array_index_83104[0];
  assign array_update_83112[1] = add_83098 == 32'h0000_0001 ? add_83110 : array_index_83104[1];
  assign array_update_83112[2] = add_83098 == 32'h0000_0002 ? add_83110 : array_index_83104[2];
  assign array_update_83112[3] = add_83098 == 32'h0000_0003 ? add_83110 : array_index_83104[3];
  assign array_update_83112[4] = add_83098 == 32'h0000_0004 ? add_83110 : array_index_83104[4];
  assign array_update_83112[5] = add_83098 == 32'h0000_0005 ? add_83110 : array_index_83104[5];
  assign array_update_83112[6] = add_83098 == 32'h0000_0006 ? add_83110 : array_index_83104[6];
  assign array_update_83112[7] = add_83098 == 32'h0000_0007 ? add_83110 : array_index_83104[7];
  assign array_update_83112[8] = add_83098 == 32'h0000_0008 ? add_83110 : array_index_83104[8];
  assign array_update_83112[9] = add_83098 == 32'h0000_0009 ? add_83110 : array_index_83104[9];
  assign add_83113 = literal_83100 + 32'h0000_0001;
  assign array_update_83114[0] = add_82825 == 32'h0000_0000 ? array_update_83112 : array_update_83101[0];
  assign array_update_83114[1] = add_82825 == 32'h0000_0001 ? array_update_83112 : array_update_83101[1];
  assign array_update_83114[2] = add_82825 == 32'h0000_0002 ? array_update_83112 : array_update_83101[2];
  assign array_update_83114[3] = add_82825 == 32'h0000_0003 ? array_update_83112 : array_update_83101[3];
  assign array_update_83114[4] = add_82825 == 32'h0000_0004 ? array_update_83112 : array_update_83101[4];
  assign array_update_83114[5] = add_82825 == 32'h0000_0005 ? array_update_83112 : array_update_83101[5];
  assign array_update_83114[6] = add_82825 == 32'h0000_0006 ? array_update_83112 : array_update_83101[6];
  assign array_update_83114[7] = add_82825 == 32'h0000_0007 ? array_update_83112 : array_update_83101[7];
  assign array_update_83114[8] = add_82825 == 32'h0000_0008 ? array_update_83112 : array_update_83101[8];
  assign array_update_83114[9] = add_82825 == 32'h0000_0009 ? array_update_83112 : array_update_83101[9];
  assign array_index_83116 = array_update_72021[add_83113 > 32'h0000_0009 ? 4'h9 : add_83113[3:0]];
  assign array_index_83117 = array_update_83114[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_83121 = smul32b_32b_x_32b(array_index_82832[add_83113 > 32'h0000_0009 ? 4'h9 : add_83113[3:0]], array_index_83116[add_83098 > 32'h0000_0009 ? 4'h9 : add_83098[3:0]]);
  assign add_83123 = array_index_83117[add_83098 > 32'h0000_0009 ? 4'h9 : add_83098[3:0]] + smul_83121;
  assign array_update_83125[0] = add_83098 == 32'h0000_0000 ? add_83123 : array_index_83117[0];
  assign array_update_83125[1] = add_83098 == 32'h0000_0001 ? add_83123 : array_index_83117[1];
  assign array_update_83125[2] = add_83098 == 32'h0000_0002 ? add_83123 : array_index_83117[2];
  assign array_update_83125[3] = add_83098 == 32'h0000_0003 ? add_83123 : array_index_83117[3];
  assign array_update_83125[4] = add_83098 == 32'h0000_0004 ? add_83123 : array_index_83117[4];
  assign array_update_83125[5] = add_83098 == 32'h0000_0005 ? add_83123 : array_index_83117[5];
  assign array_update_83125[6] = add_83098 == 32'h0000_0006 ? add_83123 : array_index_83117[6];
  assign array_update_83125[7] = add_83098 == 32'h0000_0007 ? add_83123 : array_index_83117[7];
  assign array_update_83125[8] = add_83098 == 32'h0000_0008 ? add_83123 : array_index_83117[8];
  assign array_update_83125[9] = add_83098 == 32'h0000_0009 ? add_83123 : array_index_83117[9];
  assign add_83126 = add_83113 + 32'h0000_0001;
  assign array_update_83127[0] = add_82825 == 32'h0000_0000 ? array_update_83125 : array_update_83114[0];
  assign array_update_83127[1] = add_82825 == 32'h0000_0001 ? array_update_83125 : array_update_83114[1];
  assign array_update_83127[2] = add_82825 == 32'h0000_0002 ? array_update_83125 : array_update_83114[2];
  assign array_update_83127[3] = add_82825 == 32'h0000_0003 ? array_update_83125 : array_update_83114[3];
  assign array_update_83127[4] = add_82825 == 32'h0000_0004 ? array_update_83125 : array_update_83114[4];
  assign array_update_83127[5] = add_82825 == 32'h0000_0005 ? array_update_83125 : array_update_83114[5];
  assign array_update_83127[6] = add_82825 == 32'h0000_0006 ? array_update_83125 : array_update_83114[6];
  assign array_update_83127[7] = add_82825 == 32'h0000_0007 ? array_update_83125 : array_update_83114[7];
  assign array_update_83127[8] = add_82825 == 32'h0000_0008 ? array_update_83125 : array_update_83114[8];
  assign array_update_83127[9] = add_82825 == 32'h0000_0009 ? array_update_83125 : array_update_83114[9];
  assign array_index_83129 = array_update_72021[add_83126 > 32'h0000_0009 ? 4'h9 : add_83126[3:0]];
  assign array_index_83130 = array_update_83127[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_83134 = smul32b_32b_x_32b(array_index_82832[add_83126 > 32'h0000_0009 ? 4'h9 : add_83126[3:0]], array_index_83129[add_83098 > 32'h0000_0009 ? 4'h9 : add_83098[3:0]]);
  assign add_83136 = array_index_83130[add_83098 > 32'h0000_0009 ? 4'h9 : add_83098[3:0]] + smul_83134;
  assign array_update_83138[0] = add_83098 == 32'h0000_0000 ? add_83136 : array_index_83130[0];
  assign array_update_83138[1] = add_83098 == 32'h0000_0001 ? add_83136 : array_index_83130[1];
  assign array_update_83138[2] = add_83098 == 32'h0000_0002 ? add_83136 : array_index_83130[2];
  assign array_update_83138[3] = add_83098 == 32'h0000_0003 ? add_83136 : array_index_83130[3];
  assign array_update_83138[4] = add_83098 == 32'h0000_0004 ? add_83136 : array_index_83130[4];
  assign array_update_83138[5] = add_83098 == 32'h0000_0005 ? add_83136 : array_index_83130[5];
  assign array_update_83138[6] = add_83098 == 32'h0000_0006 ? add_83136 : array_index_83130[6];
  assign array_update_83138[7] = add_83098 == 32'h0000_0007 ? add_83136 : array_index_83130[7];
  assign array_update_83138[8] = add_83098 == 32'h0000_0008 ? add_83136 : array_index_83130[8];
  assign array_update_83138[9] = add_83098 == 32'h0000_0009 ? add_83136 : array_index_83130[9];
  assign add_83139 = add_83126 + 32'h0000_0001;
  assign array_update_83140[0] = add_82825 == 32'h0000_0000 ? array_update_83138 : array_update_83127[0];
  assign array_update_83140[1] = add_82825 == 32'h0000_0001 ? array_update_83138 : array_update_83127[1];
  assign array_update_83140[2] = add_82825 == 32'h0000_0002 ? array_update_83138 : array_update_83127[2];
  assign array_update_83140[3] = add_82825 == 32'h0000_0003 ? array_update_83138 : array_update_83127[3];
  assign array_update_83140[4] = add_82825 == 32'h0000_0004 ? array_update_83138 : array_update_83127[4];
  assign array_update_83140[5] = add_82825 == 32'h0000_0005 ? array_update_83138 : array_update_83127[5];
  assign array_update_83140[6] = add_82825 == 32'h0000_0006 ? array_update_83138 : array_update_83127[6];
  assign array_update_83140[7] = add_82825 == 32'h0000_0007 ? array_update_83138 : array_update_83127[7];
  assign array_update_83140[8] = add_82825 == 32'h0000_0008 ? array_update_83138 : array_update_83127[8];
  assign array_update_83140[9] = add_82825 == 32'h0000_0009 ? array_update_83138 : array_update_83127[9];
  assign array_index_83142 = array_update_72021[add_83139 > 32'h0000_0009 ? 4'h9 : add_83139[3:0]];
  assign array_index_83143 = array_update_83140[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_83147 = smul32b_32b_x_32b(array_index_82832[add_83139 > 32'h0000_0009 ? 4'h9 : add_83139[3:0]], array_index_83142[add_83098 > 32'h0000_0009 ? 4'h9 : add_83098[3:0]]);
  assign add_83149 = array_index_83143[add_83098 > 32'h0000_0009 ? 4'h9 : add_83098[3:0]] + smul_83147;
  assign array_update_83151[0] = add_83098 == 32'h0000_0000 ? add_83149 : array_index_83143[0];
  assign array_update_83151[1] = add_83098 == 32'h0000_0001 ? add_83149 : array_index_83143[1];
  assign array_update_83151[2] = add_83098 == 32'h0000_0002 ? add_83149 : array_index_83143[2];
  assign array_update_83151[3] = add_83098 == 32'h0000_0003 ? add_83149 : array_index_83143[3];
  assign array_update_83151[4] = add_83098 == 32'h0000_0004 ? add_83149 : array_index_83143[4];
  assign array_update_83151[5] = add_83098 == 32'h0000_0005 ? add_83149 : array_index_83143[5];
  assign array_update_83151[6] = add_83098 == 32'h0000_0006 ? add_83149 : array_index_83143[6];
  assign array_update_83151[7] = add_83098 == 32'h0000_0007 ? add_83149 : array_index_83143[7];
  assign array_update_83151[8] = add_83098 == 32'h0000_0008 ? add_83149 : array_index_83143[8];
  assign array_update_83151[9] = add_83098 == 32'h0000_0009 ? add_83149 : array_index_83143[9];
  assign add_83152 = add_83139 + 32'h0000_0001;
  assign array_update_83153[0] = add_82825 == 32'h0000_0000 ? array_update_83151 : array_update_83140[0];
  assign array_update_83153[1] = add_82825 == 32'h0000_0001 ? array_update_83151 : array_update_83140[1];
  assign array_update_83153[2] = add_82825 == 32'h0000_0002 ? array_update_83151 : array_update_83140[2];
  assign array_update_83153[3] = add_82825 == 32'h0000_0003 ? array_update_83151 : array_update_83140[3];
  assign array_update_83153[4] = add_82825 == 32'h0000_0004 ? array_update_83151 : array_update_83140[4];
  assign array_update_83153[5] = add_82825 == 32'h0000_0005 ? array_update_83151 : array_update_83140[5];
  assign array_update_83153[6] = add_82825 == 32'h0000_0006 ? array_update_83151 : array_update_83140[6];
  assign array_update_83153[7] = add_82825 == 32'h0000_0007 ? array_update_83151 : array_update_83140[7];
  assign array_update_83153[8] = add_82825 == 32'h0000_0008 ? array_update_83151 : array_update_83140[8];
  assign array_update_83153[9] = add_82825 == 32'h0000_0009 ? array_update_83151 : array_update_83140[9];
  assign array_index_83155 = array_update_72021[add_83152 > 32'h0000_0009 ? 4'h9 : add_83152[3:0]];
  assign array_index_83156 = array_update_83153[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_83160 = smul32b_32b_x_32b(array_index_82832[add_83152 > 32'h0000_0009 ? 4'h9 : add_83152[3:0]], array_index_83155[add_83098 > 32'h0000_0009 ? 4'h9 : add_83098[3:0]]);
  assign add_83162 = array_index_83156[add_83098 > 32'h0000_0009 ? 4'h9 : add_83098[3:0]] + smul_83160;
  assign array_update_83164[0] = add_83098 == 32'h0000_0000 ? add_83162 : array_index_83156[0];
  assign array_update_83164[1] = add_83098 == 32'h0000_0001 ? add_83162 : array_index_83156[1];
  assign array_update_83164[2] = add_83098 == 32'h0000_0002 ? add_83162 : array_index_83156[2];
  assign array_update_83164[3] = add_83098 == 32'h0000_0003 ? add_83162 : array_index_83156[3];
  assign array_update_83164[4] = add_83098 == 32'h0000_0004 ? add_83162 : array_index_83156[4];
  assign array_update_83164[5] = add_83098 == 32'h0000_0005 ? add_83162 : array_index_83156[5];
  assign array_update_83164[6] = add_83098 == 32'h0000_0006 ? add_83162 : array_index_83156[6];
  assign array_update_83164[7] = add_83098 == 32'h0000_0007 ? add_83162 : array_index_83156[7];
  assign array_update_83164[8] = add_83098 == 32'h0000_0008 ? add_83162 : array_index_83156[8];
  assign array_update_83164[9] = add_83098 == 32'h0000_0009 ? add_83162 : array_index_83156[9];
  assign add_83165 = add_83152 + 32'h0000_0001;
  assign array_update_83166[0] = add_82825 == 32'h0000_0000 ? array_update_83164 : array_update_83153[0];
  assign array_update_83166[1] = add_82825 == 32'h0000_0001 ? array_update_83164 : array_update_83153[1];
  assign array_update_83166[2] = add_82825 == 32'h0000_0002 ? array_update_83164 : array_update_83153[2];
  assign array_update_83166[3] = add_82825 == 32'h0000_0003 ? array_update_83164 : array_update_83153[3];
  assign array_update_83166[4] = add_82825 == 32'h0000_0004 ? array_update_83164 : array_update_83153[4];
  assign array_update_83166[5] = add_82825 == 32'h0000_0005 ? array_update_83164 : array_update_83153[5];
  assign array_update_83166[6] = add_82825 == 32'h0000_0006 ? array_update_83164 : array_update_83153[6];
  assign array_update_83166[7] = add_82825 == 32'h0000_0007 ? array_update_83164 : array_update_83153[7];
  assign array_update_83166[8] = add_82825 == 32'h0000_0008 ? array_update_83164 : array_update_83153[8];
  assign array_update_83166[9] = add_82825 == 32'h0000_0009 ? array_update_83164 : array_update_83153[9];
  assign array_index_83168 = array_update_72021[add_83165 > 32'h0000_0009 ? 4'h9 : add_83165[3:0]];
  assign array_index_83169 = array_update_83166[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_83173 = smul32b_32b_x_32b(array_index_82832[add_83165 > 32'h0000_0009 ? 4'h9 : add_83165[3:0]], array_index_83168[add_83098 > 32'h0000_0009 ? 4'h9 : add_83098[3:0]]);
  assign add_83175 = array_index_83169[add_83098 > 32'h0000_0009 ? 4'h9 : add_83098[3:0]] + smul_83173;
  assign array_update_83177[0] = add_83098 == 32'h0000_0000 ? add_83175 : array_index_83169[0];
  assign array_update_83177[1] = add_83098 == 32'h0000_0001 ? add_83175 : array_index_83169[1];
  assign array_update_83177[2] = add_83098 == 32'h0000_0002 ? add_83175 : array_index_83169[2];
  assign array_update_83177[3] = add_83098 == 32'h0000_0003 ? add_83175 : array_index_83169[3];
  assign array_update_83177[4] = add_83098 == 32'h0000_0004 ? add_83175 : array_index_83169[4];
  assign array_update_83177[5] = add_83098 == 32'h0000_0005 ? add_83175 : array_index_83169[5];
  assign array_update_83177[6] = add_83098 == 32'h0000_0006 ? add_83175 : array_index_83169[6];
  assign array_update_83177[7] = add_83098 == 32'h0000_0007 ? add_83175 : array_index_83169[7];
  assign array_update_83177[8] = add_83098 == 32'h0000_0008 ? add_83175 : array_index_83169[8];
  assign array_update_83177[9] = add_83098 == 32'h0000_0009 ? add_83175 : array_index_83169[9];
  assign add_83178 = add_83165 + 32'h0000_0001;
  assign array_update_83179[0] = add_82825 == 32'h0000_0000 ? array_update_83177 : array_update_83166[0];
  assign array_update_83179[1] = add_82825 == 32'h0000_0001 ? array_update_83177 : array_update_83166[1];
  assign array_update_83179[2] = add_82825 == 32'h0000_0002 ? array_update_83177 : array_update_83166[2];
  assign array_update_83179[3] = add_82825 == 32'h0000_0003 ? array_update_83177 : array_update_83166[3];
  assign array_update_83179[4] = add_82825 == 32'h0000_0004 ? array_update_83177 : array_update_83166[4];
  assign array_update_83179[5] = add_82825 == 32'h0000_0005 ? array_update_83177 : array_update_83166[5];
  assign array_update_83179[6] = add_82825 == 32'h0000_0006 ? array_update_83177 : array_update_83166[6];
  assign array_update_83179[7] = add_82825 == 32'h0000_0007 ? array_update_83177 : array_update_83166[7];
  assign array_update_83179[8] = add_82825 == 32'h0000_0008 ? array_update_83177 : array_update_83166[8];
  assign array_update_83179[9] = add_82825 == 32'h0000_0009 ? array_update_83177 : array_update_83166[9];
  assign array_index_83181 = array_update_72021[add_83178 > 32'h0000_0009 ? 4'h9 : add_83178[3:0]];
  assign array_index_83182 = array_update_83179[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_83186 = smul32b_32b_x_32b(array_index_82832[add_83178 > 32'h0000_0009 ? 4'h9 : add_83178[3:0]], array_index_83181[add_83098 > 32'h0000_0009 ? 4'h9 : add_83098[3:0]]);
  assign add_83188 = array_index_83182[add_83098 > 32'h0000_0009 ? 4'h9 : add_83098[3:0]] + smul_83186;
  assign array_update_83190[0] = add_83098 == 32'h0000_0000 ? add_83188 : array_index_83182[0];
  assign array_update_83190[1] = add_83098 == 32'h0000_0001 ? add_83188 : array_index_83182[1];
  assign array_update_83190[2] = add_83098 == 32'h0000_0002 ? add_83188 : array_index_83182[2];
  assign array_update_83190[3] = add_83098 == 32'h0000_0003 ? add_83188 : array_index_83182[3];
  assign array_update_83190[4] = add_83098 == 32'h0000_0004 ? add_83188 : array_index_83182[4];
  assign array_update_83190[5] = add_83098 == 32'h0000_0005 ? add_83188 : array_index_83182[5];
  assign array_update_83190[6] = add_83098 == 32'h0000_0006 ? add_83188 : array_index_83182[6];
  assign array_update_83190[7] = add_83098 == 32'h0000_0007 ? add_83188 : array_index_83182[7];
  assign array_update_83190[8] = add_83098 == 32'h0000_0008 ? add_83188 : array_index_83182[8];
  assign array_update_83190[9] = add_83098 == 32'h0000_0009 ? add_83188 : array_index_83182[9];
  assign add_83191 = add_83178 + 32'h0000_0001;
  assign array_update_83192[0] = add_82825 == 32'h0000_0000 ? array_update_83190 : array_update_83179[0];
  assign array_update_83192[1] = add_82825 == 32'h0000_0001 ? array_update_83190 : array_update_83179[1];
  assign array_update_83192[2] = add_82825 == 32'h0000_0002 ? array_update_83190 : array_update_83179[2];
  assign array_update_83192[3] = add_82825 == 32'h0000_0003 ? array_update_83190 : array_update_83179[3];
  assign array_update_83192[4] = add_82825 == 32'h0000_0004 ? array_update_83190 : array_update_83179[4];
  assign array_update_83192[5] = add_82825 == 32'h0000_0005 ? array_update_83190 : array_update_83179[5];
  assign array_update_83192[6] = add_82825 == 32'h0000_0006 ? array_update_83190 : array_update_83179[6];
  assign array_update_83192[7] = add_82825 == 32'h0000_0007 ? array_update_83190 : array_update_83179[7];
  assign array_update_83192[8] = add_82825 == 32'h0000_0008 ? array_update_83190 : array_update_83179[8];
  assign array_update_83192[9] = add_82825 == 32'h0000_0009 ? array_update_83190 : array_update_83179[9];
  assign array_index_83194 = array_update_72021[add_83191 > 32'h0000_0009 ? 4'h9 : add_83191[3:0]];
  assign array_index_83195 = array_update_83192[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_83199 = smul32b_32b_x_32b(array_index_82832[add_83191 > 32'h0000_0009 ? 4'h9 : add_83191[3:0]], array_index_83194[add_83098 > 32'h0000_0009 ? 4'h9 : add_83098[3:0]]);
  assign add_83201 = array_index_83195[add_83098 > 32'h0000_0009 ? 4'h9 : add_83098[3:0]] + smul_83199;
  assign array_update_83203[0] = add_83098 == 32'h0000_0000 ? add_83201 : array_index_83195[0];
  assign array_update_83203[1] = add_83098 == 32'h0000_0001 ? add_83201 : array_index_83195[1];
  assign array_update_83203[2] = add_83098 == 32'h0000_0002 ? add_83201 : array_index_83195[2];
  assign array_update_83203[3] = add_83098 == 32'h0000_0003 ? add_83201 : array_index_83195[3];
  assign array_update_83203[4] = add_83098 == 32'h0000_0004 ? add_83201 : array_index_83195[4];
  assign array_update_83203[5] = add_83098 == 32'h0000_0005 ? add_83201 : array_index_83195[5];
  assign array_update_83203[6] = add_83098 == 32'h0000_0006 ? add_83201 : array_index_83195[6];
  assign array_update_83203[7] = add_83098 == 32'h0000_0007 ? add_83201 : array_index_83195[7];
  assign array_update_83203[8] = add_83098 == 32'h0000_0008 ? add_83201 : array_index_83195[8];
  assign array_update_83203[9] = add_83098 == 32'h0000_0009 ? add_83201 : array_index_83195[9];
  assign add_83204 = add_83191 + 32'h0000_0001;
  assign array_update_83205[0] = add_82825 == 32'h0000_0000 ? array_update_83203 : array_update_83192[0];
  assign array_update_83205[1] = add_82825 == 32'h0000_0001 ? array_update_83203 : array_update_83192[1];
  assign array_update_83205[2] = add_82825 == 32'h0000_0002 ? array_update_83203 : array_update_83192[2];
  assign array_update_83205[3] = add_82825 == 32'h0000_0003 ? array_update_83203 : array_update_83192[3];
  assign array_update_83205[4] = add_82825 == 32'h0000_0004 ? array_update_83203 : array_update_83192[4];
  assign array_update_83205[5] = add_82825 == 32'h0000_0005 ? array_update_83203 : array_update_83192[5];
  assign array_update_83205[6] = add_82825 == 32'h0000_0006 ? array_update_83203 : array_update_83192[6];
  assign array_update_83205[7] = add_82825 == 32'h0000_0007 ? array_update_83203 : array_update_83192[7];
  assign array_update_83205[8] = add_82825 == 32'h0000_0008 ? array_update_83203 : array_update_83192[8];
  assign array_update_83205[9] = add_82825 == 32'h0000_0009 ? array_update_83203 : array_update_83192[9];
  assign array_index_83207 = array_update_72021[add_83204 > 32'h0000_0009 ? 4'h9 : add_83204[3:0]];
  assign array_index_83208 = array_update_83205[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_83212 = smul32b_32b_x_32b(array_index_82832[add_83204 > 32'h0000_0009 ? 4'h9 : add_83204[3:0]], array_index_83207[add_83098 > 32'h0000_0009 ? 4'h9 : add_83098[3:0]]);
  assign add_83214 = array_index_83208[add_83098 > 32'h0000_0009 ? 4'h9 : add_83098[3:0]] + smul_83212;
  assign array_update_83216[0] = add_83098 == 32'h0000_0000 ? add_83214 : array_index_83208[0];
  assign array_update_83216[1] = add_83098 == 32'h0000_0001 ? add_83214 : array_index_83208[1];
  assign array_update_83216[2] = add_83098 == 32'h0000_0002 ? add_83214 : array_index_83208[2];
  assign array_update_83216[3] = add_83098 == 32'h0000_0003 ? add_83214 : array_index_83208[3];
  assign array_update_83216[4] = add_83098 == 32'h0000_0004 ? add_83214 : array_index_83208[4];
  assign array_update_83216[5] = add_83098 == 32'h0000_0005 ? add_83214 : array_index_83208[5];
  assign array_update_83216[6] = add_83098 == 32'h0000_0006 ? add_83214 : array_index_83208[6];
  assign array_update_83216[7] = add_83098 == 32'h0000_0007 ? add_83214 : array_index_83208[7];
  assign array_update_83216[8] = add_83098 == 32'h0000_0008 ? add_83214 : array_index_83208[8];
  assign array_update_83216[9] = add_83098 == 32'h0000_0009 ? add_83214 : array_index_83208[9];
  assign add_83217 = add_83204 + 32'h0000_0001;
  assign array_update_83218[0] = add_82825 == 32'h0000_0000 ? array_update_83216 : array_update_83205[0];
  assign array_update_83218[1] = add_82825 == 32'h0000_0001 ? array_update_83216 : array_update_83205[1];
  assign array_update_83218[2] = add_82825 == 32'h0000_0002 ? array_update_83216 : array_update_83205[2];
  assign array_update_83218[3] = add_82825 == 32'h0000_0003 ? array_update_83216 : array_update_83205[3];
  assign array_update_83218[4] = add_82825 == 32'h0000_0004 ? array_update_83216 : array_update_83205[4];
  assign array_update_83218[5] = add_82825 == 32'h0000_0005 ? array_update_83216 : array_update_83205[5];
  assign array_update_83218[6] = add_82825 == 32'h0000_0006 ? array_update_83216 : array_update_83205[6];
  assign array_update_83218[7] = add_82825 == 32'h0000_0007 ? array_update_83216 : array_update_83205[7];
  assign array_update_83218[8] = add_82825 == 32'h0000_0008 ? array_update_83216 : array_update_83205[8];
  assign array_update_83218[9] = add_82825 == 32'h0000_0009 ? array_update_83216 : array_update_83205[9];
  assign array_index_83220 = array_update_72021[add_83217 > 32'h0000_0009 ? 4'h9 : add_83217[3:0]];
  assign array_index_83221 = array_update_83218[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_83225 = smul32b_32b_x_32b(array_index_82832[add_83217 > 32'h0000_0009 ? 4'h9 : add_83217[3:0]], array_index_83220[add_83098 > 32'h0000_0009 ? 4'h9 : add_83098[3:0]]);
  assign add_83227 = array_index_83221[add_83098 > 32'h0000_0009 ? 4'h9 : add_83098[3:0]] + smul_83225;
  assign array_update_83228[0] = add_83098 == 32'h0000_0000 ? add_83227 : array_index_83221[0];
  assign array_update_83228[1] = add_83098 == 32'h0000_0001 ? add_83227 : array_index_83221[1];
  assign array_update_83228[2] = add_83098 == 32'h0000_0002 ? add_83227 : array_index_83221[2];
  assign array_update_83228[3] = add_83098 == 32'h0000_0003 ? add_83227 : array_index_83221[3];
  assign array_update_83228[4] = add_83098 == 32'h0000_0004 ? add_83227 : array_index_83221[4];
  assign array_update_83228[5] = add_83098 == 32'h0000_0005 ? add_83227 : array_index_83221[5];
  assign array_update_83228[6] = add_83098 == 32'h0000_0006 ? add_83227 : array_index_83221[6];
  assign array_update_83228[7] = add_83098 == 32'h0000_0007 ? add_83227 : array_index_83221[7];
  assign array_update_83228[8] = add_83098 == 32'h0000_0008 ? add_83227 : array_index_83221[8];
  assign array_update_83228[9] = add_83098 == 32'h0000_0009 ? add_83227 : array_index_83221[9];
  assign array_update_83229[0] = add_82825 == 32'h0000_0000 ? array_update_83228 : array_update_83218[0];
  assign array_update_83229[1] = add_82825 == 32'h0000_0001 ? array_update_83228 : array_update_83218[1];
  assign array_update_83229[2] = add_82825 == 32'h0000_0002 ? array_update_83228 : array_update_83218[2];
  assign array_update_83229[3] = add_82825 == 32'h0000_0003 ? array_update_83228 : array_update_83218[3];
  assign array_update_83229[4] = add_82825 == 32'h0000_0004 ? array_update_83228 : array_update_83218[4];
  assign array_update_83229[5] = add_82825 == 32'h0000_0005 ? array_update_83228 : array_update_83218[5];
  assign array_update_83229[6] = add_82825 == 32'h0000_0006 ? array_update_83228 : array_update_83218[6];
  assign array_update_83229[7] = add_82825 == 32'h0000_0007 ? array_update_83228 : array_update_83218[7];
  assign array_update_83229[8] = add_82825 == 32'h0000_0008 ? array_update_83228 : array_update_83218[8];
  assign array_update_83229[9] = add_82825 == 32'h0000_0009 ? array_update_83228 : array_update_83218[9];
  assign array_index_83231 = array_update_83229[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign add_83233 = add_83098 + 32'h0000_0001;
  assign array_update_83234[0] = add_83233 == 32'h0000_0000 ? 32'h0000_0000 : array_index_83231[0];
  assign array_update_83234[1] = add_83233 == 32'h0000_0001 ? 32'h0000_0000 : array_index_83231[1];
  assign array_update_83234[2] = add_83233 == 32'h0000_0002 ? 32'h0000_0000 : array_index_83231[2];
  assign array_update_83234[3] = add_83233 == 32'h0000_0003 ? 32'h0000_0000 : array_index_83231[3];
  assign array_update_83234[4] = add_83233 == 32'h0000_0004 ? 32'h0000_0000 : array_index_83231[4];
  assign array_update_83234[5] = add_83233 == 32'h0000_0005 ? 32'h0000_0000 : array_index_83231[5];
  assign array_update_83234[6] = add_83233 == 32'h0000_0006 ? 32'h0000_0000 : array_index_83231[6];
  assign array_update_83234[7] = add_83233 == 32'h0000_0007 ? 32'h0000_0000 : array_index_83231[7];
  assign array_update_83234[8] = add_83233 == 32'h0000_0008 ? 32'h0000_0000 : array_index_83231[8];
  assign array_update_83234[9] = add_83233 == 32'h0000_0009 ? 32'h0000_0000 : array_index_83231[9];
  assign literal_83235 = 32'h0000_0000;
  assign array_update_83236[0] = add_82825 == 32'h0000_0000 ? array_update_83234 : array_update_83229[0];
  assign array_update_83236[1] = add_82825 == 32'h0000_0001 ? array_update_83234 : array_update_83229[1];
  assign array_update_83236[2] = add_82825 == 32'h0000_0002 ? array_update_83234 : array_update_83229[2];
  assign array_update_83236[3] = add_82825 == 32'h0000_0003 ? array_update_83234 : array_update_83229[3];
  assign array_update_83236[4] = add_82825 == 32'h0000_0004 ? array_update_83234 : array_update_83229[4];
  assign array_update_83236[5] = add_82825 == 32'h0000_0005 ? array_update_83234 : array_update_83229[5];
  assign array_update_83236[6] = add_82825 == 32'h0000_0006 ? array_update_83234 : array_update_83229[6];
  assign array_update_83236[7] = add_82825 == 32'h0000_0007 ? array_update_83234 : array_update_83229[7];
  assign array_update_83236[8] = add_82825 == 32'h0000_0008 ? array_update_83234 : array_update_83229[8];
  assign array_update_83236[9] = add_82825 == 32'h0000_0009 ? array_update_83234 : array_update_83229[9];
  assign array_index_83238 = array_update_72021[literal_83235 > 32'h0000_0009 ? 4'h9 : literal_83235[3:0]];
  assign array_index_83239 = array_update_83236[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_83243 = smul32b_32b_x_32b(array_index_82832[literal_83235 > 32'h0000_0009 ? 4'h9 : literal_83235[3:0]], array_index_83238[add_83233 > 32'h0000_0009 ? 4'h9 : add_83233[3:0]]);
  assign add_83245 = array_index_83239[add_83233 > 32'h0000_0009 ? 4'h9 : add_83233[3:0]] + smul_83243;
  assign array_update_83247[0] = add_83233 == 32'h0000_0000 ? add_83245 : array_index_83239[0];
  assign array_update_83247[1] = add_83233 == 32'h0000_0001 ? add_83245 : array_index_83239[1];
  assign array_update_83247[2] = add_83233 == 32'h0000_0002 ? add_83245 : array_index_83239[2];
  assign array_update_83247[3] = add_83233 == 32'h0000_0003 ? add_83245 : array_index_83239[3];
  assign array_update_83247[4] = add_83233 == 32'h0000_0004 ? add_83245 : array_index_83239[4];
  assign array_update_83247[5] = add_83233 == 32'h0000_0005 ? add_83245 : array_index_83239[5];
  assign array_update_83247[6] = add_83233 == 32'h0000_0006 ? add_83245 : array_index_83239[6];
  assign array_update_83247[7] = add_83233 == 32'h0000_0007 ? add_83245 : array_index_83239[7];
  assign array_update_83247[8] = add_83233 == 32'h0000_0008 ? add_83245 : array_index_83239[8];
  assign array_update_83247[9] = add_83233 == 32'h0000_0009 ? add_83245 : array_index_83239[9];
  assign add_83248 = literal_83235 + 32'h0000_0001;
  assign array_update_83249[0] = add_82825 == 32'h0000_0000 ? array_update_83247 : array_update_83236[0];
  assign array_update_83249[1] = add_82825 == 32'h0000_0001 ? array_update_83247 : array_update_83236[1];
  assign array_update_83249[2] = add_82825 == 32'h0000_0002 ? array_update_83247 : array_update_83236[2];
  assign array_update_83249[3] = add_82825 == 32'h0000_0003 ? array_update_83247 : array_update_83236[3];
  assign array_update_83249[4] = add_82825 == 32'h0000_0004 ? array_update_83247 : array_update_83236[4];
  assign array_update_83249[5] = add_82825 == 32'h0000_0005 ? array_update_83247 : array_update_83236[5];
  assign array_update_83249[6] = add_82825 == 32'h0000_0006 ? array_update_83247 : array_update_83236[6];
  assign array_update_83249[7] = add_82825 == 32'h0000_0007 ? array_update_83247 : array_update_83236[7];
  assign array_update_83249[8] = add_82825 == 32'h0000_0008 ? array_update_83247 : array_update_83236[8];
  assign array_update_83249[9] = add_82825 == 32'h0000_0009 ? array_update_83247 : array_update_83236[9];
  assign array_index_83251 = array_update_72021[add_83248 > 32'h0000_0009 ? 4'h9 : add_83248[3:0]];
  assign array_index_83252 = array_update_83249[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_83256 = smul32b_32b_x_32b(array_index_82832[add_83248 > 32'h0000_0009 ? 4'h9 : add_83248[3:0]], array_index_83251[add_83233 > 32'h0000_0009 ? 4'h9 : add_83233[3:0]]);
  assign add_83258 = array_index_83252[add_83233 > 32'h0000_0009 ? 4'h9 : add_83233[3:0]] + smul_83256;
  assign array_update_83260[0] = add_83233 == 32'h0000_0000 ? add_83258 : array_index_83252[0];
  assign array_update_83260[1] = add_83233 == 32'h0000_0001 ? add_83258 : array_index_83252[1];
  assign array_update_83260[2] = add_83233 == 32'h0000_0002 ? add_83258 : array_index_83252[2];
  assign array_update_83260[3] = add_83233 == 32'h0000_0003 ? add_83258 : array_index_83252[3];
  assign array_update_83260[4] = add_83233 == 32'h0000_0004 ? add_83258 : array_index_83252[4];
  assign array_update_83260[5] = add_83233 == 32'h0000_0005 ? add_83258 : array_index_83252[5];
  assign array_update_83260[6] = add_83233 == 32'h0000_0006 ? add_83258 : array_index_83252[6];
  assign array_update_83260[7] = add_83233 == 32'h0000_0007 ? add_83258 : array_index_83252[7];
  assign array_update_83260[8] = add_83233 == 32'h0000_0008 ? add_83258 : array_index_83252[8];
  assign array_update_83260[9] = add_83233 == 32'h0000_0009 ? add_83258 : array_index_83252[9];
  assign add_83261 = add_83248 + 32'h0000_0001;
  assign array_update_83262[0] = add_82825 == 32'h0000_0000 ? array_update_83260 : array_update_83249[0];
  assign array_update_83262[1] = add_82825 == 32'h0000_0001 ? array_update_83260 : array_update_83249[1];
  assign array_update_83262[2] = add_82825 == 32'h0000_0002 ? array_update_83260 : array_update_83249[2];
  assign array_update_83262[3] = add_82825 == 32'h0000_0003 ? array_update_83260 : array_update_83249[3];
  assign array_update_83262[4] = add_82825 == 32'h0000_0004 ? array_update_83260 : array_update_83249[4];
  assign array_update_83262[5] = add_82825 == 32'h0000_0005 ? array_update_83260 : array_update_83249[5];
  assign array_update_83262[6] = add_82825 == 32'h0000_0006 ? array_update_83260 : array_update_83249[6];
  assign array_update_83262[7] = add_82825 == 32'h0000_0007 ? array_update_83260 : array_update_83249[7];
  assign array_update_83262[8] = add_82825 == 32'h0000_0008 ? array_update_83260 : array_update_83249[8];
  assign array_update_83262[9] = add_82825 == 32'h0000_0009 ? array_update_83260 : array_update_83249[9];
  assign array_index_83264 = array_update_72021[add_83261 > 32'h0000_0009 ? 4'h9 : add_83261[3:0]];
  assign array_index_83265 = array_update_83262[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_83269 = smul32b_32b_x_32b(array_index_82832[add_83261 > 32'h0000_0009 ? 4'h9 : add_83261[3:0]], array_index_83264[add_83233 > 32'h0000_0009 ? 4'h9 : add_83233[3:0]]);
  assign add_83271 = array_index_83265[add_83233 > 32'h0000_0009 ? 4'h9 : add_83233[3:0]] + smul_83269;
  assign array_update_83273[0] = add_83233 == 32'h0000_0000 ? add_83271 : array_index_83265[0];
  assign array_update_83273[1] = add_83233 == 32'h0000_0001 ? add_83271 : array_index_83265[1];
  assign array_update_83273[2] = add_83233 == 32'h0000_0002 ? add_83271 : array_index_83265[2];
  assign array_update_83273[3] = add_83233 == 32'h0000_0003 ? add_83271 : array_index_83265[3];
  assign array_update_83273[4] = add_83233 == 32'h0000_0004 ? add_83271 : array_index_83265[4];
  assign array_update_83273[5] = add_83233 == 32'h0000_0005 ? add_83271 : array_index_83265[5];
  assign array_update_83273[6] = add_83233 == 32'h0000_0006 ? add_83271 : array_index_83265[6];
  assign array_update_83273[7] = add_83233 == 32'h0000_0007 ? add_83271 : array_index_83265[7];
  assign array_update_83273[8] = add_83233 == 32'h0000_0008 ? add_83271 : array_index_83265[8];
  assign array_update_83273[9] = add_83233 == 32'h0000_0009 ? add_83271 : array_index_83265[9];
  assign add_83274 = add_83261 + 32'h0000_0001;
  assign array_update_83275[0] = add_82825 == 32'h0000_0000 ? array_update_83273 : array_update_83262[0];
  assign array_update_83275[1] = add_82825 == 32'h0000_0001 ? array_update_83273 : array_update_83262[1];
  assign array_update_83275[2] = add_82825 == 32'h0000_0002 ? array_update_83273 : array_update_83262[2];
  assign array_update_83275[3] = add_82825 == 32'h0000_0003 ? array_update_83273 : array_update_83262[3];
  assign array_update_83275[4] = add_82825 == 32'h0000_0004 ? array_update_83273 : array_update_83262[4];
  assign array_update_83275[5] = add_82825 == 32'h0000_0005 ? array_update_83273 : array_update_83262[5];
  assign array_update_83275[6] = add_82825 == 32'h0000_0006 ? array_update_83273 : array_update_83262[6];
  assign array_update_83275[7] = add_82825 == 32'h0000_0007 ? array_update_83273 : array_update_83262[7];
  assign array_update_83275[8] = add_82825 == 32'h0000_0008 ? array_update_83273 : array_update_83262[8];
  assign array_update_83275[9] = add_82825 == 32'h0000_0009 ? array_update_83273 : array_update_83262[9];
  assign array_index_83277 = array_update_72021[add_83274 > 32'h0000_0009 ? 4'h9 : add_83274[3:0]];
  assign array_index_83278 = array_update_83275[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_83282 = smul32b_32b_x_32b(array_index_82832[add_83274 > 32'h0000_0009 ? 4'h9 : add_83274[3:0]], array_index_83277[add_83233 > 32'h0000_0009 ? 4'h9 : add_83233[3:0]]);
  assign add_83284 = array_index_83278[add_83233 > 32'h0000_0009 ? 4'h9 : add_83233[3:0]] + smul_83282;
  assign array_update_83286[0] = add_83233 == 32'h0000_0000 ? add_83284 : array_index_83278[0];
  assign array_update_83286[1] = add_83233 == 32'h0000_0001 ? add_83284 : array_index_83278[1];
  assign array_update_83286[2] = add_83233 == 32'h0000_0002 ? add_83284 : array_index_83278[2];
  assign array_update_83286[3] = add_83233 == 32'h0000_0003 ? add_83284 : array_index_83278[3];
  assign array_update_83286[4] = add_83233 == 32'h0000_0004 ? add_83284 : array_index_83278[4];
  assign array_update_83286[5] = add_83233 == 32'h0000_0005 ? add_83284 : array_index_83278[5];
  assign array_update_83286[6] = add_83233 == 32'h0000_0006 ? add_83284 : array_index_83278[6];
  assign array_update_83286[7] = add_83233 == 32'h0000_0007 ? add_83284 : array_index_83278[7];
  assign array_update_83286[8] = add_83233 == 32'h0000_0008 ? add_83284 : array_index_83278[8];
  assign array_update_83286[9] = add_83233 == 32'h0000_0009 ? add_83284 : array_index_83278[9];
  assign add_83287 = add_83274 + 32'h0000_0001;
  assign array_update_83288[0] = add_82825 == 32'h0000_0000 ? array_update_83286 : array_update_83275[0];
  assign array_update_83288[1] = add_82825 == 32'h0000_0001 ? array_update_83286 : array_update_83275[1];
  assign array_update_83288[2] = add_82825 == 32'h0000_0002 ? array_update_83286 : array_update_83275[2];
  assign array_update_83288[3] = add_82825 == 32'h0000_0003 ? array_update_83286 : array_update_83275[3];
  assign array_update_83288[4] = add_82825 == 32'h0000_0004 ? array_update_83286 : array_update_83275[4];
  assign array_update_83288[5] = add_82825 == 32'h0000_0005 ? array_update_83286 : array_update_83275[5];
  assign array_update_83288[6] = add_82825 == 32'h0000_0006 ? array_update_83286 : array_update_83275[6];
  assign array_update_83288[7] = add_82825 == 32'h0000_0007 ? array_update_83286 : array_update_83275[7];
  assign array_update_83288[8] = add_82825 == 32'h0000_0008 ? array_update_83286 : array_update_83275[8];
  assign array_update_83288[9] = add_82825 == 32'h0000_0009 ? array_update_83286 : array_update_83275[9];
  assign array_index_83290 = array_update_72021[add_83287 > 32'h0000_0009 ? 4'h9 : add_83287[3:0]];
  assign array_index_83291 = array_update_83288[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_83295 = smul32b_32b_x_32b(array_index_82832[add_83287 > 32'h0000_0009 ? 4'h9 : add_83287[3:0]], array_index_83290[add_83233 > 32'h0000_0009 ? 4'h9 : add_83233[3:0]]);
  assign add_83297 = array_index_83291[add_83233 > 32'h0000_0009 ? 4'h9 : add_83233[3:0]] + smul_83295;
  assign array_update_83299[0] = add_83233 == 32'h0000_0000 ? add_83297 : array_index_83291[0];
  assign array_update_83299[1] = add_83233 == 32'h0000_0001 ? add_83297 : array_index_83291[1];
  assign array_update_83299[2] = add_83233 == 32'h0000_0002 ? add_83297 : array_index_83291[2];
  assign array_update_83299[3] = add_83233 == 32'h0000_0003 ? add_83297 : array_index_83291[3];
  assign array_update_83299[4] = add_83233 == 32'h0000_0004 ? add_83297 : array_index_83291[4];
  assign array_update_83299[5] = add_83233 == 32'h0000_0005 ? add_83297 : array_index_83291[5];
  assign array_update_83299[6] = add_83233 == 32'h0000_0006 ? add_83297 : array_index_83291[6];
  assign array_update_83299[7] = add_83233 == 32'h0000_0007 ? add_83297 : array_index_83291[7];
  assign array_update_83299[8] = add_83233 == 32'h0000_0008 ? add_83297 : array_index_83291[8];
  assign array_update_83299[9] = add_83233 == 32'h0000_0009 ? add_83297 : array_index_83291[9];
  assign add_83300 = add_83287 + 32'h0000_0001;
  assign array_update_83301[0] = add_82825 == 32'h0000_0000 ? array_update_83299 : array_update_83288[0];
  assign array_update_83301[1] = add_82825 == 32'h0000_0001 ? array_update_83299 : array_update_83288[1];
  assign array_update_83301[2] = add_82825 == 32'h0000_0002 ? array_update_83299 : array_update_83288[2];
  assign array_update_83301[3] = add_82825 == 32'h0000_0003 ? array_update_83299 : array_update_83288[3];
  assign array_update_83301[4] = add_82825 == 32'h0000_0004 ? array_update_83299 : array_update_83288[4];
  assign array_update_83301[5] = add_82825 == 32'h0000_0005 ? array_update_83299 : array_update_83288[5];
  assign array_update_83301[6] = add_82825 == 32'h0000_0006 ? array_update_83299 : array_update_83288[6];
  assign array_update_83301[7] = add_82825 == 32'h0000_0007 ? array_update_83299 : array_update_83288[7];
  assign array_update_83301[8] = add_82825 == 32'h0000_0008 ? array_update_83299 : array_update_83288[8];
  assign array_update_83301[9] = add_82825 == 32'h0000_0009 ? array_update_83299 : array_update_83288[9];
  assign array_index_83303 = array_update_72021[add_83300 > 32'h0000_0009 ? 4'h9 : add_83300[3:0]];
  assign array_index_83304 = array_update_83301[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_83308 = smul32b_32b_x_32b(array_index_82832[add_83300 > 32'h0000_0009 ? 4'h9 : add_83300[3:0]], array_index_83303[add_83233 > 32'h0000_0009 ? 4'h9 : add_83233[3:0]]);
  assign add_83310 = array_index_83304[add_83233 > 32'h0000_0009 ? 4'h9 : add_83233[3:0]] + smul_83308;
  assign array_update_83312[0] = add_83233 == 32'h0000_0000 ? add_83310 : array_index_83304[0];
  assign array_update_83312[1] = add_83233 == 32'h0000_0001 ? add_83310 : array_index_83304[1];
  assign array_update_83312[2] = add_83233 == 32'h0000_0002 ? add_83310 : array_index_83304[2];
  assign array_update_83312[3] = add_83233 == 32'h0000_0003 ? add_83310 : array_index_83304[3];
  assign array_update_83312[4] = add_83233 == 32'h0000_0004 ? add_83310 : array_index_83304[4];
  assign array_update_83312[5] = add_83233 == 32'h0000_0005 ? add_83310 : array_index_83304[5];
  assign array_update_83312[6] = add_83233 == 32'h0000_0006 ? add_83310 : array_index_83304[6];
  assign array_update_83312[7] = add_83233 == 32'h0000_0007 ? add_83310 : array_index_83304[7];
  assign array_update_83312[8] = add_83233 == 32'h0000_0008 ? add_83310 : array_index_83304[8];
  assign array_update_83312[9] = add_83233 == 32'h0000_0009 ? add_83310 : array_index_83304[9];
  assign add_83313 = add_83300 + 32'h0000_0001;
  assign array_update_83314[0] = add_82825 == 32'h0000_0000 ? array_update_83312 : array_update_83301[0];
  assign array_update_83314[1] = add_82825 == 32'h0000_0001 ? array_update_83312 : array_update_83301[1];
  assign array_update_83314[2] = add_82825 == 32'h0000_0002 ? array_update_83312 : array_update_83301[2];
  assign array_update_83314[3] = add_82825 == 32'h0000_0003 ? array_update_83312 : array_update_83301[3];
  assign array_update_83314[4] = add_82825 == 32'h0000_0004 ? array_update_83312 : array_update_83301[4];
  assign array_update_83314[5] = add_82825 == 32'h0000_0005 ? array_update_83312 : array_update_83301[5];
  assign array_update_83314[6] = add_82825 == 32'h0000_0006 ? array_update_83312 : array_update_83301[6];
  assign array_update_83314[7] = add_82825 == 32'h0000_0007 ? array_update_83312 : array_update_83301[7];
  assign array_update_83314[8] = add_82825 == 32'h0000_0008 ? array_update_83312 : array_update_83301[8];
  assign array_update_83314[9] = add_82825 == 32'h0000_0009 ? array_update_83312 : array_update_83301[9];
  assign array_index_83316 = array_update_72021[add_83313 > 32'h0000_0009 ? 4'h9 : add_83313[3:0]];
  assign array_index_83317 = array_update_83314[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_83321 = smul32b_32b_x_32b(array_index_82832[add_83313 > 32'h0000_0009 ? 4'h9 : add_83313[3:0]], array_index_83316[add_83233 > 32'h0000_0009 ? 4'h9 : add_83233[3:0]]);
  assign add_83323 = array_index_83317[add_83233 > 32'h0000_0009 ? 4'h9 : add_83233[3:0]] + smul_83321;
  assign array_update_83325[0] = add_83233 == 32'h0000_0000 ? add_83323 : array_index_83317[0];
  assign array_update_83325[1] = add_83233 == 32'h0000_0001 ? add_83323 : array_index_83317[1];
  assign array_update_83325[2] = add_83233 == 32'h0000_0002 ? add_83323 : array_index_83317[2];
  assign array_update_83325[3] = add_83233 == 32'h0000_0003 ? add_83323 : array_index_83317[3];
  assign array_update_83325[4] = add_83233 == 32'h0000_0004 ? add_83323 : array_index_83317[4];
  assign array_update_83325[5] = add_83233 == 32'h0000_0005 ? add_83323 : array_index_83317[5];
  assign array_update_83325[6] = add_83233 == 32'h0000_0006 ? add_83323 : array_index_83317[6];
  assign array_update_83325[7] = add_83233 == 32'h0000_0007 ? add_83323 : array_index_83317[7];
  assign array_update_83325[8] = add_83233 == 32'h0000_0008 ? add_83323 : array_index_83317[8];
  assign array_update_83325[9] = add_83233 == 32'h0000_0009 ? add_83323 : array_index_83317[9];
  assign add_83326 = add_83313 + 32'h0000_0001;
  assign array_update_83327[0] = add_82825 == 32'h0000_0000 ? array_update_83325 : array_update_83314[0];
  assign array_update_83327[1] = add_82825 == 32'h0000_0001 ? array_update_83325 : array_update_83314[1];
  assign array_update_83327[2] = add_82825 == 32'h0000_0002 ? array_update_83325 : array_update_83314[2];
  assign array_update_83327[3] = add_82825 == 32'h0000_0003 ? array_update_83325 : array_update_83314[3];
  assign array_update_83327[4] = add_82825 == 32'h0000_0004 ? array_update_83325 : array_update_83314[4];
  assign array_update_83327[5] = add_82825 == 32'h0000_0005 ? array_update_83325 : array_update_83314[5];
  assign array_update_83327[6] = add_82825 == 32'h0000_0006 ? array_update_83325 : array_update_83314[6];
  assign array_update_83327[7] = add_82825 == 32'h0000_0007 ? array_update_83325 : array_update_83314[7];
  assign array_update_83327[8] = add_82825 == 32'h0000_0008 ? array_update_83325 : array_update_83314[8];
  assign array_update_83327[9] = add_82825 == 32'h0000_0009 ? array_update_83325 : array_update_83314[9];
  assign array_index_83329 = array_update_72021[add_83326 > 32'h0000_0009 ? 4'h9 : add_83326[3:0]];
  assign array_index_83330 = array_update_83327[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_83334 = smul32b_32b_x_32b(array_index_82832[add_83326 > 32'h0000_0009 ? 4'h9 : add_83326[3:0]], array_index_83329[add_83233 > 32'h0000_0009 ? 4'h9 : add_83233[3:0]]);
  assign add_83336 = array_index_83330[add_83233 > 32'h0000_0009 ? 4'h9 : add_83233[3:0]] + smul_83334;
  assign array_update_83338[0] = add_83233 == 32'h0000_0000 ? add_83336 : array_index_83330[0];
  assign array_update_83338[1] = add_83233 == 32'h0000_0001 ? add_83336 : array_index_83330[1];
  assign array_update_83338[2] = add_83233 == 32'h0000_0002 ? add_83336 : array_index_83330[2];
  assign array_update_83338[3] = add_83233 == 32'h0000_0003 ? add_83336 : array_index_83330[3];
  assign array_update_83338[4] = add_83233 == 32'h0000_0004 ? add_83336 : array_index_83330[4];
  assign array_update_83338[5] = add_83233 == 32'h0000_0005 ? add_83336 : array_index_83330[5];
  assign array_update_83338[6] = add_83233 == 32'h0000_0006 ? add_83336 : array_index_83330[6];
  assign array_update_83338[7] = add_83233 == 32'h0000_0007 ? add_83336 : array_index_83330[7];
  assign array_update_83338[8] = add_83233 == 32'h0000_0008 ? add_83336 : array_index_83330[8];
  assign array_update_83338[9] = add_83233 == 32'h0000_0009 ? add_83336 : array_index_83330[9];
  assign add_83339 = add_83326 + 32'h0000_0001;
  assign array_update_83340[0] = add_82825 == 32'h0000_0000 ? array_update_83338 : array_update_83327[0];
  assign array_update_83340[1] = add_82825 == 32'h0000_0001 ? array_update_83338 : array_update_83327[1];
  assign array_update_83340[2] = add_82825 == 32'h0000_0002 ? array_update_83338 : array_update_83327[2];
  assign array_update_83340[3] = add_82825 == 32'h0000_0003 ? array_update_83338 : array_update_83327[3];
  assign array_update_83340[4] = add_82825 == 32'h0000_0004 ? array_update_83338 : array_update_83327[4];
  assign array_update_83340[5] = add_82825 == 32'h0000_0005 ? array_update_83338 : array_update_83327[5];
  assign array_update_83340[6] = add_82825 == 32'h0000_0006 ? array_update_83338 : array_update_83327[6];
  assign array_update_83340[7] = add_82825 == 32'h0000_0007 ? array_update_83338 : array_update_83327[7];
  assign array_update_83340[8] = add_82825 == 32'h0000_0008 ? array_update_83338 : array_update_83327[8];
  assign array_update_83340[9] = add_82825 == 32'h0000_0009 ? array_update_83338 : array_update_83327[9];
  assign array_index_83342 = array_update_72021[add_83339 > 32'h0000_0009 ? 4'h9 : add_83339[3:0]];
  assign array_index_83343 = array_update_83340[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_83347 = smul32b_32b_x_32b(array_index_82832[add_83339 > 32'h0000_0009 ? 4'h9 : add_83339[3:0]], array_index_83342[add_83233 > 32'h0000_0009 ? 4'h9 : add_83233[3:0]]);
  assign add_83349 = array_index_83343[add_83233 > 32'h0000_0009 ? 4'h9 : add_83233[3:0]] + smul_83347;
  assign array_update_83351[0] = add_83233 == 32'h0000_0000 ? add_83349 : array_index_83343[0];
  assign array_update_83351[1] = add_83233 == 32'h0000_0001 ? add_83349 : array_index_83343[1];
  assign array_update_83351[2] = add_83233 == 32'h0000_0002 ? add_83349 : array_index_83343[2];
  assign array_update_83351[3] = add_83233 == 32'h0000_0003 ? add_83349 : array_index_83343[3];
  assign array_update_83351[4] = add_83233 == 32'h0000_0004 ? add_83349 : array_index_83343[4];
  assign array_update_83351[5] = add_83233 == 32'h0000_0005 ? add_83349 : array_index_83343[5];
  assign array_update_83351[6] = add_83233 == 32'h0000_0006 ? add_83349 : array_index_83343[6];
  assign array_update_83351[7] = add_83233 == 32'h0000_0007 ? add_83349 : array_index_83343[7];
  assign array_update_83351[8] = add_83233 == 32'h0000_0008 ? add_83349 : array_index_83343[8];
  assign array_update_83351[9] = add_83233 == 32'h0000_0009 ? add_83349 : array_index_83343[9];
  assign add_83352 = add_83339 + 32'h0000_0001;
  assign array_update_83353[0] = add_82825 == 32'h0000_0000 ? array_update_83351 : array_update_83340[0];
  assign array_update_83353[1] = add_82825 == 32'h0000_0001 ? array_update_83351 : array_update_83340[1];
  assign array_update_83353[2] = add_82825 == 32'h0000_0002 ? array_update_83351 : array_update_83340[2];
  assign array_update_83353[3] = add_82825 == 32'h0000_0003 ? array_update_83351 : array_update_83340[3];
  assign array_update_83353[4] = add_82825 == 32'h0000_0004 ? array_update_83351 : array_update_83340[4];
  assign array_update_83353[5] = add_82825 == 32'h0000_0005 ? array_update_83351 : array_update_83340[5];
  assign array_update_83353[6] = add_82825 == 32'h0000_0006 ? array_update_83351 : array_update_83340[6];
  assign array_update_83353[7] = add_82825 == 32'h0000_0007 ? array_update_83351 : array_update_83340[7];
  assign array_update_83353[8] = add_82825 == 32'h0000_0008 ? array_update_83351 : array_update_83340[8];
  assign array_update_83353[9] = add_82825 == 32'h0000_0009 ? array_update_83351 : array_update_83340[9];
  assign array_index_83355 = array_update_72021[add_83352 > 32'h0000_0009 ? 4'h9 : add_83352[3:0]];
  assign array_index_83356 = array_update_83353[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_83360 = smul32b_32b_x_32b(array_index_82832[add_83352 > 32'h0000_0009 ? 4'h9 : add_83352[3:0]], array_index_83355[add_83233 > 32'h0000_0009 ? 4'h9 : add_83233[3:0]]);
  assign add_83362 = array_index_83356[add_83233 > 32'h0000_0009 ? 4'h9 : add_83233[3:0]] + smul_83360;
  assign array_update_83363[0] = add_83233 == 32'h0000_0000 ? add_83362 : array_index_83356[0];
  assign array_update_83363[1] = add_83233 == 32'h0000_0001 ? add_83362 : array_index_83356[1];
  assign array_update_83363[2] = add_83233 == 32'h0000_0002 ? add_83362 : array_index_83356[2];
  assign array_update_83363[3] = add_83233 == 32'h0000_0003 ? add_83362 : array_index_83356[3];
  assign array_update_83363[4] = add_83233 == 32'h0000_0004 ? add_83362 : array_index_83356[4];
  assign array_update_83363[5] = add_83233 == 32'h0000_0005 ? add_83362 : array_index_83356[5];
  assign array_update_83363[6] = add_83233 == 32'h0000_0006 ? add_83362 : array_index_83356[6];
  assign array_update_83363[7] = add_83233 == 32'h0000_0007 ? add_83362 : array_index_83356[7];
  assign array_update_83363[8] = add_83233 == 32'h0000_0008 ? add_83362 : array_index_83356[8];
  assign array_update_83363[9] = add_83233 == 32'h0000_0009 ? add_83362 : array_index_83356[9];
  assign array_update_83364[0] = add_82825 == 32'h0000_0000 ? array_update_83363 : array_update_83353[0];
  assign array_update_83364[1] = add_82825 == 32'h0000_0001 ? array_update_83363 : array_update_83353[1];
  assign array_update_83364[2] = add_82825 == 32'h0000_0002 ? array_update_83363 : array_update_83353[2];
  assign array_update_83364[3] = add_82825 == 32'h0000_0003 ? array_update_83363 : array_update_83353[3];
  assign array_update_83364[4] = add_82825 == 32'h0000_0004 ? array_update_83363 : array_update_83353[4];
  assign array_update_83364[5] = add_82825 == 32'h0000_0005 ? array_update_83363 : array_update_83353[5];
  assign array_update_83364[6] = add_82825 == 32'h0000_0006 ? array_update_83363 : array_update_83353[6];
  assign array_update_83364[7] = add_82825 == 32'h0000_0007 ? array_update_83363 : array_update_83353[7];
  assign array_update_83364[8] = add_82825 == 32'h0000_0008 ? array_update_83363 : array_update_83353[8];
  assign array_update_83364[9] = add_82825 == 32'h0000_0009 ? array_update_83363 : array_update_83353[9];
  assign array_index_83366 = array_update_83364[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign add_83368 = add_83233 + 32'h0000_0001;
  assign array_update_83369[0] = add_83368 == 32'h0000_0000 ? 32'h0000_0000 : array_index_83366[0];
  assign array_update_83369[1] = add_83368 == 32'h0000_0001 ? 32'h0000_0000 : array_index_83366[1];
  assign array_update_83369[2] = add_83368 == 32'h0000_0002 ? 32'h0000_0000 : array_index_83366[2];
  assign array_update_83369[3] = add_83368 == 32'h0000_0003 ? 32'h0000_0000 : array_index_83366[3];
  assign array_update_83369[4] = add_83368 == 32'h0000_0004 ? 32'h0000_0000 : array_index_83366[4];
  assign array_update_83369[5] = add_83368 == 32'h0000_0005 ? 32'h0000_0000 : array_index_83366[5];
  assign array_update_83369[6] = add_83368 == 32'h0000_0006 ? 32'h0000_0000 : array_index_83366[6];
  assign array_update_83369[7] = add_83368 == 32'h0000_0007 ? 32'h0000_0000 : array_index_83366[7];
  assign array_update_83369[8] = add_83368 == 32'h0000_0008 ? 32'h0000_0000 : array_index_83366[8];
  assign array_update_83369[9] = add_83368 == 32'h0000_0009 ? 32'h0000_0000 : array_index_83366[9];
  assign literal_83370 = 32'h0000_0000;
  assign array_update_83371[0] = add_82825 == 32'h0000_0000 ? array_update_83369 : array_update_83364[0];
  assign array_update_83371[1] = add_82825 == 32'h0000_0001 ? array_update_83369 : array_update_83364[1];
  assign array_update_83371[2] = add_82825 == 32'h0000_0002 ? array_update_83369 : array_update_83364[2];
  assign array_update_83371[3] = add_82825 == 32'h0000_0003 ? array_update_83369 : array_update_83364[3];
  assign array_update_83371[4] = add_82825 == 32'h0000_0004 ? array_update_83369 : array_update_83364[4];
  assign array_update_83371[5] = add_82825 == 32'h0000_0005 ? array_update_83369 : array_update_83364[5];
  assign array_update_83371[6] = add_82825 == 32'h0000_0006 ? array_update_83369 : array_update_83364[6];
  assign array_update_83371[7] = add_82825 == 32'h0000_0007 ? array_update_83369 : array_update_83364[7];
  assign array_update_83371[8] = add_82825 == 32'h0000_0008 ? array_update_83369 : array_update_83364[8];
  assign array_update_83371[9] = add_82825 == 32'h0000_0009 ? array_update_83369 : array_update_83364[9];
  assign array_index_83373 = array_update_72021[literal_83370 > 32'h0000_0009 ? 4'h9 : literal_83370[3:0]];
  assign array_index_83374 = array_update_83371[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_83378 = smul32b_32b_x_32b(array_index_82832[literal_83370 > 32'h0000_0009 ? 4'h9 : literal_83370[3:0]], array_index_83373[add_83368 > 32'h0000_0009 ? 4'h9 : add_83368[3:0]]);
  assign add_83380 = array_index_83374[add_83368 > 32'h0000_0009 ? 4'h9 : add_83368[3:0]] + smul_83378;
  assign array_update_83382[0] = add_83368 == 32'h0000_0000 ? add_83380 : array_index_83374[0];
  assign array_update_83382[1] = add_83368 == 32'h0000_0001 ? add_83380 : array_index_83374[1];
  assign array_update_83382[2] = add_83368 == 32'h0000_0002 ? add_83380 : array_index_83374[2];
  assign array_update_83382[3] = add_83368 == 32'h0000_0003 ? add_83380 : array_index_83374[3];
  assign array_update_83382[4] = add_83368 == 32'h0000_0004 ? add_83380 : array_index_83374[4];
  assign array_update_83382[5] = add_83368 == 32'h0000_0005 ? add_83380 : array_index_83374[5];
  assign array_update_83382[6] = add_83368 == 32'h0000_0006 ? add_83380 : array_index_83374[6];
  assign array_update_83382[7] = add_83368 == 32'h0000_0007 ? add_83380 : array_index_83374[7];
  assign array_update_83382[8] = add_83368 == 32'h0000_0008 ? add_83380 : array_index_83374[8];
  assign array_update_83382[9] = add_83368 == 32'h0000_0009 ? add_83380 : array_index_83374[9];
  assign add_83383 = literal_83370 + 32'h0000_0001;
  assign array_update_83384[0] = add_82825 == 32'h0000_0000 ? array_update_83382 : array_update_83371[0];
  assign array_update_83384[1] = add_82825 == 32'h0000_0001 ? array_update_83382 : array_update_83371[1];
  assign array_update_83384[2] = add_82825 == 32'h0000_0002 ? array_update_83382 : array_update_83371[2];
  assign array_update_83384[3] = add_82825 == 32'h0000_0003 ? array_update_83382 : array_update_83371[3];
  assign array_update_83384[4] = add_82825 == 32'h0000_0004 ? array_update_83382 : array_update_83371[4];
  assign array_update_83384[5] = add_82825 == 32'h0000_0005 ? array_update_83382 : array_update_83371[5];
  assign array_update_83384[6] = add_82825 == 32'h0000_0006 ? array_update_83382 : array_update_83371[6];
  assign array_update_83384[7] = add_82825 == 32'h0000_0007 ? array_update_83382 : array_update_83371[7];
  assign array_update_83384[8] = add_82825 == 32'h0000_0008 ? array_update_83382 : array_update_83371[8];
  assign array_update_83384[9] = add_82825 == 32'h0000_0009 ? array_update_83382 : array_update_83371[9];
  assign array_index_83386 = array_update_72021[add_83383 > 32'h0000_0009 ? 4'h9 : add_83383[3:0]];
  assign array_index_83387 = array_update_83384[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_83391 = smul32b_32b_x_32b(array_index_82832[add_83383 > 32'h0000_0009 ? 4'h9 : add_83383[3:0]], array_index_83386[add_83368 > 32'h0000_0009 ? 4'h9 : add_83368[3:0]]);
  assign add_83393 = array_index_83387[add_83368 > 32'h0000_0009 ? 4'h9 : add_83368[3:0]] + smul_83391;
  assign array_update_83395[0] = add_83368 == 32'h0000_0000 ? add_83393 : array_index_83387[0];
  assign array_update_83395[1] = add_83368 == 32'h0000_0001 ? add_83393 : array_index_83387[1];
  assign array_update_83395[2] = add_83368 == 32'h0000_0002 ? add_83393 : array_index_83387[2];
  assign array_update_83395[3] = add_83368 == 32'h0000_0003 ? add_83393 : array_index_83387[3];
  assign array_update_83395[4] = add_83368 == 32'h0000_0004 ? add_83393 : array_index_83387[4];
  assign array_update_83395[5] = add_83368 == 32'h0000_0005 ? add_83393 : array_index_83387[5];
  assign array_update_83395[6] = add_83368 == 32'h0000_0006 ? add_83393 : array_index_83387[6];
  assign array_update_83395[7] = add_83368 == 32'h0000_0007 ? add_83393 : array_index_83387[7];
  assign array_update_83395[8] = add_83368 == 32'h0000_0008 ? add_83393 : array_index_83387[8];
  assign array_update_83395[9] = add_83368 == 32'h0000_0009 ? add_83393 : array_index_83387[9];
  assign add_83396 = add_83383 + 32'h0000_0001;
  assign array_update_83397[0] = add_82825 == 32'h0000_0000 ? array_update_83395 : array_update_83384[0];
  assign array_update_83397[1] = add_82825 == 32'h0000_0001 ? array_update_83395 : array_update_83384[1];
  assign array_update_83397[2] = add_82825 == 32'h0000_0002 ? array_update_83395 : array_update_83384[2];
  assign array_update_83397[3] = add_82825 == 32'h0000_0003 ? array_update_83395 : array_update_83384[3];
  assign array_update_83397[4] = add_82825 == 32'h0000_0004 ? array_update_83395 : array_update_83384[4];
  assign array_update_83397[5] = add_82825 == 32'h0000_0005 ? array_update_83395 : array_update_83384[5];
  assign array_update_83397[6] = add_82825 == 32'h0000_0006 ? array_update_83395 : array_update_83384[6];
  assign array_update_83397[7] = add_82825 == 32'h0000_0007 ? array_update_83395 : array_update_83384[7];
  assign array_update_83397[8] = add_82825 == 32'h0000_0008 ? array_update_83395 : array_update_83384[8];
  assign array_update_83397[9] = add_82825 == 32'h0000_0009 ? array_update_83395 : array_update_83384[9];
  assign array_index_83399 = array_update_72021[add_83396 > 32'h0000_0009 ? 4'h9 : add_83396[3:0]];
  assign array_index_83400 = array_update_83397[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_83404 = smul32b_32b_x_32b(array_index_82832[add_83396 > 32'h0000_0009 ? 4'h9 : add_83396[3:0]], array_index_83399[add_83368 > 32'h0000_0009 ? 4'h9 : add_83368[3:0]]);
  assign add_83406 = array_index_83400[add_83368 > 32'h0000_0009 ? 4'h9 : add_83368[3:0]] + smul_83404;
  assign array_update_83408[0] = add_83368 == 32'h0000_0000 ? add_83406 : array_index_83400[0];
  assign array_update_83408[1] = add_83368 == 32'h0000_0001 ? add_83406 : array_index_83400[1];
  assign array_update_83408[2] = add_83368 == 32'h0000_0002 ? add_83406 : array_index_83400[2];
  assign array_update_83408[3] = add_83368 == 32'h0000_0003 ? add_83406 : array_index_83400[3];
  assign array_update_83408[4] = add_83368 == 32'h0000_0004 ? add_83406 : array_index_83400[4];
  assign array_update_83408[5] = add_83368 == 32'h0000_0005 ? add_83406 : array_index_83400[5];
  assign array_update_83408[6] = add_83368 == 32'h0000_0006 ? add_83406 : array_index_83400[6];
  assign array_update_83408[7] = add_83368 == 32'h0000_0007 ? add_83406 : array_index_83400[7];
  assign array_update_83408[8] = add_83368 == 32'h0000_0008 ? add_83406 : array_index_83400[8];
  assign array_update_83408[9] = add_83368 == 32'h0000_0009 ? add_83406 : array_index_83400[9];
  assign add_83409 = add_83396 + 32'h0000_0001;
  assign array_update_83410[0] = add_82825 == 32'h0000_0000 ? array_update_83408 : array_update_83397[0];
  assign array_update_83410[1] = add_82825 == 32'h0000_0001 ? array_update_83408 : array_update_83397[1];
  assign array_update_83410[2] = add_82825 == 32'h0000_0002 ? array_update_83408 : array_update_83397[2];
  assign array_update_83410[3] = add_82825 == 32'h0000_0003 ? array_update_83408 : array_update_83397[3];
  assign array_update_83410[4] = add_82825 == 32'h0000_0004 ? array_update_83408 : array_update_83397[4];
  assign array_update_83410[5] = add_82825 == 32'h0000_0005 ? array_update_83408 : array_update_83397[5];
  assign array_update_83410[6] = add_82825 == 32'h0000_0006 ? array_update_83408 : array_update_83397[6];
  assign array_update_83410[7] = add_82825 == 32'h0000_0007 ? array_update_83408 : array_update_83397[7];
  assign array_update_83410[8] = add_82825 == 32'h0000_0008 ? array_update_83408 : array_update_83397[8];
  assign array_update_83410[9] = add_82825 == 32'h0000_0009 ? array_update_83408 : array_update_83397[9];
  assign array_index_83412 = array_update_72021[add_83409 > 32'h0000_0009 ? 4'h9 : add_83409[3:0]];
  assign array_index_83413 = array_update_83410[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_83417 = smul32b_32b_x_32b(array_index_82832[add_83409 > 32'h0000_0009 ? 4'h9 : add_83409[3:0]], array_index_83412[add_83368 > 32'h0000_0009 ? 4'h9 : add_83368[3:0]]);
  assign add_83419 = array_index_83413[add_83368 > 32'h0000_0009 ? 4'h9 : add_83368[3:0]] + smul_83417;
  assign array_update_83421[0] = add_83368 == 32'h0000_0000 ? add_83419 : array_index_83413[0];
  assign array_update_83421[1] = add_83368 == 32'h0000_0001 ? add_83419 : array_index_83413[1];
  assign array_update_83421[2] = add_83368 == 32'h0000_0002 ? add_83419 : array_index_83413[2];
  assign array_update_83421[3] = add_83368 == 32'h0000_0003 ? add_83419 : array_index_83413[3];
  assign array_update_83421[4] = add_83368 == 32'h0000_0004 ? add_83419 : array_index_83413[4];
  assign array_update_83421[5] = add_83368 == 32'h0000_0005 ? add_83419 : array_index_83413[5];
  assign array_update_83421[6] = add_83368 == 32'h0000_0006 ? add_83419 : array_index_83413[6];
  assign array_update_83421[7] = add_83368 == 32'h0000_0007 ? add_83419 : array_index_83413[7];
  assign array_update_83421[8] = add_83368 == 32'h0000_0008 ? add_83419 : array_index_83413[8];
  assign array_update_83421[9] = add_83368 == 32'h0000_0009 ? add_83419 : array_index_83413[9];
  assign add_83422 = add_83409 + 32'h0000_0001;
  assign array_update_83423[0] = add_82825 == 32'h0000_0000 ? array_update_83421 : array_update_83410[0];
  assign array_update_83423[1] = add_82825 == 32'h0000_0001 ? array_update_83421 : array_update_83410[1];
  assign array_update_83423[2] = add_82825 == 32'h0000_0002 ? array_update_83421 : array_update_83410[2];
  assign array_update_83423[3] = add_82825 == 32'h0000_0003 ? array_update_83421 : array_update_83410[3];
  assign array_update_83423[4] = add_82825 == 32'h0000_0004 ? array_update_83421 : array_update_83410[4];
  assign array_update_83423[5] = add_82825 == 32'h0000_0005 ? array_update_83421 : array_update_83410[5];
  assign array_update_83423[6] = add_82825 == 32'h0000_0006 ? array_update_83421 : array_update_83410[6];
  assign array_update_83423[7] = add_82825 == 32'h0000_0007 ? array_update_83421 : array_update_83410[7];
  assign array_update_83423[8] = add_82825 == 32'h0000_0008 ? array_update_83421 : array_update_83410[8];
  assign array_update_83423[9] = add_82825 == 32'h0000_0009 ? array_update_83421 : array_update_83410[9];
  assign array_index_83425 = array_update_72021[add_83422 > 32'h0000_0009 ? 4'h9 : add_83422[3:0]];
  assign array_index_83426 = array_update_83423[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_83430 = smul32b_32b_x_32b(array_index_82832[add_83422 > 32'h0000_0009 ? 4'h9 : add_83422[3:0]], array_index_83425[add_83368 > 32'h0000_0009 ? 4'h9 : add_83368[3:0]]);
  assign add_83432 = array_index_83426[add_83368 > 32'h0000_0009 ? 4'h9 : add_83368[3:0]] + smul_83430;
  assign array_update_83434[0] = add_83368 == 32'h0000_0000 ? add_83432 : array_index_83426[0];
  assign array_update_83434[1] = add_83368 == 32'h0000_0001 ? add_83432 : array_index_83426[1];
  assign array_update_83434[2] = add_83368 == 32'h0000_0002 ? add_83432 : array_index_83426[2];
  assign array_update_83434[3] = add_83368 == 32'h0000_0003 ? add_83432 : array_index_83426[3];
  assign array_update_83434[4] = add_83368 == 32'h0000_0004 ? add_83432 : array_index_83426[4];
  assign array_update_83434[5] = add_83368 == 32'h0000_0005 ? add_83432 : array_index_83426[5];
  assign array_update_83434[6] = add_83368 == 32'h0000_0006 ? add_83432 : array_index_83426[6];
  assign array_update_83434[7] = add_83368 == 32'h0000_0007 ? add_83432 : array_index_83426[7];
  assign array_update_83434[8] = add_83368 == 32'h0000_0008 ? add_83432 : array_index_83426[8];
  assign array_update_83434[9] = add_83368 == 32'h0000_0009 ? add_83432 : array_index_83426[9];
  assign add_83435 = add_83422 + 32'h0000_0001;
  assign array_update_83436[0] = add_82825 == 32'h0000_0000 ? array_update_83434 : array_update_83423[0];
  assign array_update_83436[1] = add_82825 == 32'h0000_0001 ? array_update_83434 : array_update_83423[1];
  assign array_update_83436[2] = add_82825 == 32'h0000_0002 ? array_update_83434 : array_update_83423[2];
  assign array_update_83436[3] = add_82825 == 32'h0000_0003 ? array_update_83434 : array_update_83423[3];
  assign array_update_83436[4] = add_82825 == 32'h0000_0004 ? array_update_83434 : array_update_83423[4];
  assign array_update_83436[5] = add_82825 == 32'h0000_0005 ? array_update_83434 : array_update_83423[5];
  assign array_update_83436[6] = add_82825 == 32'h0000_0006 ? array_update_83434 : array_update_83423[6];
  assign array_update_83436[7] = add_82825 == 32'h0000_0007 ? array_update_83434 : array_update_83423[7];
  assign array_update_83436[8] = add_82825 == 32'h0000_0008 ? array_update_83434 : array_update_83423[8];
  assign array_update_83436[9] = add_82825 == 32'h0000_0009 ? array_update_83434 : array_update_83423[9];
  assign array_index_83438 = array_update_72021[add_83435 > 32'h0000_0009 ? 4'h9 : add_83435[3:0]];
  assign array_index_83439 = array_update_83436[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_83443 = smul32b_32b_x_32b(array_index_82832[add_83435 > 32'h0000_0009 ? 4'h9 : add_83435[3:0]], array_index_83438[add_83368 > 32'h0000_0009 ? 4'h9 : add_83368[3:0]]);
  assign add_83445 = array_index_83439[add_83368 > 32'h0000_0009 ? 4'h9 : add_83368[3:0]] + smul_83443;
  assign array_update_83447[0] = add_83368 == 32'h0000_0000 ? add_83445 : array_index_83439[0];
  assign array_update_83447[1] = add_83368 == 32'h0000_0001 ? add_83445 : array_index_83439[1];
  assign array_update_83447[2] = add_83368 == 32'h0000_0002 ? add_83445 : array_index_83439[2];
  assign array_update_83447[3] = add_83368 == 32'h0000_0003 ? add_83445 : array_index_83439[3];
  assign array_update_83447[4] = add_83368 == 32'h0000_0004 ? add_83445 : array_index_83439[4];
  assign array_update_83447[5] = add_83368 == 32'h0000_0005 ? add_83445 : array_index_83439[5];
  assign array_update_83447[6] = add_83368 == 32'h0000_0006 ? add_83445 : array_index_83439[6];
  assign array_update_83447[7] = add_83368 == 32'h0000_0007 ? add_83445 : array_index_83439[7];
  assign array_update_83447[8] = add_83368 == 32'h0000_0008 ? add_83445 : array_index_83439[8];
  assign array_update_83447[9] = add_83368 == 32'h0000_0009 ? add_83445 : array_index_83439[9];
  assign add_83448 = add_83435 + 32'h0000_0001;
  assign array_update_83449[0] = add_82825 == 32'h0000_0000 ? array_update_83447 : array_update_83436[0];
  assign array_update_83449[1] = add_82825 == 32'h0000_0001 ? array_update_83447 : array_update_83436[1];
  assign array_update_83449[2] = add_82825 == 32'h0000_0002 ? array_update_83447 : array_update_83436[2];
  assign array_update_83449[3] = add_82825 == 32'h0000_0003 ? array_update_83447 : array_update_83436[3];
  assign array_update_83449[4] = add_82825 == 32'h0000_0004 ? array_update_83447 : array_update_83436[4];
  assign array_update_83449[5] = add_82825 == 32'h0000_0005 ? array_update_83447 : array_update_83436[5];
  assign array_update_83449[6] = add_82825 == 32'h0000_0006 ? array_update_83447 : array_update_83436[6];
  assign array_update_83449[7] = add_82825 == 32'h0000_0007 ? array_update_83447 : array_update_83436[7];
  assign array_update_83449[8] = add_82825 == 32'h0000_0008 ? array_update_83447 : array_update_83436[8];
  assign array_update_83449[9] = add_82825 == 32'h0000_0009 ? array_update_83447 : array_update_83436[9];
  assign array_index_83451 = array_update_72021[add_83448 > 32'h0000_0009 ? 4'h9 : add_83448[3:0]];
  assign array_index_83452 = array_update_83449[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_83456 = smul32b_32b_x_32b(array_index_82832[add_83448 > 32'h0000_0009 ? 4'h9 : add_83448[3:0]], array_index_83451[add_83368 > 32'h0000_0009 ? 4'h9 : add_83368[3:0]]);
  assign add_83458 = array_index_83452[add_83368 > 32'h0000_0009 ? 4'h9 : add_83368[3:0]] + smul_83456;
  assign array_update_83460[0] = add_83368 == 32'h0000_0000 ? add_83458 : array_index_83452[0];
  assign array_update_83460[1] = add_83368 == 32'h0000_0001 ? add_83458 : array_index_83452[1];
  assign array_update_83460[2] = add_83368 == 32'h0000_0002 ? add_83458 : array_index_83452[2];
  assign array_update_83460[3] = add_83368 == 32'h0000_0003 ? add_83458 : array_index_83452[3];
  assign array_update_83460[4] = add_83368 == 32'h0000_0004 ? add_83458 : array_index_83452[4];
  assign array_update_83460[5] = add_83368 == 32'h0000_0005 ? add_83458 : array_index_83452[5];
  assign array_update_83460[6] = add_83368 == 32'h0000_0006 ? add_83458 : array_index_83452[6];
  assign array_update_83460[7] = add_83368 == 32'h0000_0007 ? add_83458 : array_index_83452[7];
  assign array_update_83460[8] = add_83368 == 32'h0000_0008 ? add_83458 : array_index_83452[8];
  assign array_update_83460[9] = add_83368 == 32'h0000_0009 ? add_83458 : array_index_83452[9];
  assign add_83461 = add_83448 + 32'h0000_0001;
  assign array_update_83462[0] = add_82825 == 32'h0000_0000 ? array_update_83460 : array_update_83449[0];
  assign array_update_83462[1] = add_82825 == 32'h0000_0001 ? array_update_83460 : array_update_83449[1];
  assign array_update_83462[2] = add_82825 == 32'h0000_0002 ? array_update_83460 : array_update_83449[2];
  assign array_update_83462[3] = add_82825 == 32'h0000_0003 ? array_update_83460 : array_update_83449[3];
  assign array_update_83462[4] = add_82825 == 32'h0000_0004 ? array_update_83460 : array_update_83449[4];
  assign array_update_83462[5] = add_82825 == 32'h0000_0005 ? array_update_83460 : array_update_83449[5];
  assign array_update_83462[6] = add_82825 == 32'h0000_0006 ? array_update_83460 : array_update_83449[6];
  assign array_update_83462[7] = add_82825 == 32'h0000_0007 ? array_update_83460 : array_update_83449[7];
  assign array_update_83462[8] = add_82825 == 32'h0000_0008 ? array_update_83460 : array_update_83449[8];
  assign array_update_83462[9] = add_82825 == 32'h0000_0009 ? array_update_83460 : array_update_83449[9];
  assign array_index_83464 = array_update_72021[add_83461 > 32'h0000_0009 ? 4'h9 : add_83461[3:0]];
  assign array_index_83465 = array_update_83462[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_83469 = smul32b_32b_x_32b(array_index_82832[add_83461 > 32'h0000_0009 ? 4'h9 : add_83461[3:0]], array_index_83464[add_83368 > 32'h0000_0009 ? 4'h9 : add_83368[3:0]]);
  assign add_83471 = array_index_83465[add_83368 > 32'h0000_0009 ? 4'h9 : add_83368[3:0]] + smul_83469;
  assign array_update_83473[0] = add_83368 == 32'h0000_0000 ? add_83471 : array_index_83465[0];
  assign array_update_83473[1] = add_83368 == 32'h0000_0001 ? add_83471 : array_index_83465[1];
  assign array_update_83473[2] = add_83368 == 32'h0000_0002 ? add_83471 : array_index_83465[2];
  assign array_update_83473[3] = add_83368 == 32'h0000_0003 ? add_83471 : array_index_83465[3];
  assign array_update_83473[4] = add_83368 == 32'h0000_0004 ? add_83471 : array_index_83465[4];
  assign array_update_83473[5] = add_83368 == 32'h0000_0005 ? add_83471 : array_index_83465[5];
  assign array_update_83473[6] = add_83368 == 32'h0000_0006 ? add_83471 : array_index_83465[6];
  assign array_update_83473[7] = add_83368 == 32'h0000_0007 ? add_83471 : array_index_83465[7];
  assign array_update_83473[8] = add_83368 == 32'h0000_0008 ? add_83471 : array_index_83465[8];
  assign array_update_83473[9] = add_83368 == 32'h0000_0009 ? add_83471 : array_index_83465[9];
  assign add_83474 = add_83461 + 32'h0000_0001;
  assign array_update_83475[0] = add_82825 == 32'h0000_0000 ? array_update_83473 : array_update_83462[0];
  assign array_update_83475[1] = add_82825 == 32'h0000_0001 ? array_update_83473 : array_update_83462[1];
  assign array_update_83475[2] = add_82825 == 32'h0000_0002 ? array_update_83473 : array_update_83462[2];
  assign array_update_83475[3] = add_82825 == 32'h0000_0003 ? array_update_83473 : array_update_83462[3];
  assign array_update_83475[4] = add_82825 == 32'h0000_0004 ? array_update_83473 : array_update_83462[4];
  assign array_update_83475[5] = add_82825 == 32'h0000_0005 ? array_update_83473 : array_update_83462[5];
  assign array_update_83475[6] = add_82825 == 32'h0000_0006 ? array_update_83473 : array_update_83462[6];
  assign array_update_83475[7] = add_82825 == 32'h0000_0007 ? array_update_83473 : array_update_83462[7];
  assign array_update_83475[8] = add_82825 == 32'h0000_0008 ? array_update_83473 : array_update_83462[8];
  assign array_update_83475[9] = add_82825 == 32'h0000_0009 ? array_update_83473 : array_update_83462[9];
  assign array_index_83477 = array_update_72021[add_83474 > 32'h0000_0009 ? 4'h9 : add_83474[3:0]];
  assign array_index_83478 = array_update_83475[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_83482 = smul32b_32b_x_32b(array_index_82832[add_83474 > 32'h0000_0009 ? 4'h9 : add_83474[3:0]], array_index_83477[add_83368 > 32'h0000_0009 ? 4'h9 : add_83368[3:0]]);
  assign add_83484 = array_index_83478[add_83368 > 32'h0000_0009 ? 4'h9 : add_83368[3:0]] + smul_83482;
  assign array_update_83486[0] = add_83368 == 32'h0000_0000 ? add_83484 : array_index_83478[0];
  assign array_update_83486[1] = add_83368 == 32'h0000_0001 ? add_83484 : array_index_83478[1];
  assign array_update_83486[2] = add_83368 == 32'h0000_0002 ? add_83484 : array_index_83478[2];
  assign array_update_83486[3] = add_83368 == 32'h0000_0003 ? add_83484 : array_index_83478[3];
  assign array_update_83486[4] = add_83368 == 32'h0000_0004 ? add_83484 : array_index_83478[4];
  assign array_update_83486[5] = add_83368 == 32'h0000_0005 ? add_83484 : array_index_83478[5];
  assign array_update_83486[6] = add_83368 == 32'h0000_0006 ? add_83484 : array_index_83478[6];
  assign array_update_83486[7] = add_83368 == 32'h0000_0007 ? add_83484 : array_index_83478[7];
  assign array_update_83486[8] = add_83368 == 32'h0000_0008 ? add_83484 : array_index_83478[8];
  assign array_update_83486[9] = add_83368 == 32'h0000_0009 ? add_83484 : array_index_83478[9];
  assign add_83487 = add_83474 + 32'h0000_0001;
  assign array_update_83488[0] = add_82825 == 32'h0000_0000 ? array_update_83486 : array_update_83475[0];
  assign array_update_83488[1] = add_82825 == 32'h0000_0001 ? array_update_83486 : array_update_83475[1];
  assign array_update_83488[2] = add_82825 == 32'h0000_0002 ? array_update_83486 : array_update_83475[2];
  assign array_update_83488[3] = add_82825 == 32'h0000_0003 ? array_update_83486 : array_update_83475[3];
  assign array_update_83488[4] = add_82825 == 32'h0000_0004 ? array_update_83486 : array_update_83475[4];
  assign array_update_83488[5] = add_82825 == 32'h0000_0005 ? array_update_83486 : array_update_83475[5];
  assign array_update_83488[6] = add_82825 == 32'h0000_0006 ? array_update_83486 : array_update_83475[6];
  assign array_update_83488[7] = add_82825 == 32'h0000_0007 ? array_update_83486 : array_update_83475[7];
  assign array_update_83488[8] = add_82825 == 32'h0000_0008 ? array_update_83486 : array_update_83475[8];
  assign array_update_83488[9] = add_82825 == 32'h0000_0009 ? array_update_83486 : array_update_83475[9];
  assign array_index_83490 = array_update_72021[add_83487 > 32'h0000_0009 ? 4'h9 : add_83487[3:0]];
  assign array_index_83491 = array_update_83488[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_83495 = smul32b_32b_x_32b(array_index_82832[add_83487 > 32'h0000_0009 ? 4'h9 : add_83487[3:0]], array_index_83490[add_83368 > 32'h0000_0009 ? 4'h9 : add_83368[3:0]]);
  assign add_83497 = array_index_83491[add_83368 > 32'h0000_0009 ? 4'h9 : add_83368[3:0]] + smul_83495;
  assign array_update_83498[0] = add_83368 == 32'h0000_0000 ? add_83497 : array_index_83491[0];
  assign array_update_83498[1] = add_83368 == 32'h0000_0001 ? add_83497 : array_index_83491[1];
  assign array_update_83498[2] = add_83368 == 32'h0000_0002 ? add_83497 : array_index_83491[2];
  assign array_update_83498[3] = add_83368 == 32'h0000_0003 ? add_83497 : array_index_83491[3];
  assign array_update_83498[4] = add_83368 == 32'h0000_0004 ? add_83497 : array_index_83491[4];
  assign array_update_83498[5] = add_83368 == 32'h0000_0005 ? add_83497 : array_index_83491[5];
  assign array_update_83498[6] = add_83368 == 32'h0000_0006 ? add_83497 : array_index_83491[6];
  assign array_update_83498[7] = add_83368 == 32'h0000_0007 ? add_83497 : array_index_83491[7];
  assign array_update_83498[8] = add_83368 == 32'h0000_0008 ? add_83497 : array_index_83491[8];
  assign array_update_83498[9] = add_83368 == 32'h0000_0009 ? add_83497 : array_index_83491[9];
  assign array_update_83499[0] = add_82825 == 32'h0000_0000 ? array_update_83498 : array_update_83488[0];
  assign array_update_83499[1] = add_82825 == 32'h0000_0001 ? array_update_83498 : array_update_83488[1];
  assign array_update_83499[2] = add_82825 == 32'h0000_0002 ? array_update_83498 : array_update_83488[2];
  assign array_update_83499[3] = add_82825 == 32'h0000_0003 ? array_update_83498 : array_update_83488[3];
  assign array_update_83499[4] = add_82825 == 32'h0000_0004 ? array_update_83498 : array_update_83488[4];
  assign array_update_83499[5] = add_82825 == 32'h0000_0005 ? array_update_83498 : array_update_83488[5];
  assign array_update_83499[6] = add_82825 == 32'h0000_0006 ? array_update_83498 : array_update_83488[6];
  assign array_update_83499[7] = add_82825 == 32'h0000_0007 ? array_update_83498 : array_update_83488[7];
  assign array_update_83499[8] = add_82825 == 32'h0000_0008 ? array_update_83498 : array_update_83488[8];
  assign array_update_83499[9] = add_82825 == 32'h0000_0009 ? array_update_83498 : array_update_83488[9];
  assign array_index_83501 = array_update_83499[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign add_83503 = add_83368 + 32'h0000_0001;
  assign array_update_83504[0] = add_83503 == 32'h0000_0000 ? 32'h0000_0000 : array_index_83501[0];
  assign array_update_83504[1] = add_83503 == 32'h0000_0001 ? 32'h0000_0000 : array_index_83501[1];
  assign array_update_83504[2] = add_83503 == 32'h0000_0002 ? 32'h0000_0000 : array_index_83501[2];
  assign array_update_83504[3] = add_83503 == 32'h0000_0003 ? 32'h0000_0000 : array_index_83501[3];
  assign array_update_83504[4] = add_83503 == 32'h0000_0004 ? 32'h0000_0000 : array_index_83501[4];
  assign array_update_83504[5] = add_83503 == 32'h0000_0005 ? 32'h0000_0000 : array_index_83501[5];
  assign array_update_83504[6] = add_83503 == 32'h0000_0006 ? 32'h0000_0000 : array_index_83501[6];
  assign array_update_83504[7] = add_83503 == 32'h0000_0007 ? 32'h0000_0000 : array_index_83501[7];
  assign array_update_83504[8] = add_83503 == 32'h0000_0008 ? 32'h0000_0000 : array_index_83501[8];
  assign array_update_83504[9] = add_83503 == 32'h0000_0009 ? 32'h0000_0000 : array_index_83501[9];
  assign literal_83505 = 32'h0000_0000;
  assign array_update_83506[0] = add_82825 == 32'h0000_0000 ? array_update_83504 : array_update_83499[0];
  assign array_update_83506[1] = add_82825 == 32'h0000_0001 ? array_update_83504 : array_update_83499[1];
  assign array_update_83506[2] = add_82825 == 32'h0000_0002 ? array_update_83504 : array_update_83499[2];
  assign array_update_83506[3] = add_82825 == 32'h0000_0003 ? array_update_83504 : array_update_83499[3];
  assign array_update_83506[4] = add_82825 == 32'h0000_0004 ? array_update_83504 : array_update_83499[4];
  assign array_update_83506[5] = add_82825 == 32'h0000_0005 ? array_update_83504 : array_update_83499[5];
  assign array_update_83506[6] = add_82825 == 32'h0000_0006 ? array_update_83504 : array_update_83499[6];
  assign array_update_83506[7] = add_82825 == 32'h0000_0007 ? array_update_83504 : array_update_83499[7];
  assign array_update_83506[8] = add_82825 == 32'h0000_0008 ? array_update_83504 : array_update_83499[8];
  assign array_update_83506[9] = add_82825 == 32'h0000_0009 ? array_update_83504 : array_update_83499[9];
  assign array_index_83508 = array_update_72021[literal_83505 > 32'h0000_0009 ? 4'h9 : literal_83505[3:0]];
  assign array_index_83509 = array_update_83506[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_83513 = smul32b_32b_x_32b(array_index_82832[literal_83505 > 32'h0000_0009 ? 4'h9 : literal_83505[3:0]], array_index_83508[add_83503 > 32'h0000_0009 ? 4'h9 : add_83503[3:0]]);
  assign add_83515 = array_index_83509[add_83503 > 32'h0000_0009 ? 4'h9 : add_83503[3:0]] + smul_83513;
  assign array_update_83517[0] = add_83503 == 32'h0000_0000 ? add_83515 : array_index_83509[0];
  assign array_update_83517[1] = add_83503 == 32'h0000_0001 ? add_83515 : array_index_83509[1];
  assign array_update_83517[2] = add_83503 == 32'h0000_0002 ? add_83515 : array_index_83509[2];
  assign array_update_83517[3] = add_83503 == 32'h0000_0003 ? add_83515 : array_index_83509[3];
  assign array_update_83517[4] = add_83503 == 32'h0000_0004 ? add_83515 : array_index_83509[4];
  assign array_update_83517[5] = add_83503 == 32'h0000_0005 ? add_83515 : array_index_83509[5];
  assign array_update_83517[6] = add_83503 == 32'h0000_0006 ? add_83515 : array_index_83509[6];
  assign array_update_83517[7] = add_83503 == 32'h0000_0007 ? add_83515 : array_index_83509[7];
  assign array_update_83517[8] = add_83503 == 32'h0000_0008 ? add_83515 : array_index_83509[8];
  assign array_update_83517[9] = add_83503 == 32'h0000_0009 ? add_83515 : array_index_83509[9];
  assign add_83518 = literal_83505 + 32'h0000_0001;
  assign array_update_83519[0] = add_82825 == 32'h0000_0000 ? array_update_83517 : array_update_83506[0];
  assign array_update_83519[1] = add_82825 == 32'h0000_0001 ? array_update_83517 : array_update_83506[1];
  assign array_update_83519[2] = add_82825 == 32'h0000_0002 ? array_update_83517 : array_update_83506[2];
  assign array_update_83519[3] = add_82825 == 32'h0000_0003 ? array_update_83517 : array_update_83506[3];
  assign array_update_83519[4] = add_82825 == 32'h0000_0004 ? array_update_83517 : array_update_83506[4];
  assign array_update_83519[5] = add_82825 == 32'h0000_0005 ? array_update_83517 : array_update_83506[5];
  assign array_update_83519[6] = add_82825 == 32'h0000_0006 ? array_update_83517 : array_update_83506[6];
  assign array_update_83519[7] = add_82825 == 32'h0000_0007 ? array_update_83517 : array_update_83506[7];
  assign array_update_83519[8] = add_82825 == 32'h0000_0008 ? array_update_83517 : array_update_83506[8];
  assign array_update_83519[9] = add_82825 == 32'h0000_0009 ? array_update_83517 : array_update_83506[9];
  assign array_index_83521 = array_update_72021[add_83518 > 32'h0000_0009 ? 4'h9 : add_83518[3:0]];
  assign array_index_83522 = array_update_83519[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_83526 = smul32b_32b_x_32b(array_index_82832[add_83518 > 32'h0000_0009 ? 4'h9 : add_83518[3:0]], array_index_83521[add_83503 > 32'h0000_0009 ? 4'h9 : add_83503[3:0]]);
  assign add_83528 = array_index_83522[add_83503 > 32'h0000_0009 ? 4'h9 : add_83503[3:0]] + smul_83526;
  assign array_update_83530[0] = add_83503 == 32'h0000_0000 ? add_83528 : array_index_83522[0];
  assign array_update_83530[1] = add_83503 == 32'h0000_0001 ? add_83528 : array_index_83522[1];
  assign array_update_83530[2] = add_83503 == 32'h0000_0002 ? add_83528 : array_index_83522[2];
  assign array_update_83530[3] = add_83503 == 32'h0000_0003 ? add_83528 : array_index_83522[3];
  assign array_update_83530[4] = add_83503 == 32'h0000_0004 ? add_83528 : array_index_83522[4];
  assign array_update_83530[5] = add_83503 == 32'h0000_0005 ? add_83528 : array_index_83522[5];
  assign array_update_83530[6] = add_83503 == 32'h0000_0006 ? add_83528 : array_index_83522[6];
  assign array_update_83530[7] = add_83503 == 32'h0000_0007 ? add_83528 : array_index_83522[7];
  assign array_update_83530[8] = add_83503 == 32'h0000_0008 ? add_83528 : array_index_83522[8];
  assign array_update_83530[9] = add_83503 == 32'h0000_0009 ? add_83528 : array_index_83522[9];
  assign add_83531 = add_83518 + 32'h0000_0001;
  assign array_update_83532[0] = add_82825 == 32'h0000_0000 ? array_update_83530 : array_update_83519[0];
  assign array_update_83532[1] = add_82825 == 32'h0000_0001 ? array_update_83530 : array_update_83519[1];
  assign array_update_83532[2] = add_82825 == 32'h0000_0002 ? array_update_83530 : array_update_83519[2];
  assign array_update_83532[3] = add_82825 == 32'h0000_0003 ? array_update_83530 : array_update_83519[3];
  assign array_update_83532[4] = add_82825 == 32'h0000_0004 ? array_update_83530 : array_update_83519[4];
  assign array_update_83532[5] = add_82825 == 32'h0000_0005 ? array_update_83530 : array_update_83519[5];
  assign array_update_83532[6] = add_82825 == 32'h0000_0006 ? array_update_83530 : array_update_83519[6];
  assign array_update_83532[7] = add_82825 == 32'h0000_0007 ? array_update_83530 : array_update_83519[7];
  assign array_update_83532[8] = add_82825 == 32'h0000_0008 ? array_update_83530 : array_update_83519[8];
  assign array_update_83532[9] = add_82825 == 32'h0000_0009 ? array_update_83530 : array_update_83519[9];
  assign array_index_83534 = array_update_72021[add_83531 > 32'h0000_0009 ? 4'h9 : add_83531[3:0]];
  assign array_index_83535 = array_update_83532[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_83539 = smul32b_32b_x_32b(array_index_82832[add_83531 > 32'h0000_0009 ? 4'h9 : add_83531[3:0]], array_index_83534[add_83503 > 32'h0000_0009 ? 4'h9 : add_83503[3:0]]);
  assign add_83541 = array_index_83535[add_83503 > 32'h0000_0009 ? 4'h9 : add_83503[3:0]] + smul_83539;
  assign array_update_83543[0] = add_83503 == 32'h0000_0000 ? add_83541 : array_index_83535[0];
  assign array_update_83543[1] = add_83503 == 32'h0000_0001 ? add_83541 : array_index_83535[1];
  assign array_update_83543[2] = add_83503 == 32'h0000_0002 ? add_83541 : array_index_83535[2];
  assign array_update_83543[3] = add_83503 == 32'h0000_0003 ? add_83541 : array_index_83535[3];
  assign array_update_83543[4] = add_83503 == 32'h0000_0004 ? add_83541 : array_index_83535[4];
  assign array_update_83543[5] = add_83503 == 32'h0000_0005 ? add_83541 : array_index_83535[5];
  assign array_update_83543[6] = add_83503 == 32'h0000_0006 ? add_83541 : array_index_83535[6];
  assign array_update_83543[7] = add_83503 == 32'h0000_0007 ? add_83541 : array_index_83535[7];
  assign array_update_83543[8] = add_83503 == 32'h0000_0008 ? add_83541 : array_index_83535[8];
  assign array_update_83543[9] = add_83503 == 32'h0000_0009 ? add_83541 : array_index_83535[9];
  assign add_83544 = add_83531 + 32'h0000_0001;
  assign array_update_83545[0] = add_82825 == 32'h0000_0000 ? array_update_83543 : array_update_83532[0];
  assign array_update_83545[1] = add_82825 == 32'h0000_0001 ? array_update_83543 : array_update_83532[1];
  assign array_update_83545[2] = add_82825 == 32'h0000_0002 ? array_update_83543 : array_update_83532[2];
  assign array_update_83545[3] = add_82825 == 32'h0000_0003 ? array_update_83543 : array_update_83532[3];
  assign array_update_83545[4] = add_82825 == 32'h0000_0004 ? array_update_83543 : array_update_83532[4];
  assign array_update_83545[5] = add_82825 == 32'h0000_0005 ? array_update_83543 : array_update_83532[5];
  assign array_update_83545[6] = add_82825 == 32'h0000_0006 ? array_update_83543 : array_update_83532[6];
  assign array_update_83545[7] = add_82825 == 32'h0000_0007 ? array_update_83543 : array_update_83532[7];
  assign array_update_83545[8] = add_82825 == 32'h0000_0008 ? array_update_83543 : array_update_83532[8];
  assign array_update_83545[9] = add_82825 == 32'h0000_0009 ? array_update_83543 : array_update_83532[9];
  assign array_index_83547 = array_update_72021[add_83544 > 32'h0000_0009 ? 4'h9 : add_83544[3:0]];
  assign array_index_83548 = array_update_83545[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_83552 = smul32b_32b_x_32b(array_index_82832[add_83544 > 32'h0000_0009 ? 4'h9 : add_83544[3:0]], array_index_83547[add_83503 > 32'h0000_0009 ? 4'h9 : add_83503[3:0]]);
  assign add_83554 = array_index_83548[add_83503 > 32'h0000_0009 ? 4'h9 : add_83503[3:0]] + smul_83552;
  assign array_update_83556[0] = add_83503 == 32'h0000_0000 ? add_83554 : array_index_83548[0];
  assign array_update_83556[1] = add_83503 == 32'h0000_0001 ? add_83554 : array_index_83548[1];
  assign array_update_83556[2] = add_83503 == 32'h0000_0002 ? add_83554 : array_index_83548[2];
  assign array_update_83556[3] = add_83503 == 32'h0000_0003 ? add_83554 : array_index_83548[3];
  assign array_update_83556[4] = add_83503 == 32'h0000_0004 ? add_83554 : array_index_83548[4];
  assign array_update_83556[5] = add_83503 == 32'h0000_0005 ? add_83554 : array_index_83548[5];
  assign array_update_83556[6] = add_83503 == 32'h0000_0006 ? add_83554 : array_index_83548[6];
  assign array_update_83556[7] = add_83503 == 32'h0000_0007 ? add_83554 : array_index_83548[7];
  assign array_update_83556[8] = add_83503 == 32'h0000_0008 ? add_83554 : array_index_83548[8];
  assign array_update_83556[9] = add_83503 == 32'h0000_0009 ? add_83554 : array_index_83548[9];
  assign add_83557 = add_83544 + 32'h0000_0001;
  assign array_update_83558[0] = add_82825 == 32'h0000_0000 ? array_update_83556 : array_update_83545[0];
  assign array_update_83558[1] = add_82825 == 32'h0000_0001 ? array_update_83556 : array_update_83545[1];
  assign array_update_83558[2] = add_82825 == 32'h0000_0002 ? array_update_83556 : array_update_83545[2];
  assign array_update_83558[3] = add_82825 == 32'h0000_0003 ? array_update_83556 : array_update_83545[3];
  assign array_update_83558[4] = add_82825 == 32'h0000_0004 ? array_update_83556 : array_update_83545[4];
  assign array_update_83558[5] = add_82825 == 32'h0000_0005 ? array_update_83556 : array_update_83545[5];
  assign array_update_83558[6] = add_82825 == 32'h0000_0006 ? array_update_83556 : array_update_83545[6];
  assign array_update_83558[7] = add_82825 == 32'h0000_0007 ? array_update_83556 : array_update_83545[7];
  assign array_update_83558[8] = add_82825 == 32'h0000_0008 ? array_update_83556 : array_update_83545[8];
  assign array_update_83558[9] = add_82825 == 32'h0000_0009 ? array_update_83556 : array_update_83545[9];
  assign array_index_83560 = array_update_72021[add_83557 > 32'h0000_0009 ? 4'h9 : add_83557[3:0]];
  assign array_index_83561 = array_update_83558[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_83565 = smul32b_32b_x_32b(array_index_82832[add_83557 > 32'h0000_0009 ? 4'h9 : add_83557[3:0]], array_index_83560[add_83503 > 32'h0000_0009 ? 4'h9 : add_83503[3:0]]);
  assign add_83567 = array_index_83561[add_83503 > 32'h0000_0009 ? 4'h9 : add_83503[3:0]] + smul_83565;
  assign array_update_83569[0] = add_83503 == 32'h0000_0000 ? add_83567 : array_index_83561[0];
  assign array_update_83569[1] = add_83503 == 32'h0000_0001 ? add_83567 : array_index_83561[1];
  assign array_update_83569[2] = add_83503 == 32'h0000_0002 ? add_83567 : array_index_83561[2];
  assign array_update_83569[3] = add_83503 == 32'h0000_0003 ? add_83567 : array_index_83561[3];
  assign array_update_83569[4] = add_83503 == 32'h0000_0004 ? add_83567 : array_index_83561[4];
  assign array_update_83569[5] = add_83503 == 32'h0000_0005 ? add_83567 : array_index_83561[5];
  assign array_update_83569[6] = add_83503 == 32'h0000_0006 ? add_83567 : array_index_83561[6];
  assign array_update_83569[7] = add_83503 == 32'h0000_0007 ? add_83567 : array_index_83561[7];
  assign array_update_83569[8] = add_83503 == 32'h0000_0008 ? add_83567 : array_index_83561[8];
  assign array_update_83569[9] = add_83503 == 32'h0000_0009 ? add_83567 : array_index_83561[9];
  assign add_83570 = add_83557 + 32'h0000_0001;
  assign array_update_83571[0] = add_82825 == 32'h0000_0000 ? array_update_83569 : array_update_83558[0];
  assign array_update_83571[1] = add_82825 == 32'h0000_0001 ? array_update_83569 : array_update_83558[1];
  assign array_update_83571[2] = add_82825 == 32'h0000_0002 ? array_update_83569 : array_update_83558[2];
  assign array_update_83571[3] = add_82825 == 32'h0000_0003 ? array_update_83569 : array_update_83558[3];
  assign array_update_83571[4] = add_82825 == 32'h0000_0004 ? array_update_83569 : array_update_83558[4];
  assign array_update_83571[5] = add_82825 == 32'h0000_0005 ? array_update_83569 : array_update_83558[5];
  assign array_update_83571[6] = add_82825 == 32'h0000_0006 ? array_update_83569 : array_update_83558[6];
  assign array_update_83571[7] = add_82825 == 32'h0000_0007 ? array_update_83569 : array_update_83558[7];
  assign array_update_83571[8] = add_82825 == 32'h0000_0008 ? array_update_83569 : array_update_83558[8];
  assign array_update_83571[9] = add_82825 == 32'h0000_0009 ? array_update_83569 : array_update_83558[9];
  assign array_index_83573 = array_update_72021[add_83570 > 32'h0000_0009 ? 4'h9 : add_83570[3:0]];
  assign array_index_83574 = array_update_83571[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_83578 = smul32b_32b_x_32b(array_index_82832[add_83570 > 32'h0000_0009 ? 4'h9 : add_83570[3:0]], array_index_83573[add_83503 > 32'h0000_0009 ? 4'h9 : add_83503[3:0]]);
  assign add_83580 = array_index_83574[add_83503 > 32'h0000_0009 ? 4'h9 : add_83503[3:0]] + smul_83578;
  assign array_update_83582[0] = add_83503 == 32'h0000_0000 ? add_83580 : array_index_83574[0];
  assign array_update_83582[1] = add_83503 == 32'h0000_0001 ? add_83580 : array_index_83574[1];
  assign array_update_83582[2] = add_83503 == 32'h0000_0002 ? add_83580 : array_index_83574[2];
  assign array_update_83582[3] = add_83503 == 32'h0000_0003 ? add_83580 : array_index_83574[3];
  assign array_update_83582[4] = add_83503 == 32'h0000_0004 ? add_83580 : array_index_83574[4];
  assign array_update_83582[5] = add_83503 == 32'h0000_0005 ? add_83580 : array_index_83574[5];
  assign array_update_83582[6] = add_83503 == 32'h0000_0006 ? add_83580 : array_index_83574[6];
  assign array_update_83582[7] = add_83503 == 32'h0000_0007 ? add_83580 : array_index_83574[7];
  assign array_update_83582[8] = add_83503 == 32'h0000_0008 ? add_83580 : array_index_83574[8];
  assign array_update_83582[9] = add_83503 == 32'h0000_0009 ? add_83580 : array_index_83574[9];
  assign add_83583 = add_83570 + 32'h0000_0001;
  assign array_update_83584[0] = add_82825 == 32'h0000_0000 ? array_update_83582 : array_update_83571[0];
  assign array_update_83584[1] = add_82825 == 32'h0000_0001 ? array_update_83582 : array_update_83571[1];
  assign array_update_83584[2] = add_82825 == 32'h0000_0002 ? array_update_83582 : array_update_83571[2];
  assign array_update_83584[3] = add_82825 == 32'h0000_0003 ? array_update_83582 : array_update_83571[3];
  assign array_update_83584[4] = add_82825 == 32'h0000_0004 ? array_update_83582 : array_update_83571[4];
  assign array_update_83584[5] = add_82825 == 32'h0000_0005 ? array_update_83582 : array_update_83571[5];
  assign array_update_83584[6] = add_82825 == 32'h0000_0006 ? array_update_83582 : array_update_83571[6];
  assign array_update_83584[7] = add_82825 == 32'h0000_0007 ? array_update_83582 : array_update_83571[7];
  assign array_update_83584[8] = add_82825 == 32'h0000_0008 ? array_update_83582 : array_update_83571[8];
  assign array_update_83584[9] = add_82825 == 32'h0000_0009 ? array_update_83582 : array_update_83571[9];
  assign array_index_83586 = array_update_72021[add_83583 > 32'h0000_0009 ? 4'h9 : add_83583[3:0]];
  assign array_index_83587 = array_update_83584[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_83591 = smul32b_32b_x_32b(array_index_82832[add_83583 > 32'h0000_0009 ? 4'h9 : add_83583[3:0]], array_index_83586[add_83503 > 32'h0000_0009 ? 4'h9 : add_83503[3:0]]);
  assign add_83593 = array_index_83587[add_83503 > 32'h0000_0009 ? 4'h9 : add_83503[3:0]] + smul_83591;
  assign array_update_83595[0] = add_83503 == 32'h0000_0000 ? add_83593 : array_index_83587[0];
  assign array_update_83595[1] = add_83503 == 32'h0000_0001 ? add_83593 : array_index_83587[1];
  assign array_update_83595[2] = add_83503 == 32'h0000_0002 ? add_83593 : array_index_83587[2];
  assign array_update_83595[3] = add_83503 == 32'h0000_0003 ? add_83593 : array_index_83587[3];
  assign array_update_83595[4] = add_83503 == 32'h0000_0004 ? add_83593 : array_index_83587[4];
  assign array_update_83595[5] = add_83503 == 32'h0000_0005 ? add_83593 : array_index_83587[5];
  assign array_update_83595[6] = add_83503 == 32'h0000_0006 ? add_83593 : array_index_83587[6];
  assign array_update_83595[7] = add_83503 == 32'h0000_0007 ? add_83593 : array_index_83587[7];
  assign array_update_83595[8] = add_83503 == 32'h0000_0008 ? add_83593 : array_index_83587[8];
  assign array_update_83595[9] = add_83503 == 32'h0000_0009 ? add_83593 : array_index_83587[9];
  assign add_83596 = add_83583 + 32'h0000_0001;
  assign array_update_83597[0] = add_82825 == 32'h0000_0000 ? array_update_83595 : array_update_83584[0];
  assign array_update_83597[1] = add_82825 == 32'h0000_0001 ? array_update_83595 : array_update_83584[1];
  assign array_update_83597[2] = add_82825 == 32'h0000_0002 ? array_update_83595 : array_update_83584[2];
  assign array_update_83597[3] = add_82825 == 32'h0000_0003 ? array_update_83595 : array_update_83584[3];
  assign array_update_83597[4] = add_82825 == 32'h0000_0004 ? array_update_83595 : array_update_83584[4];
  assign array_update_83597[5] = add_82825 == 32'h0000_0005 ? array_update_83595 : array_update_83584[5];
  assign array_update_83597[6] = add_82825 == 32'h0000_0006 ? array_update_83595 : array_update_83584[6];
  assign array_update_83597[7] = add_82825 == 32'h0000_0007 ? array_update_83595 : array_update_83584[7];
  assign array_update_83597[8] = add_82825 == 32'h0000_0008 ? array_update_83595 : array_update_83584[8];
  assign array_update_83597[9] = add_82825 == 32'h0000_0009 ? array_update_83595 : array_update_83584[9];
  assign array_index_83599 = array_update_72021[add_83596 > 32'h0000_0009 ? 4'h9 : add_83596[3:0]];
  assign array_index_83600 = array_update_83597[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_83604 = smul32b_32b_x_32b(array_index_82832[add_83596 > 32'h0000_0009 ? 4'h9 : add_83596[3:0]], array_index_83599[add_83503 > 32'h0000_0009 ? 4'h9 : add_83503[3:0]]);
  assign add_83606 = array_index_83600[add_83503 > 32'h0000_0009 ? 4'h9 : add_83503[3:0]] + smul_83604;
  assign array_update_83608[0] = add_83503 == 32'h0000_0000 ? add_83606 : array_index_83600[0];
  assign array_update_83608[1] = add_83503 == 32'h0000_0001 ? add_83606 : array_index_83600[1];
  assign array_update_83608[2] = add_83503 == 32'h0000_0002 ? add_83606 : array_index_83600[2];
  assign array_update_83608[3] = add_83503 == 32'h0000_0003 ? add_83606 : array_index_83600[3];
  assign array_update_83608[4] = add_83503 == 32'h0000_0004 ? add_83606 : array_index_83600[4];
  assign array_update_83608[5] = add_83503 == 32'h0000_0005 ? add_83606 : array_index_83600[5];
  assign array_update_83608[6] = add_83503 == 32'h0000_0006 ? add_83606 : array_index_83600[6];
  assign array_update_83608[7] = add_83503 == 32'h0000_0007 ? add_83606 : array_index_83600[7];
  assign array_update_83608[8] = add_83503 == 32'h0000_0008 ? add_83606 : array_index_83600[8];
  assign array_update_83608[9] = add_83503 == 32'h0000_0009 ? add_83606 : array_index_83600[9];
  assign add_83609 = add_83596 + 32'h0000_0001;
  assign array_update_83610[0] = add_82825 == 32'h0000_0000 ? array_update_83608 : array_update_83597[0];
  assign array_update_83610[1] = add_82825 == 32'h0000_0001 ? array_update_83608 : array_update_83597[1];
  assign array_update_83610[2] = add_82825 == 32'h0000_0002 ? array_update_83608 : array_update_83597[2];
  assign array_update_83610[3] = add_82825 == 32'h0000_0003 ? array_update_83608 : array_update_83597[3];
  assign array_update_83610[4] = add_82825 == 32'h0000_0004 ? array_update_83608 : array_update_83597[4];
  assign array_update_83610[5] = add_82825 == 32'h0000_0005 ? array_update_83608 : array_update_83597[5];
  assign array_update_83610[6] = add_82825 == 32'h0000_0006 ? array_update_83608 : array_update_83597[6];
  assign array_update_83610[7] = add_82825 == 32'h0000_0007 ? array_update_83608 : array_update_83597[7];
  assign array_update_83610[8] = add_82825 == 32'h0000_0008 ? array_update_83608 : array_update_83597[8];
  assign array_update_83610[9] = add_82825 == 32'h0000_0009 ? array_update_83608 : array_update_83597[9];
  assign array_index_83612 = array_update_72021[add_83609 > 32'h0000_0009 ? 4'h9 : add_83609[3:0]];
  assign array_index_83613 = array_update_83610[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_83617 = smul32b_32b_x_32b(array_index_82832[add_83609 > 32'h0000_0009 ? 4'h9 : add_83609[3:0]], array_index_83612[add_83503 > 32'h0000_0009 ? 4'h9 : add_83503[3:0]]);
  assign add_83619 = array_index_83613[add_83503 > 32'h0000_0009 ? 4'h9 : add_83503[3:0]] + smul_83617;
  assign array_update_83621[0] = add_83503 == 32'h0000_0000 ? add_83619 : array_index_83613[0];
  assign array_update_83621[1] = add_83503 == 32'h0000_0001 ? add_83619 : array_index_83613[1];
  assign array_update_83621[2] = add_83503 == 32'h0000_0002 ? add_83619 : array_index_83613[2];
  assign array_update_83621[3] = add_83503 == 32'h0000_0003 ? add_83619 : array_index_83613[3];
  assign array_update_83621[4] = add_83503 == 32'h0000_0004 ? add_83619 : array_index_83613[4];
  assign array_update_83621[5] = add_83503 == 32'h0000_0005 ? add_83619 : array_index_83613[5];
  assign array_update_83621[6] = add_83503 == 32'h0000_0006 ? add_83619 : array_index_83613[6];
  assign array_update_83621[7] = add_83503 == 32'h0000_0007 ? add_83619 : array_index_83613[7];
  assign array_update_83621[8] = add_83503 == 32'h0000_0008 ? add_83619 : array_index_83613[8];
  assign array_update_83621[9] = add_83503 == 32'h0000_0009 ? add_83619 : array_index_83613[9];
  assign add_83622 = add_83609 + 32'h0000_0001;
  assign array_update_83623[0] = add_82825 == 32'h0000_0000 ? array_update_83621 : array_update_83610[0];
  assign array_update_83623[1] = add_82825 == 32'h0000_0001 ? array_update_83621 : array_update_83610[1];
  assign array_update_83623[2] = add_82825 == 32'h0000_0002 ? array_update_83621 : array_update_83610[2];
  assign array_update_83623[3] = add_82825 == 32'h0000_0003 ? array_update_83621 : array_update_83610[3];
  assign array_update_83623[4] = add_82825 == 32'h0000_0004 ? array_update_83621 : array_update_83610[4];
  assign array_update_83623[5] = add_82825 == 32'h0000_0005 ? array_update_83621 : array_update_83610[5];
  assign array_update_83623[6] = add_82825 == 32'h0000_0006 ? array_update_83621 : array_update_83610[6];
  assign array_update_83623[7] = add_82825 == 32'h0000_0007 ? array_update_83621 : array_update_83610[7];
  assign array_update_83623[8] = add_82825 == 32'h0000_0008 ? array_update_83621 : array_update_83610[8];
  assign array_update_83623[9] = add_82825 == 32'h0000_0009 ? array_update_83621 : array_update_83610[9];
  assign array_index_83625 = array_update_72021[add_83622 > 32'h0000_0009 ? 4'h9 : add_83622[3:0]];
  assign array_index_83626 = array_update_83623[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_83630 = smul32b_32b_x_32b(array_index_82832[add_83622 > 32'h0000_0009 ? 4'h9 : add_83622[3:0]], array_index_83625[add_83503 > 32'h0000_0009 ? 4'h9 : add_83503[3:0]]);
  assign add_83632 = array_index_83626[add_83503 > 32'h0000_0009 ? 4'h9 : add_83503[3:0]] + smul_83630;
  assign array_update_83633[0] = add_83503 == 32'h0000_0000 ? add_83632 : array_index_83626[0];
  assign array_update_83633[1] = add_83503 == 32'h0000_0001 ? add_83632 : array_index_83626[1];
  assign array_update_83633[2] = add_83503 == 32'h0000_0002 ? add_83632 : array_index_83626[2];
  assign array_update_83633[3] = add_83503 == 32'h0000_0003 ? add_83632 : array_index_83626[3];
  assign array_update_83633[4] = add_83503 == 32'h0000_0004 ? add_83632 : array_index_83626[4];
  assign array_update_83633[5] = add_83503 == 32'h0000_0005 ? add_83632 : array_index_83626[5];
  assign array_update_83633[6] = add_83503 == 32'h0000_0006 ? add_83632 : array_index_83626[6];
  assign array_update_83633[7] = add_83503 == 32'h0000_0007 ? add_83632 : array_index_83626[7];
  assign array_update_83633[8] = add_83503 == 32'h0000_0008 ? add_83632 : array_index_83626[8];
  assign array_update_83633[9] = add_83503 == 32'h0000_0009 ? add_83632 : array_index_83626[9];
  assign array_update_83634[0] = add_82825 == 32'h0000_0000 ? array_update_83633 : array_update_83623[0];
  assign array_update_83634[1] = add_82825 == 32'h0000_0001 ? array_update_83633 : array_update_83623[1];
  assign array_update_83634[2] = add_82825 == 32'h0000_0002 ? array_update_83633 : array_update_83623[2];
  assign array_update_83634[3] = add_82825 == 32'h0000_0003 ? array_update_83633 : array_update_83623[3];
  assign array_update_83634[4] = add_82825 == 32'h0000_0004 ? array_update_83633 : array_update_83623[4];
  assign array_update_83634[5] = add_82825 == 32'h0000_0005 ? array_update_83633 : array_update_83623[5];
  assign array_update_83634[6] = add_82825 == 32'h0000_0006 ? array_update_83633 : array_update_83623[6];
  assign array_update_83634[7] = add_82825 == 32'h0000_0007 ? array_update_83633 : array_update_83623[7];
  assign array_update_83634[8] = add_82825 == 32'h0000_0008 ? array_update_83633 : array_update_83623[8];
  assign array_update_83634[9] = add_82825 == 32'h0000_0009 ? array_update_83633 : array_update_83623[9];
  assign array_index_83636 = array_update_83634[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign add_83638 = add_83503 + 32'h0000_0001;
  assign array_update_83639[0] = add_83638 == 32'h0000_0000 ? 32'h0000_0000 : array_index_83636[0];
  assign array_update_83639[1] = add_83638 == 32'h0000_0001 ? 32'h0000_0000 : array_index_83636[1];
  assign array_update_83639[2] = add_83638 == 32'h0000_0002 ? 32'h0000_0000 : array_index_83636[2];
  assign array_update_83639[3] = add_83638 == 32'h0000_0003 ? 32'h0000_0000 : array_index_83636[3];
  assign array_update_83639[4] = add_83638 == 32'h0000_0004 ? 32'h0000_0000 : array_index_83636[4];
  assign array_update_83639[5] = add_83638 == 32'h0000_0005 ? 32'h0000_0000 : array_index_83636[5];
  assign array_update_83639[6] = add_83638 == 32'h0000_0006 ? 32'h0000_0000 : array_index_83636[6];
  assign array_update_83639[7] = add_83638 == 32'h0000_0007 ? 32'h0000_0000 : array_index_83636[7];
  assign array_update_83639[8] = add_83638 == 32'h0000_0008 ? 32'h0000_0000 : array_index_83636[8];
  assign array_update_83639[9] = add_83638 == 32'h0000_0009 ? 32'h0000_0000 : array_index_83636[9];
  assign literal_83640 = 32'h0000_0000;
  assign array_update_83641[0] = add_82825 == 32'h0000_0000 ? array_update_83639 : array_update_83634[0];
  assign array_update_83641[1] = add_82825 == 32'h0000_0001 ? array_update_83639 : array_update_83634[1];
  assign array_update_83641[2] = add_82825 == 32'h0000_0002 ? array_update_83639 : array_update_83634[2];
  assign array_update_83641[3] = add_82825 == 32'h0000_0003 ? array_update_83639 : array_update_83634[3];
  assign array_update_83641[4] = add_82825 == 32'h0000_0004 ? array_update_83639 : array_update_83634[4];
  assign array_update_83641[5] = add_82825 == 32'h0000_0005 ? array_update_83639 : array_update_83634[5];
  assign array_update_83641[6] = add_82825 == 32'h0000_0006 ? array_update_83639 : array_update_83634[6];
  assign array_update_83641[7] = add_82825 == 32'h0000_0007 ? array_update_83639 : array_update_83634[7];
  assign array_update_83641[8] = add_82825 == 32'h0000_0008 ? array_update_83639 : array_update_83634[8];
  assign array_update_83641[9] = add_82825 == 32'h0000_0009 ? array_update_83639 : array_update_83634[9];
  assign array_index_83643 = array_update_72021[literal_83640 > 32'h0000_0009 ? 4'h9 : literal_83640[3:0]];
  assign array_index_83644 = array_update_83641[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_83648 = smul32b_32b_x_32b(array_index_82832[literal_83640 > 32'h0000_0009 ? 4'h9 : literal_83640[3:0]], array_index_83643[add_83638 > 32'h0000_0009 ? 4'h9 : add_83638[3:0]]);
  assign add_83650 = array_index_83644[add_83638 > 32'h0000_0009 ? 4'h9 : add_83638[3:0]] + smul_83648;
  assign array_update_83652[0] = add_83638 == 32'h0000_0000 ? add_83650 : array_index_83644[0];
  assign array_update_83652[1] = add_83638 == 32'h0000_0001 ? add_83650 : array_index_83644[1];
  assign array_update_83652[2] = add_83638 == 32'h0000_0002 ? add_83650 : array_index_83644[2];
  assign array_update_83652[3] = add_83638 == 32'h0000_0003 ? add_83650 : array_index_83644[3];
  assign array_update_83652[4] = add_83638 == 32'h0000_0004 ? add_83650 : array_index_83644[4];
  assign array_update_83652[5] = add_83638 == 32'h0000_0005 ? add_83650 : array_index_83644[5];
  assign array_update_83652[6] = add_83638 == 32'h0000_0006 ? add_83650 : array_index_83644[6];
  assign array_update_83652[7] = add_83638 == 32'h0000_0007 ? add_83650 : array_index_83644[7];
  assign array_update_83652[8] = add_83638 == 32'h0000_0008 ? add_83650 : array_index_83644[8];
  assign array_update_83652[9] = add_83638 == 32'h0000_0009 ? add_83650 : array_index_83644[9];
  assign add_83653 = literal_83640 + 32'h0000_0001;
  assign array_update_83654[0] = add_82825 == 32'h0000_0000 ? array_update_83652 : array_update_83641[0];
  assign array_update_83654[1] = add_82825 == 32'h0000_0001 ? array_update_83652 : array_update_83641[1];
  assign array_update_83654[2] = add_82825 == 32'h0000_0002 ? array_update_83652 : array_update_83641[2];
  assign array_update_83654[3] = add_82825 == 32'h0000_0003 ? array_update_83652 : array_update_83641[3];
  assign array_update_83654[4] = add_82825 == 32'h0000_0004 ? array_update_83652 : array_update_83641[4];
  assign array_update_83654[5] = add_82825 == 32'h0000_0005 ? array_update_83652 : array_update_83641[5];
  assign array_update_83654[6] = add_82825 == 32'h0000_0006 ? array_update_83652 : array_update_83641[6];
  assign array_update_83654[7] = add_82825 == 32'h0000_0007 ? array_update_83652 : array_update_83641[7];
  assign array_update_83654[8] = add_82825 == 32'h0000_0008 ? array_update_83652 : array_update_83641[8];
  assign array_update_83654[9] = add_82825 == 32'h0000_0009 ? array_update_83652 : array_update_83641[9];
  assign array_index_83656 = array_update_72021[add_83653 > 32'h0000_0009 ? 4'h9 : add_83653[3:0]];
  assign array_index_83657 = array_update_83654[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_83661 = smul32b_32b_x_32b(array_index_82832[add_83653 > 32'h0000_0009 ? 4'h9 : add_83653[3:0]], array_index_83656[add_83638 > 32'h0000_0009 ? 4'h9 : add_83638[3:0]]);
  assign add_83663 = array_index_83657[add_83638 > 32'h0000_0009 ? 4'h9 : add_83638[3:0]] + smul_83661;
  assign array_update_83665[0] = add_83638 == 32'h0000_0000 ? add_83663 : array_index_83657[0];
  assign array_update_83665[1] = add_83638 == 32'h0000_0001 ? add_83663 : array_index_83657[1];
  assign array_update_83665[2] = add_83638 == 32'h0000_0002 ? add_83663 : array_index_83657[2];
  assign array_update_83665[3] = add_83638 == 32'h0000_0003 ? add_83663 : array_index_83657[3];
  assign array_update_83665[4] = add_83638 == 32'h0000_0004 ? add_83663 : array_index_83657[4];
  assign array_update_83665[5] = add_83638 == 32'h0000_0005 ? add_83663 : array_index_83657[5];
  assign array_update_83665[6] = add_83638 == 32'h0000_0006 ? add_83663 : array_index_83657[6];
  assign array_update_83665[7] = add_83638 == 32'h0000_0007 ? add_83663 : array_index_83657[7];
  assign array_update_83665[8] = add_83638 == 32'h0000_0008 ? add_83663 : array_index_83657[8];
  assign array_update_83665[9] = add_83638 == 32'h0000_0009 ? add_83663 : array_index_83657[9];
  assign add_83666 = add_83653 + 32'h0000_0001;
  assign array_update_83667[0] = add_82825 == 32'h0000_0000 ? array_update_83665 : array_update_83654[0];
  assign array_update_83667[1] = add_82825 == 32'h0000_0001 ? array_update_83665 : array_update_83654[1];
  assign array_update_83667[2] = add_82825 == 32'h0000_0002 ? array_update_83665 : array_update_83654[2];
  assign array_update_83667[3] = add_82825 == 32'h0000_0003 ? array_update_83665 : array_update_83654[3];
  assign array_update_83667[4] = add_82825 == 32'h0000_0004 ? array_update_83665 : array_update_83654[4];
  assign array_update_83667[5] = add_82825 == 32'h0000_0005 ? array_update_83665 : array_update_83654[5];
  assign array_update_83667[6] = add_82825 == 32'h0000_0006 ? array_update_83665 : array_update_83654[6];
  assign array_update_83667[7] = add_82825 == 32'h0000_0007 ? array_update_83665 : array_update_83654[7];
  assign array_update_83667[8] = add_82825 == 32'h0000_0008 ? array_update_83665 : array_update_83654[8];
  assign array_update_83667[9] = add_82825 == 32'h0000_0009 ? array_update_83665 : array_update_83654[9];
  assign array_index_83669 = array_update_72021[add_83666 > 32'h0000_0009 ? 4'h9 : add_83666[3:0]];
  assign array_index_83670 = array_update_83667[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_83674 = smul32b_32b_x_32b(array_index_82832[add_83666 > 32'h0000_0009 ? 4'h9 : add_83666[3:0]], array_index_83669[add_83638 > 32'h0000_0009 ? 4'h9 : add_83638[3:0]]);
  assign add_83676 = array_index_83670[add_83638 > 32'h0000_0009 ? 4'h9 : add_83638[3:0]] + smul_83674;
  assign array_update_83678[0] = add_83638 == 32'h0000_0000 ? add_83676 : array_index_83670[0];
  assign array_update_83678[1] = add_83638 == 32'h0000_0001 ? add_83676 : array_index_83670[1];
  assign array_update_83678[2] = add_83638 == 32'h0000_0002 ? add_83676 : array_index_83670[2];
  assign array_update_83678[3] = add_83638 == 32'h0000_0003 ? add_83676 : array_index_83670[3];
  assign array_update_83678[4] = add_83638 == 32'h0000_0004 ? add_83676 : array_index_83670[4];
  assign array_update_83678[5] = add_83638 == 32'h0000_0005 ? add_83676 : array_index_83670[5];
  assign array_update_83678[6] = add_83638 == 32'h0000_0006 ? add_83676 : array_index_83670[6];
  assign array_update_83678[7] = add_83638 == 32'h0000_0007 ? add_83676 : array_index_83670[7];
  assign array_update_83678[8] = add_83638 == 32'h0000_0008 ? add_83676 : array_index_83670[8];
  assign array_update_83678[9] = add_83638 == 32'h0000_0009 ? add_83676 : array_index_83670[9];
  assign add_83679 = add_83666 + 32'h0000_0001;
  assign array_update_83680[0] = add_82825 == 32'h0000_0000 ? array_update_83678 : array_update_83667[0];
  assign array_update_83680[1] = add_82825 == 32'h0000_0001 ? array_update_83678 : array_update_83667[1];
  assign array_update_83680[2] = add_82825 == 32'h0000_0002 ? array_update_83678 : array_update_83667[2];
  assign array_update_83680[3] = add_82825 == 32'h0000_0003 ? array_update_83678 : array_update_83667[3];
  assign array_update_83680[4] = add_82825 == 32'h0000_0004 ? array_update_83678 : array_update_83667[4];
  assign array_update_83680[5] = add_82825 == 32'h0000_0005 ? array_update_83678 : array_update_83667[5];
  assign array_update_83680[6] = add_82825 == 32'h0000_0006 ? array_update_83678 : array_update_83667[6];
  assign array_update_83680[7] = add_82825 == 32'h0000_0007 ? array_update_83678 : array_update_83667[7];
  assign array_update_83680[8] = add_82825 == 32'h0000_0008 ? array_update_83678 : array_update_83667[8];
  assign array_update_83680[9] = add_82825 == 32'h0000_0009 ? array_update_83678 : array_update_83667[9];
  assign array_index_83682 = array_update_72021[add_83679 > 32'h0000_0009 ? 4'h9 : add_83679[3:0]];
  assign array_index_83683 = array_update_83680[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_83687 = smul32b_32b_x_32b(array_index_82832[add_83679 > 32'h0000_0009 ? 4'h9 : add_83679[3:0]], array_index_83682[add_83638 > 32'h0000_0009 ? 4'h9 : add_83638[3:0]]);
  assign add_83689 = array_index_83683[add_83638 > 32'h0000_0009 ? 4'h9 : add_83638[3:0]] + smul_83687;
  assign array_update_83691[0] = add_83638 == 32'h0000_0000 ? add_83689 : array_index_83683[0];
  assign array_update_83691[1] = add_83638 == 32'h0000_0001 ? add_83689 : array_index_83683[1];
  assign array_update_83691[2] = add_83638 == 32'h0000_0002 ? add_83689 : array_index_83683[2];
  assign array_update_83691[3] = add_83638 == 32'h0000_0003 ? add_83689 : array_index_83683[3];
  assign array_update_83691[4] = add_83638 == 32'h0000_0004 ? add_83689 : array_index_83683[4];
  assign array_update_83691[5] = add_83638 == 32'h0000_0005 ? add_83689 : array_index_83683[5];
  assign array_update_83691[6] = add_83638 == 32'h0000_0006 ? add_83689 : array_index_83683[6];
  assign array_update_83691[7] = add_83638 == 32'h0000_0007 ? add_83689 : array_index_83683[7];
  assign array_update_83691[8] = add_83638 == 32'h0000_0008 ? add_83689 : array_index_83683[8];
  assign array_update_83691[9] = add_83638 == 32'h0000_0009 ? add_83689 : array_index_83683[9];
  assign add_83692 = add_83679 + 32'h0000_0001;
  assign array_update_83693[0] = add_82825 == 32'h0000_0000 ? array_update_83691 : array_update_83680[0];
  assign array_update_83693[1] = add_82825 == 32'h0000_0001 ? array_update_83691 : array_update_83680[1];
  assign array_update_83693[2] = add_82825 == 32'h0000_0002 ? array_update_83691 : array_update_83680[2];
  assign array_update_83693[3] = add_82825 == 32'h0000_0003 ? array_update_83691 : array_update_83680[3];
  assign array_update_83693[4] = add_82825 == 32'h0000_0004 ? array_update_83691 : array_update_83680[4];
  assign array_update_83693[5] = add_82825 == 32'h0000_0005 ? array_update_83691 : array_update_83680[5];
  assign array_update_83693[6] = add_82825 == 32'h0000_0006 ? array_update_83691 : array_update_83680[6];
  assign array_update_83693[7] = add_82825 == 32'h0000_0007 ? array_update_83691 : array_update_83680[7];
  assign array_update_83693[8] = add_82825 == 32'h0000_0008 ? array_update_83691 : array_update_83680[8];
  assign array_update_83693[9] = add_82825 == 32'h0000_0009 ? array_update_83691 : array_update_83680[9];
  assign array_index_83695 = array_update_72021[add_83692 > 32'h0000_0009 ? 4'h9 : add_83692[3:0]];
  assign array_index_83696 = array_update_83693[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_83700 = smul32b_32b_x_32b(array_index_82832[add_83692 > 32'h0000_0009 ? 4'h9 : add_83692[3:0]], array_index_83695[add_83638 > 32'h0000_0009 ? 4'h9 : add_83638[3:0]]);
  assign add_83702 = array_index_83696[add_83638 > 32'h0000_0009 ? 4'h9 : add_83638[3:0]] + smul_83700;
  assign array_update_83704[0] = add_83638 == 32'h0000_0000 ? add_83702 : array_index_83696[0];
  assign array_update_83704[1] = add_83638 == 32'h0000_0001 ? add_83702 : array_index_83696[1];
  assign array_update_83704[2] = add_83638 == 32'h0000_0002 ? add_83702 : array_index_83696[2];
  assign array_update_83704[3] = add_83638 == 32'h0000_0003 ? add_83702 : array_index_83696[3];
  assign array_update_83704[4] = add_83638 == 32'h0000_0004 ? add_83702 : array_index_83696[4];
  assign array_update_83704[5] = add_83638 == 32'h0000_0005 ? add_83702 : array_index_83696[5];
  assign array_update_83704[6] = add_83638 == 32'h0000_0006 ? add_83702 : array_index_83696[6];
  assign array_update_83704[7] = add_83638 == 32'h0000_0007 ? add_83702 : array_index_83696[7];
  assign array_update_83704[8] = add_83638 == 32'h0000_0008 ? add_83702 : array_index_83696[8];
  assign array_update_83704[9] = add_83638 == 32'h0000_0009 ? add_83702 : array_index_83696[9];
  assign add_83705 = add_83692 + 32'h0000_0001;
  assign array_update_83706[0] = add_82825 == 32'h0000_0000 ? array_update_83704 : array_update_83693[0];
  assign array_update_83706[1] = add_82825 == 32'h0000_0001 ? array_update_83704 : array_update_83693[1];
  assign array_update_83706[2] = add_82825 == 32'h0000_0002 ? array_update_83704 : array_update_83693[2];
  assign array_update_83706[3] = add_82825 == 32'h0000_0003 ? array_update_83704 : array_update_83693[3];
  assign array_update_83706[4] = add_82825 == 32'h0000_0004 ? array_update_83704 : array_update_83693[4];
  assign array_update_83706[5] = add_82825 == 32'h0000_0005 ? array_update_83704 : array_update_83693[5];
  assign array_update_83706[6] = add_82825 == 32'h0000_0006 ? array_update_83704 : array_update_83693[6];
  assign array_update_83706[7] = add_82825 == 32'h0000_0007 ? array_update_83704 : array_update_83693[7];
  assign array_update_83706[8] = add_82825 == 32'h0000_0008 ? array_update_83704 : array_update_83693[8];
  assign array_update_83706[9] = add_82825 == 32'h0000_0009 ? array_update_83704 : array_update_83693[9];
  assign array_index_83708 = array_update_72021[add_83705 > 32'h0000_0009 ? 4'h9 : add_83705[3:0]];
  assign array_index_83709 = array_update_83706[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_83713 = smul32b_32b_x_32b(array_index_82832[add_83705 > 32'h0000_0009 ? 4'h9 : add_83705[3:0]], array_index_83708[add_83638 > 32'h0000_0009 ? 4'h9 : add_83638[3:0]]);
  assign add_83715 = array_index_83709[add_83638 > 32'h0000_0009 ? 4'h9 : add_83638[3:0]] + smul_83713;
  assign array_update_83717[0] = add_83638 == 32'h0000_0000 ? add_83715 : array_index_83709[0];
  assign array_update_83717[1] = add_83638 == 32'h0000_0001 ? add_83715 : array_index_83709[1];
  assign array_update_83717[2] = add_83638 == 32'h0000_0002 ? add_83715 : array_index_83709[2];
  assign array_update_83717[3] = add_83638 == 32'h0000_0003 ? add_83715 : array_index_83709[3];
  assign array_update_83717[4] = add_83638 == 32'h0000_0004 ? add_83715 : array_index_83709[4];
  assign array_update_83717[5] = add_83638 == 32'h0000_0005 ? add_83715 : array_index_83709[5];
  assign array_update_83717[6] = add_83638 == 32'h0000_0006 ? add_83715 : array_index_83709[6];
  assign array_update_83717[7] = add_83638 == 32'h0000_0007 ? add_83715 : array_index_83709[7];
  assign array_update_83717[8] = add_83638 == 32'h0000_0008 ? add_83715 : array_index_83709[8];
  assign array_update_83717[9] = add_83638 == 32'h0000_0009 ? add_83715 : array_index_83709[9];
  assign add_83718 = add_83705 + 32'h0000_0001;
  assign array_update_83719[0] = add_82825 == 32'h0000_0000 ? array_update_83717 : array_update_83706[0];
  assign array_update_83719[1] = add_82825 == 32'h0000_0001 ? array_update_83717 : array_update_83706[1];
  assign array_update_83719[2] = add_82825 == 32'h0000_0002 ? array_update_83717 : array_update_83706[2];
  assign array_update_83719[3] = add_82825 == 32'h0000_0003 ? array_update_83717 : array_update_83706[3];
  assign array_update_83719[4] = add_82825 == 32'h0000_0004 ? array_update_83717 : array_update_83706[4];
  assign array_update_83719[5] = add_82825 == 32'h0000_0005 ? array_update_83717 : array_update_83706[5];
  assign array_update_83719[6] = add_82825 == 32'h0000_0006 ? array_update_83717 : array_update_83706[6];
  assign array_update_83719[7] = add_82825 == 32'h0000_0007 ? array_update_83717 : array_update_83706[7];
  assign array_update_83719[8] = add_82825 == 32'h0000_0008 ? array_update_83717 : array_update_83706[8];
  assign array_update_83719[9] = add_82825 == 32'h0000_0009 ? array_update_83717 : array_update_83706[9];
  assign array_index_83721 = array_update_72021[add_83718 > 32'h0000_0009 ? 4'h9 : add_83718[3:0]];
  assign array_index_83722 = array_update_83719[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_83726 = smul32b_32b_x_32b(array_index_82832[add_83718 > 32'h0000_0009 ? 4'h9 : add_83718[3:0]], array_index_83721[add_83638 > 32'h0000_0009 ? 4'h9 : add_83638[3:0]]);
  assign add_83728 = array_index_83722[add_83638 > 32'h0000_0009 ? 4'h9 : add_83638[3:0]] + smul_83726;
  assign array_update_83730[0] = add_83638 == 32'h0000_0000 ? add_83728 : array_index_83722[0];
  assign array_update_83730[1] = add_83638 == 32'h0000_0001 ? add_83728 : array_index_83722[1];
  assign array_update_83730[2] = add_83638 == 32'h0000_0002 ? add_83728 : array_index_83722[2];
  assign array_update_83730[3] = add_83638 == 32'h0000_0003 ? add_83728 : array_index_83722[3];
  assign array_update_83730[4] = add_83638 == 32'h0000_0004 ? add_83728 : array_index_83722[4];
  assign array_update_83730[5] = add_83638 == 32'h0000_0005 ? add_83728 : array_index_83722[5];
  assign array_update_83730[6] = add_83638 == 32'h0000_0006 ? add_83728 : array_index_83722[6];
  assign array_update_83730[7] = add_83638 == 32'h0000_0007 ? add_83728 : array_index_83722[7];
  assign array_update_83730[8] = add_83638 == 32'h0000_0008 ? add_83728 : array_index_83722[8];
  assign array_update_83730[9] = add_83638 == 32'h0000_0009 ? add_83728 : array_index_83722[9];
  assign add_83731 = add_83718 + 32'h0000_0001;
  assign array_update_83732[0] = add_82825 == 32'h0000_0000 ? array_update_83730 : array_update_83719[0];
  assign array_update_83732[1] = add_82825 == 32'h0000_0001 ? array_update_83730 : array_update_83719[1];
  assign array_update_83732[2] = add_82825 == 32'h0000_0002 ? array_update_83730 : array_update_83719[2];
  assign array_update_83732[3] = add_82825 == 32'h0000_0003 ? array_update_83730 : array_update_83719[3];
  assign array_update_83732[4] = add_82825 == 32'h0000_0004 ? array_update_83730 : array_update_83719[4];
  assign array_update_83732[5] = add_82825 == 32'h0000_0005 ? array_update_83730 : array_update_83719[5];
  assign array_update_83732[6] = add_82825 == 32'h0000_0006 ? array_update_83730 : array_update_83719[6];
  assign array_update_83732[7] = add_82825 == 32'h0000_0007 ? array_update_83730 : array_update_83719[7];
  assign array_update_83732[8] = add_82825 == 32'h0000_0008 ? array_update_83730 : array_update_83719[8];
  assign array_update_83732[9] = add_82825 == 32'h0000_0009 ? array_update_83730 : array_update_83719[9];
  assign array_index_83734 = array_update_72021[add_83731 > 32'h0000_0009 ? 4'h9 : add_83731[3:0]];
  assign array_index_83735 = array_update_83732[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_83739 = smul32b_32b_x_32b(array_index_82832[add_83731 > 32'h0000_0009 ? 4'h9 : add_83731[3:0]], array_index_83734[add_83638 > 32'h0000_0009 ? 4'h9 : add_83638[3:0]]);
  assign add_83741 = array_index_83735[add_83638 > 32'h0000_0009 ? 4'h9 : add_83638[3:0]] + smul_83739;
  assign array_update_83743[0] = add_83638 == 32'h0000_0000 ? add_83741 : array_index_83735[0];
  assign array_update_83743[1] = add_83638 == 32'h0000_0001 ? add_83741 : array_index_83735[1];
  assign array_update_83743[2] = add_83638 == 32'h0000_0002 ? add_83741 : array_index_83735[2];
  assign array_update_83743[3] = add_83638 == 32'h0000_0003 ? add_83741 : array_index_83735[3];
  assign array_update_83743[4] = add_83638 == 32'h0000_0004 ? add_83741 : array_index_83735[4];
  assign array_update_83743[5] = add_83638 == 32'h0000_0005 ? add_83741 : array_index_83735[5];
  assign array_update_83743[6] = add_83638 == 32'h0000_0006 ? add_83741 : array_index_83735[6];
  assign array_update_83743[7] = add_83638 == 32'h0000_0007 ? add_83741 : array_index_83735[7];
  assign array_update_83743[8] = add_83638 == 32'h0000_0008 ? add_83741 : array_index_83735[8];
  assign array_update_83743[9] = add_83638 == 32'h0000_0009 ? add_83741 : array_index_83735[9];
  assign add_83744 = add_83731 + 32'h0000_0001;
  assign array_update_83745[0] = add_82825 == 32'h0000_0000 ? array_update_83743 : array_update_83732[0];
  assign array_update_83745[1] = add_82825 == 32'h0000_0001 ? array_update_83743 : array_update_83732[1];
  assign array_update_83745[2] = add_82825 == 32'h0000_0002 ? array_update_83743 : array_update_83732[2];
  assign array_update_83745[3] = add_82825 == 32'h0000_0003 ? array_update_83743 : array_update_83732[3];
  assign array_update_83745[4] = add_82825 == 32'h0000_0004 ? array_update_83743 : array_update_83732[4];
  assign array_update_83745[5] = add_82825 == 32'h0000_0005 ? array_update_83743 : array_update_83732[5];
  assign array_update_83745[6] = add_82825 == 32'h0000_0006 ? array_update_83743 : array_update_83732[6];
  assign array_update_83745[7] = add_82825 == 32'h0000_0007 ? array_update_83743 : array_update_83732[7];
  assign array_update_83745[8] = add_82825 == 32'h0000_0008 ? array_update_83743 : array_update_83732[8];
  assign array_update_83745[9] = add_82825 == 32'h0000_0009 ? array_update_83743 : array_update_83732[9];
  assign array_index_83747 = array_update_72021[add_83744 > 32'h0000_0009 ? 4'h9 : add_83744[3:0]];
  assign array_index_83748 = array_update_83745[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_83752 = smul32b_32b_x_32b(array_index_82832[add_83744 > 32'h0000_0009 ? 4'h9 : add_83744[3:0]], array_index_83747[add_83638 > 32'h0000_0009 ? 4'h9 : add_83638[3:0]]);
  assign add_83754 = array_index_83748[add_83638 > 32'h0000_0009 ? 4'h9 : add_83638[3:0]] + smul_83752;
  assign array_update_83756[0] = add_83638 == 32'h0000_0000 ? add_83754 : array_index_83748[0];
  assign array_update_83756[1] = add_83638 == 32'h0000_0001 ? add_83754 : array_index_83748[1];
  assign array_update_83756[2] = add_83638 == 32'h0000_0002 ? add_83754 : array_index_83748[2];
  assign array_update_83756[3] = add_83638 == 32'h0000_0003 ? add_83754 : array_index_83748[3];
  assign array_update_83756[4] = add_83638 == 32'h0000_0004 ? add_83754 : array_index_83748[4];
  assign array_update_83756[5] = add_83638 == 32'h0000_0005 ? add_83754 : array_index_83748[5];
  assign array_update_83756[6] = add_83638 == 32'h0000_0006 ? add_83754 : array_index_83748[6];
  assign array_update_83756[7] = add_83638 == 32'h0000_0007 ? add_83754 : array_index_83748[7];
  assign array_update_83756[8] = add_83638 == 32'h0000_0008 ? add_83754 : array_index_83748[8];
  assign array_update_83756[9] = add_83638 == 32'h0000_0009 ? add_83754 : array_index_83748[9];
  assign add_83757 = add_83744 + 32'h0000_0001;
  assign array_update_83758[0] = add_82825 == 32'h0000_0000 ? array_update_83756 : array_update_83745[0];
  assign array_update_83758[1] = add_82825 == 32'h0000_0001 ? array_update_83756 : array_update_83745[1];
  assign array_update_83758[2] = add_82825 == 32'h0000_0002 ? array_update_83756 : array_update_83745[2];
  assign array_update_83758[3] = add_82825 == 32'h0000_0003 ? array_update_83756 : array_update_83745[3];
  assign array_update_83758[4] = add_82825 == 32'h0000_0004 ? array_update_83756 : array_update_83745[4];
  assign array_update_83758[5] = add_82825 == 32'h0000_0005 ? array_update_83756 : array_update_83745[5];
  assign array_update_83758[6] = add_82825 == 32'h0000_0006 ? array_update_83756 : array_update_83745[6];
  assign array_update_83758[7] = add_82825 == 32'h0000_0007 ? array_update_83756 : array_update_83745[7];
  assign array_update_83758[8] = add_82825 == 32'h0000_0008 ? array_update_83756 : array_update_83745[8];
  assign array_update_83758[9] = add_82825 == 32'h0000_0009 ? array_update_83756 : array_update_83745[9];
  assign array_index_83760 = array_update_72021[add_83757 > 32'h0000_0009 ? 4'h9 : add_83757[3:0]];
  assign array_index_83761 = array_update_83758[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_83765 = smul32b_32b_x_32b(array_index_82832[add_83757 > 32'h0000_0009 ? 4'h9 : add_83757[3:0]], array_index_83760[add_83638 > 32'h0000_0009 ? 4'h9 : add_83638[3:0]]);
  assign add_83767 = array_index_83761[add_83638 > 32'h0000_0009 ? 4'h9 : add_83638[3:0]] + smul_83765;
  assign array_update_83768[0] = add_83638 == 32'h0000_0000 ? add_83767 : array_index_83761[0];
  assign array_update_83768[1] = add_83638 == 32'h0000_0001 ? add_83767 : array_index_83761[1];
  assign array_update_83768[2] = add_83638 == 32'h0000_0002 ? add_83767 : array_index_83761[2];
  assign array_update_83768[3] = add_83638 == 32'h0000_0003 ? add_83767 : array_index_83761[3];
  assign array_update_83768[4] = add_83638 == 32'h0000_0004 ? add_83767 : array_index_83761[4];
  assign array_update_83768[5] = add_83638 == 32'h0000_0005 ? add_83767 : array_index_83761[5];
  assign array_update_83768[6] = add_83638 == 32'h0000_0006 ? add_83767 : array_index_83761[6];
  assign array_update_83768[7] = add_83638 == 32'h0000_0007 ? add_83767 : array_index_83761[7];
  assign array_update_83768[8] = add_83638 == 32'h0000_0008 ? add_83767 : array_index_83761[8];
  assign array_update_83768[9] = add_83638 == 32'h0000_0009 ? add_83767 : array_index_83761[9];
  assign array_update_83769[0] = add_82825 == 32'h0000_0000 ? array_update_83768 : array_update_83758[0];
  assign array_update_83769[1] = add_82825 == 32'h0000_0001 ? array_update_83768 : array_update_83758[1];
  assign array_update_83769[2] = add_82825 == 32'h0000_0002 ? array_update_83768 : array_update_83758[2];
  assign array_update_83769[3] = add_82825 == 32'h0000_0003 ? array_update_83768 : array_update_83758[3];
  assign array_update_83769[4] = add_82825 == 32'h0000_0004 ? array_update_83768 : array_update_83758[4];
  assign array_update_83769[5] = add_82825 == 32'h0000_0005 ? array_update_83768 : array_update_83758[5];
  assign array_update_83769[6] = add_82825 == 32'h0000_0006 ? array_update_83768 : array_update_83758[6];
  assign array_update_83769[7] = add_82825 == 32'h0000_0007 ? array_update_83768 : array_update_83758[7];
  assign array_update_83769[8] = add_82825 == 32'h0000_0008 ? array_update_83768 : array_update_83758[8];
  assign array_update_83769[9] = add_82825 == 32'h0000_0009 ? array_update_83768 : array_update_83758[9];
  assign array_index_83771 = array_update_83769[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign add_83773 = add_83638 + 32'h0000_0001;
  assign array_update_83774[0] = add_83773 == 32'h0000_0000 ? 32'h0000_0000 : array_index_83771[0];
  assign array_update_83774[1] = add_83773 == 32'h0000_0001 ? 32'h0000_0000 : array_index_83771[1];
  assign array_update_83774[2] = add_83773 == 32'h0000_0002 ? 32'h0000_0000 : array_index_83771[2];
  assign array_update_83774[3] = add_83773 == 32'h0000_0003 ? 32'h0000_0000 : array_index_83771[3];
  assign array_update_83774[4] = add_83773 == 32'h0000_0004 ? 32'h0000_0000 : array_index_83771[4];
  assign array_update_83774[5] = add_83773 == 32'h0000_0005 ? 32'h0000_0000 : array_index_83771[5];
  assign array_update_83774[6] = add_83773 == 32'h0000_0006 ? 32'h0000_0000 : array_index_83771[6];
  assign array_update_83774[7] = add_83773 == 32'h0000_0007 ? 32'h0000_0000 : array_index_83771[7];
  assign array_update_83774[8] = add_83773 == 32'h0000_0008 ? 32'h0000_0000 : array_index_83771[8];
  assign array_update_83774[9] = add_83773 == 32'h0000_0009 ? 32'h0000_0000 : array_index_83771[9];
  assign literal_83775 = 32'h0000_0000;
  assign array_update_83776[0] = add_82825 == 32'h0000_0000 ? array_update_83774 : array_update_83769[0];
  assign array_update_83776[1] = add_82825 == 32'h0000_0001 ? array_update_83774 : array_update_83769[1];
  assign array_update_83776[2] = add_82825 == 32'h0000_0002 ? array_update_83774 : array_update_83769[2];
  assign array_update_83776[3] = add_82825 == 32'h0000_0003 ? array_update_83774 : array_update_83769[3];
  assign array_update_83776[4] = add_82825 == 32'h0000_0004 ? array_update_83774 : array_update_83769[4];
  assign array_update_83776[5] = add_82825 == 32'h0000_0005 ? array_update_83774 : array_update_83769[5];
  assign array_update_83776[6] = add_82825 == 32'h0000_0006 ? array_update_83774 : array_update_83769[6];
  assign array_update_83776[7] = add_82825 == 32'h0000_0007 ? array_update_83774 : array_update_83769[7];
  assign array_update_83776[8] = add_82825 == 32'h0000_0008 ? array_update_83774 : array_update_83769[8];
  assign array_update_83776[9] = add_82825 == 32'h0000_0009 ? array_update_83774 : array_update_83769[9];
  assign array_index_83778 = array_update_72021[literal_83775 > 32'h0000_0009 ? 4'h9 : literal_83775[3:0]];
  assign array_index_83779 = array_update_83776[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_83783 = smul32b_32b_x_32b(array_index_82832[literal_83775 > 32'h0000_0009 ? 4'h9 : literal_83775[3:0]], array_index_83778[add_83773 > 32'h0000_0009 ? 4'h9 : add_83773[3:0]]);
  assign add_83785 = array_index_83779[add_83773 > 32'h0000_0009 ? 4'h9 : add_83773[3:0]] + smul_83783;
  assign array_update_83787[0] = add_83773 == 32'h0000_0000 ? add_83785 : array_index_83779[0];
  assign array_update_83787[1] = add_83773 == 32'h0000_0001 ? add_83785 : array_index_83779[1];
  assign array_update_83787[2] = add_83773 == 32'h0000_0002 ? add_83785 : array_index_83779[2];
  assign array_update_83787[3] = add_83773 == 32'h0000_0003 ? add_83785 : array_index_83779[3];
  assign array_update_83787[4] = add_83773 == 32'h0000_0004 ? add_83785 : array_index_83779[4];
  assign array_update_83787[5] = add_83773 == 32'h0000_0005 ? add_83785 : array_index_83779[5];
  assign array_update_83787[6] = add_83773 == 32'h0000_0006 ? add_83785 : array_index_83779[6];
  assign array_update_83787[7] = add_83773 == 32'h0000_0007 ? add_83785 : array_index_83779[7];
  assign array_update_83787[8] = add_83773 == 32'h0000_0008 ? add_83785 : array_index_83779[8];
  assign array_update_83787[9] = add_83773 == 32'h0000_0009 ? add_83785 : array_index_83779[9];
  assign add_83788 = literal_83775 + 32'h0000_0001;
  assign array_update_83789[0] = add_82825 == 32'h0000_0000 ? array_update_83787 : array_update_83776[0];
  assign array_update_83789[1] = add_82825 == 32'h0000_0001 ? array_update_83787 : array_update_83776[1];
  assign array_update_83789[2] = add_82825 == 32'h0000_0002 ? array_update_83787 : array_update_83776[2];
  assign array_update_83789[3] = add_82825 == 32'h0000_0003 ? array_update_83787 : array_update_83776[3];
  assign array_update_83789[4] = add_82825 == 32'h0000_0004 ? array_update_83787 : array_update_83776[4];
  assign array_update_83789[5] = add_82825 == 32'h0000_0005 ? array_update_83787 : array_update_83776[5];
  assign array_update_83789[6] = add_82825 == 32'h0000_0006 ? array_update_83787 : array_update_83776[6];
  assign array_update_83789[7] = add_82825 == 32'h0000_0007 ? array_update_83787 : array_update_83776[7];
  assign array_update_83789[8] = add_82825 == 32'h0000_0008 ? array_update_83787 : array_update_83776[8];
  assign array_update_83789[9] = add_82825 == 32'h0000_0009 ? array_update_83787 : array_update_83776[9];
  assign array_index_83791 = array_update_72021[add_83788 > 32'h0000_0009 ? 4'h9 : add_83788[3:0]];
  assign array_index_83792 = array_update_83789[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_83796 = smul32b_32b_x_32b(array_index_82832[add_83788 > 32'h0000_0009 ? 4'h9 : add_83788[3:0]], array_index_83791[add_83773 > 32'h0000_0009 ? 4'h9 : add_83773[3:0]]);
  assign add_83798 = array_index_83792[add_83773 > 32'h0000_0009 ? 4'h9 : add_83773[3:0]] + smul_83796;
  assign array_update_83800[0] = add_83773 == 32'h0000_0000 ? add_83798 : array_index_83792[0];
  assign array_update_83800[1] = add_83773 == 32'h0000_0001 ? add_83798 : array_index_83792[1];
  assign array_update_83800[2] = add_83773 == 32'h0000_0002 ? add_83798 : array_index_83792[2];
  assign array_update_83800[3] = add_83773 == 32'h0000_0003 ? add_83798 : array_index_83792[3];
  assign array_update_83800[4] = add_83773 == 32'h0000_0004 ? add_83798 : array_index_83792[4];
  assign array_update_83800[5] = add_83773 == 32'h0000_0005 ? add_83798 : array_index_83792[5];
  assign array_update_83800[6] = add_83773 == 32'h0000_0006 ? add_83798 : array_index_83792[6];
  assign array_update_83800[7] = add_83773 == 32'h0000_0007 ? add_83798 : array_index_83792[7];
  assign array_update_83800[8] = add_83773 == 32'h0000_0008 ? add_83798 : array_index_83792[8];
  assign array_update_83800[9] = add_83773 == 32'h0000_0009 ? add_83798 : array_index_83792[9];
  assign add_83801 = add_83788 + 32'h0000_0001;
  assign array_update_83802[0] = add_82825 == 32'h0000_0000 ? array_update_83800 : array_update_83789[0];
  assign array_update_83802[1] = add_82825 == 32'h0000_0001 ? array_update_83800 : array_update_83789[1];
  assign array_update_83802[2] = add_82825 == 32'h0000_0002 ? array_update_83800 : array_update_83789[2];
  assign array_update_83802[3] = add_82825 == 32'h0000_0003 ? array_update_83800 : array_update_83789[3];
  assign array_update_83802[4] = add_82825 == 32'h0000_0004 ? array_update_83800 : array_update_83789[4];
  assign array_update_83802[5] = add_82825 == 32'h0000_0005 ? array_update_83800 : array_update_83789[5];
  assign array_update_83802[6] = add_82825 == 32'h0000_0006 ? array_update_83800 : array_update_83789[6];
  assign array_update_83802[7] = add_82825 == 32'h0000_0007 ? array_update_83800 : array_update_83789[7];
  assign array_update_83802[8] = add_82825 == 32'h0000_0008 ? array_update_83800 : array_update_83789[8];
  assign array_update_83802[9] = add_82825 == 32'h0000_0009 ? array_update_83800 : array_update_83789[9];
  assign array_index_83804 = array_update_72021[add_83801 > 32'h0000_0009 ? 4'h9 : add_83801[3:0]];
  assign array_index_83805 = array_update_83802[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_83809 = smul32b_32b_x_32b(array_index_82832[add_83801 > 32'h0000_0009 ? 4'h9 : add_83801[3:0]], array_index_83804[add_83773 > 32'h0000_0009 ? 4'h9 : add_83773[3:0]]);
  assign add_83811 = array_index_83805[add_83773 > 32'h0000_0009 ? 4'h9 : add_83773[3:0]] + smul_83809;
  assign array_update_83813[0] = add_83773 == 32'h0000_0000 ? add_83811 : array_index_83805[0];
  assign array_update_83813[1] = add_83773 == 32'h0000_0001 ? add_83811 : array_index_83805[1];
  assign array_update_83813[2] = add_83773 == 32'h0000_0002 ? add_83811 : array_index_83805[2];
  assign array_update_83813[3] = add_83773 == 32'h0000_0003 ? add_83811 : array_index_83805[3];
  assign array_update_83813[4] = add_83773 == 32'h0000_0004 ? add_83811 : array_index_83805[4];
  assign array_update_83813[5] = add_83773 == 32'h0000_0005 ? add_83811 : array_index_83805[5];
  assign array_update_83813[6] = add_83773 == 32'h0000_0006 ? add_83811 : array_index_83805[6];
  assign array_update_83813[7] = add_83773 == 32'h0000_0007 ? add_83811 : array_index_83805[7];
  assign array_update_83813[8] = add_83773 == 32'h0000_0008 ? add_83811 : array_index_83805[8];
  assign array_update_83813[9] = add_83773 == 32'h0000_0009 ? add_83811 : array_index_83805[9];
  assign add_83814 = add_83801 + 32'h0000_0001;
  assign array_update_83815[0] = add_82825 == 32'h0000_0000 ? array_update_83813 : array_update_83802[0];
  assign array_update_83815[1] = add_82825 == 32'h0000_0001 ? array_update_83813 : array_update_83802[1];
  assign array_update_83815[2] = add_82825 == 32'h0000_0002 ? array_update_83813 : array_update_83802[2];
  assign array_update_83815[3] = add_82825 == 32'h0000_0003 ? array_update_83813 : array_update_83802[3];
  assign array_update_83815[4] = add_82825 == 32'h0000_0004 ? array_update_83813 : array_update_83802[4];
  assign array_update_83815[5] = add_82825 == 32'h0000_0005 ? array_update_83813 : array_update_83802[5];
  assign array_update_83815[6] = add_82825 == 32'h0000_0006 ? array_update_83813 : array_update_83802[6];
  assign array_update_83815[7] = add_82825 == 32'h0000_0007 ? array_update_83813 : array_update_83802[7];
  assign array_update_83815[8] = add_82825 == 32'h0000_0008 ? array_update_83813 : array_update_83802[8];
  assign array_update_83815[9] = add_82825 == 32'h0000_0009 ? array_update_83813 : array_update_83802[9];
  assign array_index_83817 = array_update_72021[add_83814 > 32'h0000_0009 ? 4'h9 : add_83814[3:0]];
  assign array_index_83818 = array_update_83815[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_83822 = smul32b_32b_x_32b(array_index_82832[add_83814 > 32'h0000_0009 ? 4'h9 : add_83814[3:0]], array_index_83817[add_83773 > 32'h0000_0009 ? 4'h9 : add_83773[3:0]]);
  assign add_83824 = array_index_83818[add_83773 > 32'h0000_0009 ? 4'h9 : add_83773[3:0]] + smul_83822;
  assign array_update_83826[0] = add_83773 == 32'h0000_0000 ? add_83824 : array_index_83818[0];
  assign array_update_83826[1] = add_83773 == 32'h0000_0001 ? add_83824 : array_index_83818[1];
  assign array_update_83826[2] = add_83773 == 32'h0000_0002 ? add_83824 : array_index_83818[2];
  assign array_update_83826[3] = add_83773 == 32'h0000_0003 ? add_83824 : array_index_83818[3];
  assign array_update_83826[4] = add_83773 == 32'h0000_0004 ? add_83824 : array_index_83818[4];
  assign array_update_83826[5] = add_83773 == 32'h0000_0005 ? add_83824 : array_index_83818[5];
  assign array_update_83826[6] = add_83773 == 32'h0000_0006 ? add_83824 : array_index_83818[6];
  assign array_update_83826[7] = add_83773 == 32'h0000_0007 ? add_83824 : array_index_83818[7];
  assign array_update_83826[8] = add_83773 == 32'h0000_0008 ? add_83824 : array_index_83818[8];
  assign array_update_83826[9] = add_83773 == 32'h0000_0009 ? add_83824 : array_index_83818[9];
  assign add_83827 = add_83814 + 32'h0000_0001;
  assign array_update_83828[0] = add_82825 == 32'h0000_0000 ? array_update_83826 : array_update_83815[0];
  assign array_update_83828[1] = add_82825 == 32'h0000_0001 ? array_update_83826 : array_update_83815[1];
  assign array_update_83828[2] = add_82825 == 32'h0000_0002 ? array_update_83826 : array_update_83815[2];
  assign array_update_83828[3] = add_82825 == 32'h0000_0003 ? array_update_83826 : array_update_83815[3];
  assign array_update_83828[4] = add_82825 == 32'h0000_0004 ? array_update_83826 : array_update_83815[4];
  assign array_update_83828[5] = add_82825 == 32'h0000_0005 ? array_update_83826 : array_update_83815[5];
  assign array_update_83828[6] = add_82825 == 32'h0000_0006 ? array_update_83826 : array_update_83815[6];
  assign array_update_83828[7] = add_82825 == 32'h0000_0007 ? array_update_83826 : array_update_83815[7];
  assign array_update_83828[8] = add_82825 == 32'h0000_0008 ? array_update_83826 : array_update_83815[8];
  assign array_update_83828[9] = add_82825 == 32'h0000_0009 ? array_update_83826 : array_update_83815[9];
  assign array_index_83830 = array_update_72021[add_83827 > 32'h0000_0009 ? 4'h9 : add_83827[3:0]];
  assign array_index_83831 = array_update_83828[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_83835 = smul32b_32b_x_32b(array_index_82832[add_83827 > 32'h0000_0009 ? 4'h9 : add_83827[3:0]], array_index_83830[add_83773 > 32'h0000_0009 ? 4'h9 : add_83773[3:0]]);
  assign add_83837 = array_index_83831[add_83773 > 32'h0000_0009 ? 4'h9 : add_83773[3:0]] + smul_83835;
  assign array_update_83839[0] = add_83773 == 32'h0000_0000 ? add_83837 : array_index_83831[0];
  assign array_update_83839[1] = add_83773 == 32'h0000_0001 ? add_83837 : array_index_83831[1];
  assign array_update_83839[2] = add_83773 == 32'h0000_0002 ? add_83837 : array_index_83831[2];
  assign array_update_83839[3] = add_83773 == 32'h0000_0003 ? add_83837 : array_index_83831[3];
  assign array_update_83839[4] = add_83773 == 32'h0000_0004 ? add_83837 : array_index_83831[4];
  assign array_update_83839[5] = add_83773 == 32'h0000_0005 ? add_83837 : array_index_83831[5];
  assign array_update_83839[6] = add_83773 == 32'h0000_0006 ? add_83837 : array_index_83831[6];
  assign array_update_83839[7] = add_83773 == 32'h0000_0007 ? add_83837 : array_index_83831[7];
  assign array_update_83839[8] = add_83773 == 32'h0000_0008 ? add_83837 : array_index_83831[8];
  assign array_update_83839[9] = add_83773 == 32'h0000_0009 ? add_83837 : array_index_83831[9];
  assign add_83840 = add_83827 + 32'h0000_0001;
  assign array_update_83841[0] = add_82825 == 32'h0000_0000 ? array_update_83839 : array_update_83828[0];
  assign array_update_83841[1] = add_82825 == 32'h0000_0001 ? array_update_83839 : array_update_83828[1];
  assign array_update_83841[2] = add_82825 == 32'h0000_0002 ? array_update_83839 : array_update_83828[2];
  assign array_update_83841[3] = add_82825 == 32'h0000_0003 ? array_update_83839 : array_update_83828[3];
  assign array_update_83841[4] = add_82825 == 32'h0000_0004 ? array_update_83839 : array_update_83828[4];
  assign array_update_83841[5] = add_82825 == 32'h0000_0005 ? array_update_83839 : array_update_83828[5];
  assign array_update_83841[6] = add_82825 == 32'h0000_0006 ? array_update_83839 : array_update_83828[6];
  assign array_update_83841[7] = add_82825 == 32'h0000_0007 ? array_update_83839 : array_update_83828[7];
  assign array_update_83841[8] = add_82825 == 32'h0000_0008 ? array_update_83839 : array_update_83828[8];
  assign array_update_83841[9] = add_82825 == 32'h0000_0009 ? array_update_83839 : array_update_83828[9];
  assign array_index_83843 = array_update_72021[add_83840 > 32'h0000_0009 ? 4'h9 : add_83840[3:0]];
  assign array_index_83844 = array_update_83841[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_83848 = smul32b_32b_x_32b(array_index_82832[add_83840 > 32'h0000_0009 ? 4'h9 : add_83840[3:0]], array_index_83843[add_83773 > 32'h0000_0009 ? 4'h9 : add_83773[3:0]]);
  assign add_83850 = array_index_83844[add_83773 > 32'h0000_0009 ? 4'h9 : add_83773[3:0]] + smul_83848;
  assign array_update_83852[0] = add_83773 == 32'h0000_0000 ? add_83850 : array_index_83844[0];
  assign array_update_83852[1] = add_83773 == 32'h0000_0001 ? add_83850 : array_index_83844[1];
  assign array_update_83852[2] = add_83773 == 32'h0000_0002 ? add_83850 : array_index_83844[2];
  assign array_update_83852[3] = add_83773 == 32'h0000_0003 ? add_83850 : array_index_83844[3];
  assign array_update_83852[4] = add_83773 == 32'h0000_0004 ? add_83850 : array_index_83844[4];
  assign array_update_83852[5] = add_83773 == 32'h0000_0005 ? add_83850 : array_index_83844[5];
  assign array_update_83852[6] = add_83773 == 32'h0000_0006 ? add_83850 : array_index_83844[6];
  assign array_update_83852[7] = add_83773 == 32'h0000_0007 ? add_83850 : array_index_83844[7];
  assign array_update_83852[8] = add_83773 == 32'h0000_0008 ? add_83850 : array_index_83844[8];
  assign array_update_83852[9] = add_83773 == 32'h0000_0009 ? add_83850 : array_index_83844[9];
  assign add_83853 = add_83840 + 32'h0000_0001;
  assign array_update_83854[0] = add_82825 == 32'h0000_0000 ? array_update_83852 : array_update_83841[0];
  assign array_update_83854[1] = add_82825 == 32'h0000_0001 ? array_update_83852 : array_update_83841[1];
  assign array_update_83854[2] = add_82825 == 32'h0000_0002 ? array_update_83852 : array_update_83841[2];
  assign array_update_83854[3] = add_82825 == 32'h0000_0003 ? array_update_83852 : array_update_83841[3];
  assign array_update_83854[4] = add_82825 == 32'h0000_0004 ? array_update_83852 : array_update_83841[4];
  assign array_update_83854[5] = add_82825 == 32'h0000_0005 ? array_update_83852 : array_update_83841[5];
  assign array_update_83854[6] = add_82825 == 32'h0000_0006 ? array_update_83852 : array_update_83841[6];
  assign array_update_83854[7] = add_82825 == 32'h0000_0007 ? array_update_83852 : array_update_83841[7];
  assign array_update_83854[8] = add_82825 == 32'h0000_0008 ? array_update_83852 : array_update_83841[8];
  assign array_update_83854[9] = add_82825 == 32'h0000_0009 ? array_update_83852 : array_update_83841[9];
  assign array_index_83856 = array_update_72021[add_83853 > 32'h0000_0009 ? 4'h9 : add_83853[3:0]];
  assign array_index_83857 = array_update_83854[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_83861 = smul32b_32b_x_32b(array_index_82832[add_83853 > 32'h0000_0009 ? 4'h9 : add_83853[3:0]], array_index_83856[add_83773 > 32'h0000_0009 ? 4'h9 : add_83773[3:0]]);
  assign add_83863 = array_index_83857[add_83773 > 32'h0000_0009 ? 4'h9 : add_83773[3:0]] + smul_83861;
  assign array_update_83865[0] = add_83773 == 32'h0000_0000 ? add_83863 : array_index_83857[0];
  assign array_update_83865[1] = add_83773 == 32'h0000_0001 ? add_83863 : array_index_83857[1];
  assign array_update_83865[2] = add_83773 == 32'h0000_0002 ? add_83863 : array_index_83857[2];
  assign array_update_83865[3] = add_83773 == 32'h0000_0003 ? add_83863 : array_index_83857[3];
  assign array_update_83865[4] = add_83773 == 32'h0000_0004 ? add_83863 : array_index_83857[4];
  assign array_update_83865[5] = add_83773 == 32'h0000_0005 ? add_83863 : array_index_83857[5];
  assign array_update_83865[6] = add_83773 == 32'h0000_0006 ? add_83863 : array_index_83857[6];
  assign array_update_83865[7] = add_83773 == 32'h0000_0007 ? add_83863 : array_index_83857[7];
  assign array_update_83865[8] = add_83773 == 32'h0000_0008 ? add_83863 : array_index_83857[8];
  assign array_update_83865[9] = add_83773 == 32'h0000_0009 ? add_83863 : array_index_83857[9];
  assign add_83866 = add_83853 + 32'h0000_0001;
  assign array_update_83867[0] = add_82825 == 32'h0000_0000 ? array_update_83865 : array_update_83854[0];
  assign array_update_83867[1] = add_82825 == 32'h0000_0001 ? array_update_83865 : array_update_83854[1];
  assign array_update_83867[2] = add_82825 == 32'h0000_0002 ? array_update_83865 : array_update_83854[2];
  assign array_update_83867[3] = add_82825 == 32'h0000_0003 ? array_update_83865 : array_update_83854[3];
  assign array_update_83867[4] = add_82825 == 32'h0000_0004 ? array_update_83865 : array_update_83854[4];
  assign array_update_83867[5] = add_82825 == 32'h0000_0005 ? array_update_83865 : array_update_83854[5];
  assign array_update_83867[6] = add_82825 == 32'h0000_0006 ? array_update_83865 : array_update_83854[6];
  assign array_update_83867[7] = add_82825 == 32'h0000_0007 ? array_update_83865 : array_update_83854[7];
  assign array_update_83867[8] = add_82825 == 32'h0000_0008 ? array_update_83865 : array_update_83854[8];
  assign array_update_83867[9] = add_82825 == 32'h0000_0009 ? array_update_83865 : array_update_83854[9];
  assign array_index_83869 = array_update_72021[add_83866 > 32'h0000_0009 ? 4'h9 : add_83866[3:0]];
  assign array_index_83870 = array_update_83867[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_83874 = smul32b_32b_x_32b(array_index_82832[add_83866 > 32'h0000_0009 ? 4'h9 : add_83866[3:0]], array_index_83869[add_83773 > 32'h0000_0009 ? 4'h9 : add_83773[3:0]]);
  assign add_83876 = array_index_83870[add_83773 > 32'h0000_0009 ? 4'h9 : add_83773[3:0]] + smul_83874;
  assign array_update_83878[0] = add_83773 == 32'h0000_0000 ? add_83876 : array_index_83870[0];
  assign array_update_83878[1] = add_83773 == 32'h0000_0001 ? add_83876 : array_index_83870[1];
  assign array_update_83878[2] = add_83773 == 32'h0000_0002 ? add_83876 : array_index_83870[2];
  assign array_update_83878[3] = add_83773 == 32'h0000_0003 ? add_83876 : array_index_83870[3];
  assign array_update_83878[4] = add_83773 == 32'h0000_0004 ? add_83876 : array_index_83870[4];
  assign array_update_83878[5] = add_83773 == 32'h0000_0005 ? add_83876 : array_index_83870[5];
  assign array_update_83878[6] = add_83773 == 32'h0000_0006 ? add_83876 : array_index_83870[6];
  assign array_update_83878[7] = add_83773 == 32'h0000_0007 ? add_83876 : array_index_83870[7];
  assign array_update_83878[8] = add_83773 == 32'h0000_0008 ? add_83876 : array_index_83870[8];
  assign array_update_83878[9] = add_83773 == 32'h0000_0009 ? add_83876 : array_index_83870[9];
  assign add_83879 = add_83866 + 32'h0000_0001;
  assign array_update_83880[0] = add_82825 == 32'h0000_0000 ? array_update_83878 : array_update_83867[0];
  assign array_update_83880[1] = add_82825 == 32'h0000_0001 ? array_update_83878 : array_update_83867[1];
  assign array_update_83880[2] = add_82825 == 32'h0000_0002 ? array_update_83878 : array_update_83867[2];
  assign array_update_83880[3] = add_82825 == 32'h0000_0003 ? array_update_83878 : array_update_83867[3];
  assign array_update_83880[4] = add_82825 == 32'h0000_0004 ? array_update_83878 : array_update_83867[4];
  assign array_update_83880[5] = add_82825 == 32'h0000_0005 ? array_update_83878 : array_update_83867[5];
  assign array_update_83880[6] = add_82825 == 32'h0000_0006 ? array_update_83878 : array_update_83867[6];
  assign array_update_83880[7] = add_82825 == 32'h0000_0007 ? array_update_83878 : array_update_83867[7];
  assign array_update_83880[8] = add_82825 == 32'h0000_0008 ? array_update_83878 : array_update_83867[8];
  assign array_update_83880[9] = add_82825 == 32'h0000_0009 ? array_update_83878 : array_update_83867[9];
  assign array_index_83882 = array_update_72021[add_83879 > 32'h0000_0009 ? 4'h9 : add_83879[3:0]];
  assign array_index_83883 = array_update_83880[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_83887 = smul32b_32b_x_32b(array_index_82832[add_83879 > 32'h0000_0009 ? 4'h9 : add_83879[3:0]], array_index_83882[add_83773 > 32'h0000_0009 ? 4'h9 : add_83773[3:0]]);
  assign add_83889 = array_index_83883[add_83773 > 32'h0000_0009 ? 4'h9 : add_83773[3:0]] + smul_83887;
  assign array_update_83891[0] = add_83773 == 32'h0000_0000 ? add_83889 : array_index_83883[0];
  assign array_update_83891[1] = add_83773 == 32'h0000_0001 ? add_83889 : array_index_83883[1];
  assign array_update_83891[2] = add_83773 == 32'h0000_0002 ? add_83889 : array_index_83883[2];
  assign array_update_83891[3] = add_83773 == 32'h0000_0003 ? add_83889 : array_index_83883[3];
  assign array_update_83891[4] = add_83773 == 32'h0000_0004 ? add_83889 : array_index_83883[4];
  assign array_update_83891[5] = add_83773 == 32'h0000_0005 ? add_83889 : array_index_83883[5];
  assign array_update_83891[6] = add_83773 == 32'h0000_0006 ? add_83889 : array_index_83883[6];
  assign array_update_83891[7] = add_83773 == 32'h0000_0007 ? add_83889 : array_index_83883[7];
  assign array_update_83891[8] = add_83773 == 32'h0000_0008 ? add_83889 : array_index_83883[8];
  assign array_update_83891[9] = add_83773 == 32'h0000_0009 ? add_83889 : array_index_83883[9];
  assign add_83892 = add_83879 + 32'h0000_0001;
  assign array_update_83893[0] = add_82825 == 32'h0000_0000 ? array_update_83891 : array_update_83880[0];
  assign array_update_83893[1] = add_82825 == 32'h0000_0001 ? array_update_83891 : array_update_83880[1];
  assign array_update_83893[2] = add_82825 == 32'h0000_0002 ? array_update_83891 : array_update_83880[2];
  assign array_update_83893[3] = add_82825 == 32'h0000_0003 ? array_update_83891 : array_update_83880[3];
  assign array_update_83893[4] = add_82825 == 32'h0000_0004 ? array_update_83891 : array_update_83880[4];
  assign array_update_83893[5] = add_82825 == 32'h0000_0005 ? array_update_83891 : array_update_83880[5];
  assign array_update_83893[6] = add_82825 == 32'h0000_0006 ? array_update_83891 : array_update_83880[6];
  assign array_update_83893[7] = add_82825 == 32'h0000_0007 ? array_update_83891 : array_update_83880[7];
  assign array_update_83893[8] = add_82825 == 32'h0000_0008 ? array_update_83891 : array_update_83880[8];
  assign array_update_83893[9] = add_82825 == 32'h0000_0009 ? array_update_83891 : array_update_83880[9];
  assign array_index_83895 = array_update_72021[add_83892 > 32'h0000_0009 ? 4'h9 : add_83892[3:0]];
  assign array_index_83896 = array_update_83893[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_83900 = smul32b_32b_x_32b(array_index_82832[add_83892 > 32'h0000_0009 ? 4'h9 : add_83892[3:0]], array_index_83895[add_83773 > 32'h0000_0009 ? 4'h9 : add_83773[3:0]]);
  assign add_83902 = array_index_83896[add_83773 > 32'h0000_0009 ? 4'h9 : add_83773[3:0]] + smul_83900;
  assign array_update_83903[0] = add_83773 == 32'h0000_0000 ? add_83902 : array_index_83896[0];
  assign array_update_83903[1] = add_83773 == 32'h0000_0001 ? add_83902 : array_index_83896[1];
  assign array_update_83903[2] = add_83773 == 32'h0000_0002 ? add_83902 : array_index_83896[2];
  assign array_update_83903[3] = add_83773 == 32'h0000_0003 ? add_83902 : array_index_83896[3];
  assign array_update_83903[4] = add_83773 == 32'h0000_0004 ? add_83902 : array_index_83896[4];
  assign array_update_83903[5] = add_83773 == 32'h0000_0005 ? add_83902 : array_index_83896[5];
  assign array_update_83903[6] = add_83773 == 32'h0000_0006 ? add_83902 : array_index_83896[6];
  assign array_update_83903[7] = add_83773 == 32'h0000_0007 ? add_83902 : array_index_83896[7];
  assign array_update_83903[8] = add_83773 == 32'h0000_0008 ? add_83902 : array_index_83896[8];
  assign array_update_83903[9] = add_83773 == 32'h0000_0009 ? add_83902 : array_index_83896[9];
  assign array_update_83904[0] = add_82825 == 32'h0000_0000 ? array_update_83903 : array_update_83893[0];
  assign array_update_83904[1] = add_82825 == 32'h0000_0001 ? array_update_83903 : array_update_83893[1];
  assign array_update_83904[2] = add_82825 == 32'h0000_0002 ? array_update_83903 : array_update_83893[2];
  assign array_update_83904[3] = add_82825 == 32'h0000_0003 ? array_update_83903 : array_update_83893[3];
  assign array_update_83904[4] = add_82825 == 32'h0000_0004 ? array_update_83903 : array_update_83893[4];
  assign array_update_83904[5] = add_82825 == 32'h0000_0005 ? array_update_83903 : array_update_83893[5];
  assign array_update_83904[6] = add_82825 == 32'h0000_0006 ? array_update_83903 : array_update_83893[6];
  assign array_update_83904[7] = add_82825 == 32'h0000_0007 ? array_update_83903 : array_update_83893[7];
  assign array_update_83904[8] = add_82825 == 32'h0000_0008 ? array_update_83903 : array_update_83893[8];
  assign array_update_83904[9] = add_82825 == 32'h0000_0009 ? array_update_83903 : array_update_83893[9];
  assign array_index_83906 = array_update_83904[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign add_83908 = add_83773 + 32'h0000_0001;
  assign array_update_83909[0] = add_83908 == 32'h0000_0000 ? 32'h0000_0000 : array_index_83906[0];
  assign array_update_83909[1] = add_83908 == 32'h0000_0001 ? 32'h0000_0000 : array_index_83906[1];
  assign array_update_83909[2] = add_83908 == 32'h0000_0002 ? 32'h0000_0000 : array_index_83906[2];
  assign array_update_83909[3] = add_83908 == 32'h0000_0003 ? 32'h0000_0000 : array_index_83906[3];
  assign array_update_83909[4] = add_83908 == 32'h0000_0004 ? 32'h0000_0000 : array_index_83906[4];
  assign array_update_83909[5] = add_83908 == 32'h0000_0005 ? 32'h0000_0000 : array_index_83906[5];
  assign array_update_83909[6] = add_83908 == 32'h0000_0006 ? 32'h0000_0000 : array_index_83906[6];
  assign array_update_83909[7] = add_83908 == 32'h0000_0007 ? 32'h0000_0000 : array_index_83906[7];
  assign array_update_83909[8] = add_83908 == 32'h0000_0008 ? 32'h0000_0000 : array_index_83906[8];
  assign array_update_83909[9] = add_83908 == 32'h0000_0009 ? 32'h0000_0000 : array_index_83906[9];
  assign literal_83910 = 32'h0000_0000;
  assign array_update_83911[0] = add_82825 == 32'h0000_0000 ? array_update_83909 : array_update_83904[0];
  assign array_update_83911[1] = add_82825 == 32'h0000_0001 ? array_update_83909 : array_update_83904[1];
  assign array_update_83911[2] = add_82825 == 32'h0000_0002 ? array_update_83909 : array_update_83904[2];
  assign array_update_83911[3] = add_82825 == 32'h0000_0003 ? array_update_83909 : array_update_83904[3];
  assign array_update_83911[4] = add_82825 == 32'h0000_0004 ? array_update_83909 : array_update_83904[4];
  assign array_update_83911[5] = add_82825 == 32'h0000_0005 ? array_update_83909 : array_update_83904[5];
  assign array_update_83911[6] = add_82825 == 32'h0000_0006 ? array_update_83909 : array_update_83904[6];
  assign array_update_83911[7] = add_82825 == 32'h0000_0007 ? array_update_83909 : array_update_83904[7];
  assign array_update_83911[8] = add_82825 == 32'h0000_0008 ? array_update_83909 : array_update_83904[8];
  assign array_update_83911[9] = add_82825 == 32'h0000_0009 ? array_update_83909 : array_update_83904[9];
  assign array_index_83913 = array_update_72021[literal_83910 > 32'h0000_0009 ? 4'h9 : literal_83910[3:0]];
  assign array_index_83914 = array_update_83911[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_83918 = smul32b_32b_x_32b(array_index_82832[literal_83910 > 32'h0000_0009 ? 4'h9 : literal_83910[3:0]], array_index_83913[add_83908 > 32'h0000_0009 ? 4'h9 : add_83908[3:0]]);
  assign add_83920 = array_index_83914[add_83908 > 32'h0000_0009 ? 4'h9 : add_83908[3:0]] + smul_83918;
  assign array_update_83922[0] = add_83908 == 32'h0000_0000 ? add_83920 : array_index_83914[0];
  assign array_update_83922[1] = add_83908 == 32'h0000_0001 ? add_83920 : array_index_83914[1];
  assign array_update_83922[2] = add_83908 == 32'h0000_0002 ? add_83920 : array_index_83914[2];
  assign array_update_83922[3] = add_83908 == 32'h0000_0003 ? add_83920 : array_index_83914[3];
  assign array_update_83922[4] = add_83908 == 32'h0000_0004 ? add_83920 : array_index_83914[4];
  assign array_update_83922[5] = add_83908 == 32'h0000_0005 ? add_83920 : array_index_83914[5];
  assign array_update_83922[6] = add_83908 == 32'h0000_0006 ? add_83920 : array_index_83914[6];
  assign array_update_83922[7] = add_83908 == 32'h0000_0007 ? add_83920 : array_index_83914[7];
  assign array_update_83922[8] = add_83908 == 32'h0000_0008 ? add_83920 : array_index_83914[8];
  assign array_update_83922[9] = add_83908 == 32'h0000_0009 ? add_83920 : array_index_83914[9];
  assign add_83923 = literal_83910 + 32'h0000_0001;
  assign array_update_83924[0] = add_82825 == 32'h0000_0000 ? array_update_83922 : array_update_83911[0];
  assign array_update_83924[1] = add_82825 == 32'h0000_0001 ? array_update_83922 : array_update_83911[1];
  assign array_update_83924[2] = add_82825 == 32'h0000_0002 ? array_update_83922 : array_update_83911[2];
  assign array_update_83924[3] = add_82825 == 32'h0000_0003 ? array_update_83922 : array_update_83911[3];
  assign array_update_83924[4] = add_82825 == 32'h0000_0004 ? array_update_83922 : array_update_83911[4];
  assign array_update_83924[5] = add_82825 == 32'h0000_0005 ? array_update_83922 : array_update_83911[5];
  assign array_update_83924[6] = add_82825 == 32'h0000_0006 ? array_update_83922 : array_update_83911[6];
  assign array_update_83924[7] = add_82825 == 32'h0000_0007 ? array_update_83922 : array_update_83911[7];
  assign array_update_83924[8] = add_82825 == 32'h0000_0008 ? array_update_83922 : array_update_83911[8];
  assign array_update_83924[9] = add_82825 == 32'h0000_0009 ? array_update_83922 : array_update_83911[9];
  assign array_index_83926 = array_update_72021[add_83923 > 32'h0000_0009 ? 4'h9 : add_83923[3:0]];
  assign array_index_83927 = array_update_83924[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_83931 = smul32b_32b_x_32b(array_index_82832[add_83923 > 32'h0000_0009 ? 4'h9 : add_83923[3:0]], array_index_83926[add_83908 > 32'h0000_0009 ? 4'h9 : add_83908[3:0]]);
  assign add_83933 = array_index_83927[add_83908 > 32'h0000_0009 ? 4'h9 : add_83908[3:0]] + smul_83931;
  assign array_update_83935[0] = add_83908 == 32'h0000_0000 ? add_83933 : array_index_83927[0];
  assign array_update_83935[1] = add_83908 == 32'h0000_0001 ? add_83933 : array_index_83927[1];
  assign array_update_83935[2] = add_83908 == 32'h0000_0002 ? add_83933 : array_index_83927[2];
  assign array_update_83935[3] = add_83908 == 32'h0000_0003 ? add_83933 : array_index_83927[3];
  assign array_update_83935[4] = add_83908 == 32'h0000_0004 ? add_83933 : array_index_83927[4];
  assign array_update_83935[5] = add_83908 == 32'h0000_0005 ? add_83933 : array_index_83927[5];
  assign array_update_83935[6] = add_83908 == 32'h0000_0006 ? add_83933 : array_index_83927[6];
  assign array_update_83935[7] = add_83908 == 32'h0000_0007 ? add_83933 : array_index_83927[7];
  assign array_update_83935[8] = add_83908 == 32'h0000_0008 ? add_83933 : array_index_83927[8];
  assign array_update_83935[9] = add_83908 == 32'h0000_0009 ? add_83933 : array_index_83927[9];
  assign add_83936 = add_83923 + 32'h0000_0001;
  assign array_update_83937[0] = add_82825 == 32'h0000_0000 ? array_update_83935 : array_update_83924[0];
  assign array_update_83937[1] = add_82825 == 32'h0000_0001 ? array_update_83935 : array_update_83924[1];
  assign array_update_83937[2] = add_82825 == 32'h0000_0002 ? array_update_83935 : array_update_83924[2];
  assign array_update_83937[3] = add_82825 == 32'h0000_0003 ? array_update_83935 : array_update_83924[3];
  assign array_update_83937[4] = add_82825 == 32'h0000_0004 ? array_update_83935 : array_update_83924[4];
  assign array_update_83937[5] = add_82825 == 32'h0000_0005 ? array_update_83935 : array_update_83924[5];
  assign array_update_83937[6] = add_82825 == 32'h0000_0006 ? array_update_83935 : array_update_83924[6];
  assign array_update_83937[7] = add_82825 == 32'h0000_0007 ? array_update_83935 : array_update_83924[7];
  assign array_update_83937[8] = add_82825 == 32'h0000_0008 ? array_update_83935 : array_update_83924[8];
  assign array_update_83937[9] = add_82825 == 32'h0000_0009 ? array_update_83935 : array_update_83924[9];
  assign array_index_83939 = array_update_72021[add_83936 > 32'h0000_0009 ? 4'h9 : add_83936[3:0]];
  assign array_index_83940 = array_update_83937[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_83944 = smul32b_32b_x_32b(array_index_82832[add_83936 > 32'h0000_0009 ? 4'h9 : add_83936[3:0]], array_index_83939[add_83908 > 32'h0000_0009 ? 4'h9 : add_83908[3:0]]);
  assign add_83946 = array_index_83940[add_83908 > 32'h0000_0009 ? 4'h9 : add_83908[3:0]] + smul_83944;
  assign array_update_83948[0] = add_83908 == 32'h0000_0000 ? add_83946 : array_index_83940[0];
  assign array_update_83948[1] = add_83908 == 32'h0000_0001 ? add_83946 : array_index_83940[1];
  assign array_update_83948[2] = add_83908 == 32'h0000_0002 ? add_83946 : array_index_83940[2];
  assign array_update_83948[3] = add_83908 == 32'h0000_0003 ? add_83946 : array_index_83940[3];
  assign array_update_83948[4] = add_83908 == 32'h0000_0004 ? add_83946 : array_index_83940[4];
  assign array_update_83948[5] = add_83908 == 32'h0000_0005 ? add_83946 : array_index_83940[5];
  assign array_update_83948[6] = add_83908 == 32'h0000_0006 ? add_83946 : array_index_83940[6];
  assign array_update_83948[7] = add_83908 == 32'h0000_0007 ? add_83946 : array_index_83940[7];
  assign array_update_83948[8] = add_83908 == 32'h0000_0008 ? add_83946 : array_index_83940[8];
  assign array_update_83948[9] = add_83908 == 32'h0000_0009 ? add_83946 : array_index_83940[9];
  assign add_83949 = add_83936 + 32'h0000_0001;
  assign array_update_83950[0] = add_82825 == 32'h0000_0000 ? array_update_83948 : array_update_83937[0];
  assign array_update_83950[1] = add_82825 == 32'h0000_0001 ? array_update_83948 : array_update_83937[1];
  assign array_update_83950[2] = add_82825 == 32'h0000_0002 ? array_update_83948 : array_update_83937[2];
  assign array_update_83950[3] = add_82825 == 32'h0000_0003 ? array_update_83948 : array_update_83937[3];
  assign array_update_83950[4] = add_82825 == 32'h0000_0004 ? array_update_83948 : array_update_83937[4];
  assign array_update_83950[5] = add_82825 == 32'h0000_0005 ? array_update_83948 : array_update_83937[5];
  assign array_update_83950[6] = add_82825 == 32'h0000_0006 ? array_update_83948 : array_update_83937[6];
  assign array_update_83950[7] = add_82825 == 32'h0000_0007 ? array_update_83948 : array_update_83937[7];
  assign array_update_83950[8] = add_82825 == 32'h0000_0008 ? array_update_83948 : array_update_83937[8];
  assign array_update_83950[9] = add_82825 == 32'h0000_0009 ? array_update_83948 : array_update_83937[9];
  assign array_index_83952 = array_update_72021[add_83949 > 32'h0000_0009 ? 4'h9 : add_83949[3:0]];
  assign array_index_83953 = array_update_83950[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_83957 = smul32b_32b_x_32b(array_index_82832[add_83949 > 32'h0000_0009 ? 4'h9 : add_83949[3:0]], array_index_83952[add_83908 > 32'h0000_0009 ? 4'h9 : add_83908[3:0]]);
  assign add_83959 = array_index_83953[add_83908 > 32'h0000_0009 ? 4'h9 : add_83908[3:0]] + smul_83957;
  assign array_update_83961[0] = add_83908 == 32'h0000_0000 ? add_83959 : array_index_83953[0];
  assign array_update_83961[1] = add_83908 == 32'h0000_0001 ? add_83959 : array_index_83953[1];
  assign array_update_83961[2] = add_83908 == 32'h0000_0002 ? add_83959 : array_index_83953[2];
  assign array_update_83961[3] = add_83908 == 32'h0000_0003 ? add_83959 : array_index_83953[3];
  assign array_update_83961[4] = add_83908 == 32'h0000_0004 ? add_83959 : array_index_83953[4];
  assign array_update_83961[5] = add_83908 == 32'h0000_0005 ? add_83959 : array_index_83953[5];
  assign array_update_83961[6] = add_83908 == 32'h0000_0006 ? add_83959 : array_index_83953[6];
  assign array_update_83961[7] = add_83908 == 32'h0000_0007 ? add_83959 : array_index_83953[7];
  assign array_update_83961[8] = add_83908 == 32'h0000_0008 ? add_83959 : array_index_83953[8];
  assign array_update_83961[9] = add_83908 == 32'h0000_0009 ? add_83959 : array_index_83953[9];
  assign add_83962 = add_83949 + 32'h0000_0001;
  assign array_update_83963[0] = add_82825 == 32'h0000_0000 ? array_update_83961 : array_update_83950[0];
  assign array_update_83963[1] = add_82825 == 32'h0000_0001 ? array_update_83961 : array_update_83950[1];
  assign array_update_83963[2] = add_82825 == 32'h0000_0002 ? array_update_83961 : array_update_83950[2];
  assign array_update_83963[3] = add_82825 == 32'h0000_0003 ? array_update_83961 : array_update_83950[3];
  assign array_update_83963[4] = add_82825 == 32'h0000_0004 ? array_update_83961 : array_update_83950[4];
  assign array_update_83963[5] = add_82825 == 32'h0000_0005 ? array_update_83961 : array_update_83950[5];
  assign array_update_83963[6] = add_82825 == 32'h0000_0006 ? array_update_83961 : array_update_83950[6];
  assign array_update_83963[7] = add_82825 == 32'h0000_0007 ? array_update_83961 : array_update_83950[7];
  assign array_update_83963[8] = add_82825 == 32'h0000_0008 ? array_update_83961 : array_update_83950[8];
  assign array_update_83963[9] = add_82825 == 32'h0000_0009 ? array_update_83961 : array_update_83950[9];
  assign array_index_83965 = array_update_72021[add_83962 > 32'h0000_0009 ? 4'h9 : add_83962[3:0]];
  assign array_index_83966 = array_update_83963[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_83970 = smul32b_32b_x_32b(array_index_82832[add_83962 > 32'h0000_0009 ? 4'h9 : add_83962[3:0]], array_index_83965[add_83908 > 32'h0000_0009 ? 4'h9 : add_83908[3:0]]);
  assign add_83972 = array_index_83966[add_83908 > 32'h0000_0009 ? 4'h9 : add_83908[3:0]] + smul_83970;
  assign array_update_83974[0] = add_83908 == 32'h0000_0000 ? add_83972 : array_index_83966[0];
  assign array_update_83974[1] = add_83908 == 32'h0000_0001 ? add_83972 : array_index_83966[1];
  assign array_update_83974[2] = add_83908 == 32'h0000_0002 ? add_83972 : array_index_83966[2];
  assign array_update_83974[3] = add_83908 == 32'h0000_0003 ? add_83972 : array_index_83966[3];
  assign array_update_83974[4] = add_83908 == 32'h0000_0004 ? add_83972 : array_index_83966[4];
  assign array_update_83974[5] = add_83908 == 32'h0000_0005 ? add_83972 : array_index_83966[5];
  assign array_update_83974[6] = add_83908 == 32'h0000_0006 ? add_83972 : array_index_83966[6];
  assign array_update_83974[7] = add_83908 == 32'h0000_0007 ? add_83972 : array_index_83966[7];
  assign array_update_83974[8] = add_83908 == 32'h0000_0008 ? add_83972 : array_index_83966[8];
  assign array_update_83974[9] = add_83908 == 32'h0000_0009 ? add_83972 : array_index_83966[9];
  assign add_83975 = add_83962 + 32'h0000_0001;
  assign array_update_83976[0] = add_82825 == 32'h0000_0000 ? array_update_83974 : array_update_83963[0];
  assign array_update_83976[1] = add_82825 == 32'h0000_0001 ? array_update_83974 : array_update_83963[1];
  assign array_update_83976[2] = add_82825 == 32'h0000_0002 ? array_update_83974 : array_update_83963[2];
  assign array_update_83976[3] = add_82825 == 32'h0000_0003 ? array_update_83974 : array_update_83963[3];
  assign array_update_83976[4] = add_82825 == 32'h0000_0004 ? array_update_83974 : array_update_83963[4];
  assign array_update_83976[5] = add_82825 == 32'h0000_0005 ? array_update_83974 : array_update_83963[5];
  assign array_update_83976[6] = add_82825 == 32'h0000_0006 ? array_update_83974 : array_update_83963[6];
  assign array_update_83976[7] = add_82825 == 32'h0000_0007 ? array_update_83974 : array_update_83963[7];
  assign array_update_83976[8] = add_82825 == 32'h0000_0008 ? array_update_83974 : array_update_83963[8];
  assign array_update_83976[9] = add_82825 == 32'h0000_0009 ? array_update_83974 : array_update_83963[9];
  assign array_index_83978 = array_update_72021[add_83975 > 32'h0000_0009 ? 4'h9 : add_83975[3:0]];
  assign array_index_83979 = array_update_83976[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_83983 = smul32b_32b_x_32b(array_index_82832[add_83975 > 32'h0000_0009 ? 4'h9 : add_83975[3:0]], array_index_83978[add_83908 > 32'h0000_0009 ? 4'h9 : add_83908[3:0]]);
  assign add_83985 = array_index_83979[add_83908 > 32'h0000_0009 ? 4'h9 : add_83908[3:0]] + smul_83983;
  assign array_update_83987[0] = add_83908 == 32'h0000_0000 ? add_83985 : array_index_83979[0];
  assign array_update_83987[1] = add_83908 == 32'h0000_0001 ? add_83985 : array_index_83979[1];
  assign array_update_83987[2] = add_83908 == 32'h0000_0002 ? add_83985 : array_index_83979[2];
  assign array_update_83987[3] = add_83908 == 32'h0000_0003 ? add_83985 : array_index_83979[3];
  assign array_update_83987[4] = add_83908 == 32'h0000_0004 ? add_83985 : array_index_83979[4];
  assign array_update_83987[5] = add_83908 == 32'h0000_0005 ? add_83985 : array_index_83979[5];
  assign array_update_83987[6] = add_83908 == 32'h0000_0006 ? add_83985 : array_index_83979[6];
  assign array_update_83987[7] = add_83908 == 32'h0000_0007 ? add_83985 : array_index_83979[7];
  assign array_update_83987[8] = add_83908 == 32'h0000_0008 ? add_83985 : array_index_83979[8];
  assign array_update_83987[9] = add_83908 == 32'h0000_0009 ? add_83985 : array_index_83979[9];
  assign add_83988 = add_83975 + 32'h0000_0001;
  assign array_update_83989[0] = add_82825 == 32'h0000_0000 ? array_update_83987 : array_update_83976[0];
  assign array_update_83989[1] = add_82825 == 32'h0000_0001 ? array_update_83987 : array_update_83976[1];
  assign array_update_83989[2] = add_82825 == 32'h0000_0002 ? array_update_83987 : array_update_83976[2];
  assign array_update_83989[3] = add_82825 == 32'h0000_0003 ? array_update_83987 : array_update_83976[3];
  assign array_update_83989[4] = add_82825 == 32'h0000_0004 ? array_update_83987 : array_update_83976[4];
  assign array_update_83989[5] = add_82825 == 32'h0000_0005 ? array_update_83987 : array_update_83976[5];
  assign array_update_83989[6] = add_82825 == 32'h0000_0006 ? array_update_83987 : array_update_83976[6];
  assign array_update_83989[7] = add_82825 == 32'h0000_0007 ? array_update_83987 : array_update_83976[7];
  assign array_update_83989[8] = add_82825 == 32'h0000_0008 ? array_update_83987 : array_update_83976[8];
  assign array_update_83989[9] = add_82825 == 32'h0000_0009 ? array_update_83987 : array_update_83976[9];
  assign array_index_83991 = array_update_72021[add_83988 > 32'h0000_0009 ? 4'h9 : add_83988[3:0]];
  assign array_index_83992 = array_update_83989[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_83996 = smul32b_32b_x_32b(array_index_82832[add_83988 > 32'h0000_0009 ? 4'h9 : add_83988[3:0]], array_index_83991[add_83908 > 32'h0000_0009 ? 4'h9 : add_83908[3:0]]);
  assign add_83998 = array_index_83992[add_83908 > 32'h0000_0009 ? 4'h9 : add_83908[3:0]] + smul_83996;
  assign array_update_84000[0] = add_83908 == 32'h0000_0000 ? add_83998 : array_index_83992[0];
  assign array_update_84000[1] = add_83908 == 32'h0000_0001 ? add_83998 : array_index_83992[1];
  assign array_update_84000[2] = add_83908 == 32'h0000_0002 ? add_83998 : array_index_83992[2];
  assign array_update_84000[3] = add_83908 == 32'h0000_0003 ? add_83998 : array_index_83992[3];
  assign array_update_84000[4] = add_83908 == 32'h0000_0004 ? add_83998 : array_index_83992[4];
  assign array_update_84000[5] = add_83908 == 32'h0000_0005 ? add_83998 : array_index_83992[5];
  assign array_update_84000[6] = add_83908 == 32'h0000_0006 ? add_83998 : array_index_83992[6];
  assign array_update_84000[7] = add_83908 == 32'h0000_0007 ? add_83998 : array_index_83992[7];
  assign array_update_84000[8] = add_83908 == 32'h0000_0008 ? add_83998 : array_index_83992[8];
  assign array_update_84000[9] = add_83908 == 32'h0000_0009 ? add_83998 : array_index_83992[9];
  assign add_84001 = add_83988 + 32'h0000_0001;
  assign array_update_84002[0] = add_82825 == 32'h0000_0000 ? array_update_84000 : array_update_83989[0];
  assign array_update_84002[1] = add_82825 == 32'h0000_0001 ? array_update_84000 : array_update_83989[1];
  assign array_update_84002[2] = add_82825 == 32'h0000_0002 ? array_update_84000 : array_update_83989[2];
  assign array_update_84002[3] = add_82825 == 32'h0000_0003 ? array_update_84000 : array_update_83989[3];
  assign array_update_84002[4] = add_82825 == 32'h0000_0004 ? array_update_84000 : array_update_83989[4];
  assign array_update_84002[5] = add_82825 == 32'h0000_0005 ? array_update_84000 : array_update_83989[5];
  assign array_update_84002[6] = add_82825 == 32'h0000_0006 ? array_update_84000 : array_update_83989[6];
  assign array_update_84002[7] = add_82825 == 32'h0000_0007 ? array_update_84000 : array_update_83989[7];
  assign array_update_84002[8] = add_82825 == 32'h0000_0008 ? array_update_84000 : array_update_83989[8];
  assign array_update_84002[9] = add_82825 == 32'h0000_0009 ? array_update_84000 : array_update_83989[9];
  assign array_index_84004 = array_update_72021[add_84001 > 32'h0000_0009 ? 4'h9 : add_84001[3:0]];
  assign array_index_84005 = array_update_84002[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_84009 = smul32b_32b_x_32b(array_index_82832[add_84001 > 32'h0000_0009 ? 4'h9 : add_84001[3:0]], array_index_84004[add_83908 > 32'h0000_0009 ? 4'h9 : add_83908[3:0]]);
  assign add_84011 = array_index_84005[add_83908 > 32'h0000_0009 ? 4'h9 : add_83908[3:0]] + smul_84009;
  assign array_update_84013[0] = add_83908 == 32'h0000_0000 ? add_84011 : array_index_84005[0];
  assign array_update_84013[1] = add_83908 == 32'h0000_0001 ? add_84011 : array_index_84005[1];
  assign array_update_84013[2] = add_83908 == 32'h0000_0002 ? add_84011 : array_index_84005[2];
  assign array_update_84013[3] = add_83908 == 32'h0000_0003 ? add_84011 : array_index_84005[3];
  assign array_update_84013[4] = add_83908 == 32'h0000_0004 ? add_84011 : array_index_84005[4];
  assign array_update_84013[5] = add_83908 == 32'h0000_0005 ? add_84011 : array_index_84005[5];
  assign array_update_84013[6] = add_83908 == 32'h0000_0006 ? add_84011 : array_index_84005[6];
  assign array_update_84013[7] = add_83908 == 32'h0000_0007 ? add_84011 : array_index_84005[7];
  assign array_update_84013[8] = add_83908 == 32'h0000_0008 ? add_84011 : array_index_84005[8];
  assign array_update_84013[9] = add_83908 == 32'h0000_0009 ? add_84011 : array_index_84005[9];
  assign add_84014 = add_84001 + 32'h0000_0001;
  assign array_update_84015[0] = add_82825 == 32'h0000_0000 ? array_update_84013 : array_update_84002[0];
  assign array_update_84015[1] = add_82825 == 32'h0000_0001 ? array_update_84013 : array_update_84002[1];
  assign array_update_84015[2] = add_82825 == 32'h0000_0002 ? array_update_84013 : array_update_84002[2];
  assign array_update_84015[3] = add_82825 == 32'h0000_0003 ? array_update_84013 : array_update_84002[3];
  assign array_update_84015[4] = add_82825 == 32'h0000_0004 ? array_update_84013 : array_update_84002[4];
  assign array_update_84015[5] = add_82825 == 32'h0000_0005 ? array_update_84013 : array_update_84002[5];
  assign array_update_84015[6] = add_82825 == 32'h0000_0006 ? array_update_84013 : array_update_84002[6];
  assign array_update_84015[7] = add_82825 == 32'h0000_0007 ? array_update_84013 : array_update_84002[7];
  assign array_update_84015[8] = add_82825 == 32'h0000_0008 ? array_update_84013 : array_update_84002[8];
  assign array_update_84015[9] = add_82825 == 32'h0000_0009 ? array_update_84013 : array_update_84002[9];
  assign array_index_84017 = array_update_72021[add_84014 > 32'h0000_0009 ? 4'h9 : add_84014[3:0]];
  assign array_index_84018 = array_update_84015[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_84022 = smul32b_32b_x_32b(array_index_82832[add_84014 > 32'h0000_0009 ? 4'h9 : add_84014[3:0]], array_index_84017[add_83908 > 32'h0000_0009 ? 4'h9 : add_83908[3:0]]);
  assign add_84024 = array_index_84018[add_83908 > 32'h0000_0009 ? 4'h9 : add_83908[3:0]] + smul_84022;
  assign array_update_84026[0] = add_83908 == 32'h0000_0000 ? add_84024 : array_index_84018[0];
  assign array_update_84026[1] = add_83908 == 32'h0000_0001 ? add_84024 : array_index_84018[1];
  assign array_update_84026[2] = add_83908 == 32'h0000_0002 ? add_84024 : array_index_84018[2];
  assign array_update_84026[3] = add_83908 == 32'h0000_0003 ? add_84024 : array_index_84018[3];
  assign array_update_84026[4] = add_83908 == 32'h0000_0004 ? add_84024 : array_index_84018[4];
  assign array_update_84026[5] = add_83908 == 32'h0000_0005 ? add_84024 : array_index_84018[5];
  assign array_update_84026[6] = add_83908 == 32'h0000_0006 ? add_84024 : array_index_84018[6];
  assign array_update_84026[7] = add_83908 == 32'h0000_0007 ? add_84024 : array_index_84018[7];
  assign array_update_84026[8] = add_83908 == 32'h0000_0008 ? add_84024 : array_index_84018[8];
  assign array_update_84026[9] = add_83908 == 32'h0000_0009 ? add_84024 : array_index_84018[9];
  assign add_84027 = add_84014 + 32'h0000_0001;
  assign array_update_84028[0] = add_82825 == 32'h0000_0000 ? array_update_84026 : array_update_84015[0];
  assign array_update_84028[1] = add_82825 == 32'h0000_0001 ? array_update_84026 : array_update_84015[1];
  assign array_update_84028[2] = add_82825 == 32'h0000_0002 ? array_update_84026 : array_update_84015[2];
  assign array_update_84028[3] = add_82825 == 32'h0000_0003 ? array_update_84026 : array_update_84015[3];
  assign array_update_84028[4] = add_82825 == 32'h0000_0004 ? array_update_84026 : array_update_84015[4];
  assign array_update_84028[5] = add_82825 == 32'h0000_0005 ? array_update_84026 : array_update_84015[5];
  assign array_update_84028[6] = add_82825 == 32'h0000_0006 ? array_update_84026 : array_update_84015[6];
  assign array_update_84028[7] = add_82825 == 32'h0000_0007 ? array_update_84026 : array_update_84015[7];
  assign array_update_84028[8] = add_82825 == 32'h0000_0008 ? array_update_84026 : array_update_84015[8];
  assign array_update_84028[9] = add_82825 == 32'h0000_0009 ? array_update_84026 : array_update_84015[9];
  assign array_index_84030 = array_update_72021[add_84027 > 32'h0000_0009 ? 4'h9 : add_84027[3:0]];
  assign array_index_84031 = array_update_84028[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_84035 = smul32b_32b_x_32b(array_index_82832[add_84027 > 32'h0000_0009 ? 4'h9 : add_84027[3:0]], array_index_84030[add_83908 > 32'h0000_0009 ? 4'h9 : add_83908[3:0]]);
  assign add_84037 = array_index_84031[add_83908 > 32'h0000_0009 ? 4'h9 : add_83908[3:0]] + smul_84035;
  assign array_update_84038[0] = add_83908 == 32'h0000_0000 ? add_84037 : array_index_84031[0];
  assign array_update_84038[1] = add_83908 == 32'h0000_0001 ? add_84037 : array_index_84031[1];
  assign array_update_84038[2] = add_83908 == 32'h0000_0002 ? add_84037 : array_index_84031[2];
  assign array_update_84038[3] = add_83908 == 32'h0000_0003 ? add_84037 : array_index_84031[3];
  assign array_update_84038[4] = add_83908 == 32'h0000_0004 ? add_84037 : array_index_84031[4];
  assign array_update_84038[5] = add_83908 == 32'h0000_0005 ? add_84037 : array_index_84031[5];
  assign array_update_84038[6] = add_83908 == 32'h0000_0006 ? add_84037 : array_index_84031[6];
  assign array_update_84038[7] = add_83908 == 32'h0000_0007 ? add_84037 : array_index_84031[7];
  assign array_update_84038[8] = add_83908 == 32'h0000_0008 ? add_84037 : array_index_84031[8];
  assign array_update_84038[9] = add_83908 == 32'h0000_0009 ? add_84037 : array_index_84031[9];
  assign array_update_84039[0] = add_82825 == 32'h0000_0000 ? array_update_84038 : array_update_84028[0];
  assign array_update_84039[1] = add_82825 == 32'h0000_0001 ? array_update_84038 : array_update_84028[1];
  assign array_update_84039[2] = add_82825 == 32'h0000_0002 ? array_update_84038 : array_update_84028[2];
  assign array_update_84039[3] = add_82825 == 32'h0000_0003 ? array_update_84038 : array_update_84028[3];
  assign array_update_84039[4] = add_82825 == 32'h0000_0004 ? array_update_84038 : array_update_84028[4];
  assign array_update_84039[5] = add_82825 == 32'h0000_0005 ? array_update_84038 : array_update_84028[5];
  assign array_update_84039[6] = add_82825 == 32'h0000_0006 ? array_update_84038 : array_update_84028[6];
  assign array_update_84039[7] = add_82825 == 32'h0000_0007 ? array_update_84038 : array_update_84028[7];
  assign array_update_84039[8] = add_82825 == 32'h0000_0008 ? array_update_84038 : array_update_84028[8];
  assign array_update_84039[9] = add_82825 == 32'h0000_0009 ? array_update_84038 : array_update_84028[9];
  assign array_index_84041 = array_update_84039[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign add_84043 = add_83908 + 32'h0000_0001;
  assign array_update_84044[0] = add_84043 == 32'h0000_0000 ? 32'h0000_0000 : array_index_84041[0];
  assign array_update_84044[1] = add_84043 == 32'h0000_0001 ? 32'h0000_0000 : array_index_84041[1];
  assign array_update_84044[2] = add_84043 == 32'h0000_0002 ? 32'h0000_0000 : array_index_84041[2];
  assign array_update_84044[3] = add_84043 == 32'h0000_0003 ? 32'h0000_0000 : array_index_84041[3];
  assign array_update_84044[4] = add_84043 == 32'h0000_0004 ? 32'h0000_0000 : array_index_84041[4];
  assign array_update_84044[5] = add_84043 == 32'h0000_0005 ? 32'h0000_0000 : array_index_84041[5];
  assign array_update_84044[6] = add_84043 == 32'h0000_0006 ? 32'h0000_0000 : array_index_84041[6];
  assign array_update_84044[7] = add_84043 == 32'h0000_0007 ? 32'h0000_0000 : array_index_84041[7];
  assign array_update_84044[8] = add_84043 == 32'h0000_0008 ? 32'h0000_0000 : array_index_84041[8];
  assign array_update_84044[9] = add_84043 == 32'h0000_0009 ? 32'h0000_0000 : array_index_84041[9];
  assign literal_84045 = 32'h0000_0000;
  assign array_update_84046[0] = add_82825 == 32'h0000_0000 ? array_update_84044 : array_update_84039[0];
  assign array_update_84046[1] = add_82825 == 32'h0000_0001 ? array_update_84044 : array_update_84039[1];
  assign array_update_84046[2] = add_82825 == 32'h0000_0002 ? array_update_84044 : array_update_84039[2];
  assign array_update_84046[3] = add_82825 == 32'h0000_0003 ? array_update_84044 : array_update_84039[3];
  assign array_update_84046[4] = add_82825 == 32'h0000_0004 ? array_update_84044 : array_update_84039[4];
  assign array_update_84046[5] = add_82825 == 32'h0000_0005 ? array_update_84044 : array_update_84039[5];
  assign array_update_84046[6] = add_82825 == 32'h0000_0006 ? array_update_84044 : array_update_84039[6];
  assign array_update_84046[7] = add_82825 == 32'h0000_0007 ? array_update_84044 : array_update_84039[7];
  assign array_update_84046[8] = add_82825 == 32'h0000_0008 ? array_update_84044 : array_update_84039[8];
  assign array_update_84046[9] = add_82825 == 32'h0000_0009 ? array_update_84044 : array_update_84039[9];
  assign array_index_84048 = array_update_72021[literal_84045 > 32'h0000_0009 ? 4'h9 : literal_84045[3:0]];
  assign array_index_84049 = array_update_84046[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_84053 = smul32b_32b_x_32b(array_index_82832[literal_84045 > 32'h0000_0009 ? 4'h9 : literal_84045[3:0]], array_index_84048[add_84043 > 32'h0000_0009 ? 4'h9 : add_84043[3:0]]);
  assign add_84055 = array_index_84049[add_84043 > 32'h0000_0009 ? 4'h9 : add_84043[3:0]] + smul_84053;
  assign array_update_84057[0] = add_84043 == 32'h0000_0000 ? add_84055 : array_index_84049[0];
  assign array_update_84057[1] = add_84043 == 32'h0000_0001 ? add_84055 : array_index_84049[1];
  assign array_update_84057[2] = add_84043 == 32'h0000_0002 ? add_84055 : array_index_84049[2];
  assign array_update_84057[3] = add_84043 == 32'h0000_0003 ? add_84055 : array_index_84049[3];
  assign array_update_84057[4] = add_84043 == 32'h0000_0004 ? add_84055 : array_index_84049[4];
  assign array_update_84057[5] = add_84043 == 32'h0000_0005 ? add_84055 : array_index_84049[5];
  assign array_update_84057[6] = add_84043 == 32'h0000_0006 ? add_84055 : array_index_84049[6];
  assign array_update_84057[7] = add_84043 == 32'h0000_0007 ? add_84055 : array_index_84049[7];
  assign array_update_84057[8] = add_84043 == 32'h0000_0008 ? add_84055 : array_index_84049[8];
  assign array_update_84057[9] = add_84043 == 32'h0000_0009 ? add_84055 : array_index_84049[9];
  assign add_84058 = literal_84045 + 32'h0000_0001;
  assign array_update_84059[0] = add_82825 == 32'h0000_0000 ? array_update_84057 : array_update_84046[0];
  assign array_update_84059[1] = add_82825 == 32'h0000_0001 ? array_update_84057 : array_update_84046[1];
  assign array_update_84059[2] = add_82825 == 32'h0000_0002 ? array_update_84057 : array_update_84046[2];
  assign array_update_84059[3] = add_82825 == 32'h0000_0003 ? array_update_84057 : array_update_84046[3];
  assign array_update_84059[4] = add_82825 == 32'h0000_0004 ? array_update_84057 : array_update_84046[4];
  assign array_update_84059[5] = add_82825 == 32'h0000_0005 ? array_update_84057 : array_update_84046[5];
  assign array_update_84059[6] = add_82825 == 32'h0000_0006 ? array_update_84057 : array_update_84046[6];
  assign array_update_84059[7] = add_82825 == 32'h0000_0007 ? array_update_84057 : array_update_84046[7];
  assign array_update_84059[8] = add_82825 == 32'h0000_0008 ? array_update_84057 : array_update_84046[8];
  assign array_update_84059[9] = add_82825 == 32'h0000_0009 ? array_update_84057 : array_update_84046[9];
  assign array_index_84061 = array_update_72021[add_84058 > 32'h0000_0009 ? 4'h9 : add_84058[3:0]];
  assign array_index_84062 = array_update_84059[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_84066 = smul32b_32b_x_32b(array_index_82832[add_84058 > 32'h0000_0009 ? 4'h9 : add_84058[3:0]], array_index_84061[add_84043 > 32'h0000_0009 ? 4'h9 : add_84043[3:0]]);
  assign add_84068 = array_index_84062[add_84043 > 32'h0000_0009 ? 4'h9 : add_84043[3:0]] + smul_84066;
  assign array_update_84070[0] = add_84043 == 32'h0000_0000 ? add_84068 : array_index_84062[0];
  assign array_update_84070[1] = add_84043 == 32'h0000_0001 ? add_84068 : array_index_84062[1];
  assign array_update_84070[2] = add_84043 == 32'h0000_0002 ? add_84068 : array_index_84062[2];
  assign array_update_84070[3] = add_84043 == 32'h0000_0003 ? add_84068 : array_index_84062[3];
  assign array_update_84070[4] = add_84043 == 32'h0000_0004 ? add_84068 : array_index_84062[4];
  assign array_update_84070[5] = add_84043 == 32'h0000_0005 ? add_84068 : array_index_84062[5];
  assign array_update_84070[6] = add_84043 == 32'h0000_0006 ? add_84068 : array_index_84062[6];
  assign array_update_84070[7] = add_84043 == 32'h0000_0007 ? add_84068 : array_index_84062[7];
  assign array_update_84070[8] = add_84043 == 32'h0000_0008 ? add_84068 : array_index_84062[8];
  assign array_update_84070[9] = add_84043 == 32'h0000_0009 ? add_84068 : array_index_84062[9];
  assign add_84071 = add_84058 + 32'h0000_0001;
  assign array_update_84072[0] = add_82825 == 32'h0000_0000 ? array_update_84070 : array_update_84059[0];
  assign array_update_84072[1] = add_82825 == 32'h0000_0001 ? array_update_84070 : array_update_84059[1];
  assign array_update_84072[2] = add_82825 == 32'h0000_0002 ? array_update_84070 : array_update_84059[2];
  assign array_update_84072[3] = add_82825 == 32'h0000_0003 ? array_update_84070 : array_update_84059[3];
  assign array_update_84072[4] = add_82825 == 32'h0000_0004 ? array_update_84070 : array_update_84059[4];
  assign array_update_84072[5] = add_82825 == 32'h0000_0005 ? array_update_84070 : array_update_84059[5];
  assign array_update_84072[6] = add_82825 == 32'h0000_0006 ? array_update_84070 : array_update_84059[6];
  assign array_update_84072[7] = add_82825 == 32'h0000_0007 ? array_update_84070 : array_update_84059[7];
  assign array_update_84072[8] = add_82825 == 32'h0000_0008 ? array_update_84070 : array_update_84059[8];
  assign array_update_84072[9] = add_82825 == 32'h0000_0009 ? array_update_84070 : array_update_84059[9];
  assign array_index_84074 = array_update_72021[add_84071 > 32'h0000_0009 ? 4'h9 : add_84071[3:0]];
  assign array_index_84075 = array_update_84072[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_84079 = smul32b_32b_x_32b(array_index_82832[add_84071 > 32'h0000_0009 ? 4'h9 : add_84071[3:0]], array_index_84074[add_84043 > 32'h0000_0009 ? 4'h9 : add_84043[3:0]]);
  assign add_84081 = array_index_84075[add_84043 > 32'h0000_0009 ? 4'h9 : add_84043[3:0]] + smul_84079;
  assign array_update_84083[0] = add_84043 == 32'h0000_0000 ? add_84081 : array_index_84075[0];
  assign array_update_84083[1] = add_84043 == 32'h0000_0001 ? add_84081 : array_index_84075[1];
  assign array_update_84083[2] = add_84043 == 32'h0000_0002 ? add_84081 : array_index_84075[2];
  assign array_update_84083[3] = add_84043 == 32'h0000_0003 ? add_84081 : array_index_84075[3];
  assign array_update_84083[4] = add_84043 == 32'h0000_0004 ? add_84081 : array_index_84075[4];
  assign array_update_84083[5] = add_84043 == 32'h0000_0005 ? add_84081 : array_index_84075[5];
  assign array_update_84083[6] = add_84043 == 32'h0000_0006 ? add_84081 : array_index_84075[6];
  assign array_update_84083[7] = add_84043 == 32'h0000_0007 ? add_84081 : array_index_84075[7];
  assign array_update_84083[8] = add_84043 == 32'h0000_0008 ? add_84081 : array_index_84075[8];
  assign array_update_84083[9] = add_84043 == 32'h0000_0009 ? add_84081 : array_index_84075[9];
  assign add_84084 = add_84071 + 32'h0000_0001;
  assign array_update_84085[0] = add_82825 == 32'h0000_0000 ? array_update_84083 : array_update_84072[0];
  assign array_update_84085[1] = add_82825 == 32'h0000_0001 ? array_update_84083 : array_update_84072[1];
  assign array_update_84085[2] = add_82825 == 32'h0000_0002 ? array_update_84083 : array_update_84072[2];
  assign array_update_84085[3] = add_82825 == 32'h0000_0003 ? array_update_84083 : array_update_84072[3];
  assign array_update_84085[4] = add_82825 == 32'h0000_0004 ? array_update_84083 : array_update_84072[4];
  assign array_update_84085[5] = add_82825 == 32'h0000_0005 ? array_update_84083 : array_update_84072[5];
  assign array_update_84085[6] = add_82825 == 32'h0000_0006 ? array_update_84083 : array_update_84072[6];
  assign array_update_84085[7] = add_82825 == 32'h0000_0007 ? array_update_84083 : array_update_84072[7];
  assign array_update_84085[8] = add_82825 == 32'h0000_0008 ? array_update_84083 : array_update_84072[8];
  assign array_update_84085[9] = add_82825 == 32'h0000_0009 ? array_update_84083 : array_update_84072[9];
  assign array_index_84087 = array_update_72021[add_84084 > 32'h0000_0009 ? 4'h9 : add_84084[3:0]];
  assign array_index_84088 = array_update_84085[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_84092 = smul32b_32b_x_32b(array_index_82832[add_84084 > 32'h0000_0009 ? 4'h9 : add_84084[3:0]], array_index_84087[add_84043 > 32'h0000_0009 ? 4'h9 : add_84043[3:0]]);
  assign add_84094 = array_index_84088[add_84043 > 32'h0000_0009 ? 4'h9 : add_84043[3:0]] + smul_84092;
  assign array_update_84096[0] = add_84043 == 32'h0000_0000 ? add_84094 : array_index_84088[0];
  assign array_update_84096[1] = add_84043 == 32'h0000_0001 ? add_84094 : array_index_84088[1];
  assign array_update_84096[2] = add_84043 == 32'h0000_0002 ? add_84094 : array_index_84088[2];
  assign array_update_84096[3] = add_84043 == 32'h0000_0003 ? add_84094 : array_index_84088[3];
  assign array_update_84096[4] = add_84043 == 32'h0000_0004 ? add_84094 : array_index_84088[4];
  assign array_update_84096[5] = add_84043 == 32'h0000_0005 ? add_84094 : array_index_84088[5];
  assign array_update_84096[6] = add_84043 == 32'h0000_0006 ? add_84094 : array_index_84088[6];
  assign array_update_84096[7] = add_84043 == 32'h0000_0007 ? add_84094 : array_index_84088[7];
  assign array_update_84096[8] = add_84043 == 32'h0000_0008 ? add_84094 : array_index_84088[8];
  assign array_update_84096[9] = add_84043 == 32'h0000_0009 ? add_84094 : array_index_84088[9];
  assign add_84097 = add_84084 + 32'h0000_0001;
  assign array_update_84098[0] = add_82825 == 32'h0000_0000 ? array_update_84096 : array_update_84085[0];
  assign array_update_84098[1] = add_82825 == 32'h0000_0001 ? array_update_84096 : array_update_84085[1];
  assign array_update_84098[2] = add_82825 == 32'h0000_0002 ? array_update_84096 : array_update_84085[2];
  assign array_update_84098[3] = add_82825 == 32'h0000_0003 ? array_update_84096 : array_update_84085[3];
  assign array_update_84098[4] = add_82825 == 32'h0000_0004 ? array_update_84096 : array_update_84085[4];
  assign array_update_84098[5] = add_82825 == 32'h0000_0005 ? array_update_84096 : array_update_84085[5];
  assign array_update_84098[6] = add_82825 == 32'h0000_0006 ? array_update_84096 : array_update_84085[6];
  assign array_update_84098[7] = add_82825 == 32'h0000_0007 ? array_update_84096 : array_update_84085[7];
  assign array_update_84098[8] = add_82825 == 32'h0000_0008 ? array_update_84096 : array_update_84085[8];
  assign array_update_84098[9] = add_82825 == 32'h0000_0009 ? array_update_84096 : array_update_84085[9];
  assign array_index_84100 = array_update_72021[add_84097 > 32'h0000_0009 ? 4'h9 : add_84097[3:0]];
  assign array_index_84101 = array_update_84098[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_84105 = smul32b_32b_x_32b(array_index_82832[add_84097 > 32'h0000_0009 ? 4'h9 : add_84097[3:0]], array_index_84100[add_84043 > 32'h0000_0009 ? 4'h9 : add_84043[3:0]]);
  assign add_84107 = array_index_84101[add_84043 > 32'h0000_0009 ? 4'h9 : add_84043[3:0]] + smul_84105;
  assign array_update_84109[0] = add_84043 == 32'h0000_0000 ? add_84107 : array_index_84101[0];
  assign array_update_84109[1] = add_84043 == 32'h0000_0001 ? add_84107 : array_index_84101[1];
  assign array_update_84109[2] = add_84043 == 32'h0000_0002 ? add_84107 : array_index_84101[2];
  assign array_update_84109[3] = add_84043 == 32'h0000_0003 ? add_84107 : array_index_84101[3];
  assign array_update_84109[4] = add_84043 == 32'h0000_0004 ? add_84107 : array_index_84101[4];
  assign array_update_84109[5] = add_84043 == 32'h0000_0005 ? add_84107 : array_index_84101[5];
  assign array_update_84109[6] = add_84043 == 32'h0000_0006 ? add_84107 : array_index_84101[6];
  assign array_update_84109[7] = add_84043 == 32'h0000_0007 ? add_84107 : array_index_84101[7];
  assign array_update_84109[8] = add_84043 == 32'h0000_0008 ? add_84107 : array_index_84101[8];
  assign array_update_84109[9] = add_84043 == 32'h0000_0009 ? add_84107 : array_index_84101[9];
  assign add_84110 = add_84097 + 32'h0000_0001;
  assign array_update_84111[0] = add_82825 == 32'h0000_0000 ? array_update_84109 : array_update_84098[0];
  assign array_update_84111[1] = add_82825 == 32'h0000_0001 ? array_update_84109 : array_update_84098[1];
  assign array_update_84111[2] = add_82825 == 32'h0000_0002 ? array_update_84109 : array_update_84098[2];
  assign array_update_84111[3] = add_82825 == 32'h0000_0003 ? array_update_84109 : array_update_84098[3];
  assign array_update_84111[4] = add_82825 == 32'h0000_0004 ? array_update_84109 : array_update_84098[4];
  assign array_update_84111[5] = add_82825 == 32'h0000_0005 ? array_update_84109 : array_update_84098[5];
  assign array_update_84111[6] = add_82825 == 32'h0000_0006 ? array_update_84109 : array_update_84098[6];
  assign array_update_84111[7] = add_82825 == 32'h0000_0007 ? array_update_84109 : array_update_84098[7];
  assign array_update_84111[8] = add_82825 == 32'h0000_0008 ? array_update_84109 : array_update_84098[8];
  assign array_update_84111[9] = add_82825 == 32'h0000_0009 ? array_update_84109 : array_update_84098[9];
  assign array_index_84113 = array_update_72021[add_84110 > 32'h0000_0009 ? 4'h9 : add_84110[3:0]];
  assign array_index_84114 = array_update_84111[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_84118 = smul32b_32b_x_32b(array_index_82832[add_84110 > 32'h0000_0009 ? 4'h9 : add_84110[3:0]], array_index_84113[add_84043 > 32'h0000_0009 ? 4'h9 : add_84043[3:0]]);
  assign add_84120 = array_index_84114[add_84043 > 32'h0000_0009 ? 4'h9 : add_84043[3:0]] + smul_84118;
  assign array_update_84122[0] = add_84043 == 32'h0000_0000 ? add_84120 : array_index_84114[0];
  assign array_update_84122[1] = add_84043 == 32'h0000_0001 ? add_84120 : array_index_84114[1];
  assign array_update_84122[2] = add_84043 == 32'h0000_0002 ? add_84120 : array_index_84114[2];
  assign array_update_84122[3] = add_84043 == 32'h0000_0003 ? add_84120 : array_index_84114[3];
  assign array_update_84122[4] = add_84043 == 32'h0000_0004 ? add_84120 : array_index_84114[4];
  assign array_update_84122[5] = add_84043 == 32'h0000_0005 ? add_84120 : array_index_84114[5];
  assign array_update_84122[6] = add_84043 == 32'h0000_0006 ? add_84120 : array_index_84114[6];
  assign array_update_84122[7] = add_84043 == 32'h0000_0007 ? add_84120 : array_index_84114[7];
  assign array_update_84122[8] = add_84043 == 32'h0000_0008 ? add_84120 : array_index_84114[8];
  assign array_update_84122[9] = add_84043 == 32'h0000_0009 ? add_84120 : array_index_84114[9];
  assign add_84123 = add_84110 + 32'h0000_0001;
  assign array_update_84124[0] = add_82825 == 32'h0000_0000 ? array_update_84122 : array_update_84111[0];
  assign array_update_84124[1] = add_82825 == 32'h0000_0001 ? array_update_84122 : array_update_84111[1];
  assign array_update_84124[2] = add_82825 == 32'h0000_0002 ? array_update_84122 : array_update_84111[2];
  assign array_update_84124[3] = add_82825 == 32'h0000_0003 ? array_update_84122 : array_update_84111[3];
  assign array_update_84124[4] = add_82825 == 32'h0000_0004 ? array_update_84122 : array_update_84111[4];
  assign array_update_84124[5] = add_82825 == 32'h0000_0005 ? array_update_84122 : array_update_84111[5];
  assign array_update_84124[6] = add_82825 == 32'h0000_0006 ? array_update_84122 : array_update_84111[6];
  assign array_update_84124[7] = add_82825 == 32'h0000_0007 ? array_update_84122 : array_update_84111[7];
  assign array_update_84124[8] = add_82825 == 32'h0000_0008 ? array_update_84122 : array_update_84111[8];
  assign array_update_84124[9] = add_82825 == 32'h0000_0009 ? array_update_84122 : array_update_84111[9];
  assign array_index_84126 = array_update_72021[add_84123 > 32'h0000_0009 ? 4'h9 : add_84123[3:0]];
  assign array_index_84127 = array_update_84124[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_84131 = smul32b_32b_x_32b(array_index_82832[add_84123 > 32'h0000_0009 ? 4'h9 : add_84123[3:0]], array_index_84126[add_84043 > 32'h0000_0009 ? 4'h9 : add_84043[3:0]]);
  assign add_84133 = array_index_84127[add_84043 > 32'h0000_0009 ? 4'h9 : add_84043[3:0]] + smul_84131;
  assign array_update_84135[0] = add_84043 == 32'h0000_0000 ? add_84133 : array_index_84127[0];
  assign array_update_84135[1] = add_84043 == 32'h0000_0001 ? add_84133 : array_index_84127[1];
  assign array_update_84135[2] = add_84043 == 32'h0000_0002 ? add_84133 : array_index_84127[2];
  assign array_update_84135[3] = add_84043 == 32'h0000_0003 ? add_84133 : array_index_84127[3];
  assign array_update_84135[4] = add_84043 == 32'h0000_0004 ? add_84133 : array_index_84127[4];
  assign array_update_84135[5] = add_84043 == 32'h0000_0005 ? add_84133 : array_index_84127[5];
  assign array_update_84135[6] = add_84043 == 32'h0000_0006 ? add_84133 : array_index_84127[6];
  assign array_update_84135[7] = add_84043 == 32'h0000_0007 ? add_84133 : array_index_84127[7];
  assign array_update_84135[8] = add_84043 == 32'h0000_0008 ? add_84133 : array_index_84127[8];
  assign array_update_84135[9] = add_84043 == 32'h0000_0009 ? add_84133 : array_index_84127[9];
  assign add_84136 = add_84123 + 32'h0000_0001;
  assign array_update_84137[0] = add_82825 == 32'h0000_0000 ? array_update_84135 : array_update_84124[0];
  assign array_update_84137[1] = add_82825 == 32'h0000_0001 ? array_update_84135 : array_update_84124[1];
  assign array_update_84137[2] = add_82825 == 32'h0000_0002 ? array_update_84135 : array_update_84124[2];
  assign array_update_84137[3] = add_82825 == 32'h0000_0003 ? array_update_84135 : array_update_84124[3];
  assign array_update_84137[4] = add_82825 == 32'h0000_0004 ? array_update_84135 : array_update_84124[4];
  assign array_update_84137[5] = add_82825 == 32'h0000_0005 ? array_update_84135 : array_update_84124[5];
  assign array_update_84137[6] = add_82825 == 32'h0000_0006 ? array_update_84135 : array_update_84124[6];
  assign array_update_84137[7] = add_82825 == 32'h0000_0007 ? array_update_84135 : array_update_84124[7];
  assign array_update_84137[8] = add_82825 == 32'h0000_0008 ? array_update_84135 : array_update_84124[8];
  assign array_update_84137[9] = add_82825 == 32'h0000_0009 ? array_update_84135 : array_update_84124[9];
  assign array_index_84139 = array_update_72021[add_84136 > 32'h0000_0009 ? 4'h9 : add_84136[3:0]];
  assign array_index_84140 = array_update_84137[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_84144 = smul32b_32b_x_32b(array_index_82832[add_84136 > 32'h0000_0009 ? 4'h9 : add_84136[3:0]], array_index_84139[add_84043 > 32'h0000_0009 ? 4'h9 : add_84043[3:0]]);
  assign add_84146 = array_index_84140[add_84043 > 32'h0000_0009 ? 4'h9 : add_84043[3:0]] + smul_84144;
  assign array_update_84148[0] = add_84043 == 32'h0000_0000 ? add_84146 : array_index_84140[0];
  assign array_update_84148[1] = add_84043 == 32'h0000_0001 ? add_84146 : array_index_84140[1];
  assign array_update_84148[2] = add_84043 == 32'h0000_0002 ? add_84146 : array_index_84140[2];
  assign array_update_84148[3] = add_84043 == 32'h0000_0003 ? add_84146 : array_index_84140[3];
  assign array_update_84148[4] = add_84043 == 32'h0000_0004 ? add_84146 : array_index_84140[4];
  assign array_update_84148[5] = add_84043 == 32'h0000_0005 ? add_84146 : array_index_84140[5];
  assign array_update_84148[6] = add_84043 == 32'h0000_0006 ? add_84146 : array_index_84140[6];
  assign array_update_84148[7] = add_84043 == 32'h0000_0007 ? add_84146 : array_index_84140[7];
  assign array_update_84148[8] = add_84043 == 32'h0000_0008 ? add_84146 : array_index_84140[8];
  assign array_update_84148[9] = add_84043 == 32'h0000_0009 ? add_84146 : array_index_84140[9];
  assign add_84149 = add_84136 + 32'h0000_0001;
  assign array_update_84150[0] = add_82825 == 32'h0000_0000 ? array_update_84148 : array_update_84137[0];
  assign array_update_84150[1] = add_82825 == 32'h0000_0001 ? array_update_84148 : array_update_84137[1];
  assign array_update_84150[2] = add_82825 == 32'h0000_0002 ? array_update_84148 : array_update_84137[2];
  assign array_update_84150[3] = add_82825 == 32'h0000_0003 ? array_update_84148 : array_update_84137[3];
  assign array_update_84150[4] = add_82825 == 32'h0000_0004 ? array_update_84148 : array_update_84137[4];
  assign array_update_84150[5] = add_82825 == 32'h0000_0005 ? array_update_84148 : array_update_84137[5];
  assign array_update_84150[6] = add_82825 == 32'h0000_0006 ? array_update_84148 : array_update_84137[6];
  assign array_update_84150[7] = add_82825 == 32'h0000_0007 ? array_update_84148 : array_update_84137[7];
  assign array_update_84150[8] = add_82825 == 32'h0000_0008 ? array_update_84148 : array_update_84137[8];
  assign array_update_84150[9] = add_82825 == 32'h0000_0009 ? array_update_84148 : array_update_84137[9];
  assign array_index_84152 = array_update_72021[add_84149 > 32'h0000_0009 ? 4'h9 : add_84149[3:0]];
  assign array_index_84153 = array_update_84150[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_84157 = smul32b_32b_x_32b(array_index_82832[add_84149 > 32'h0000_0009 ? 4'h9 : add_84149[3:0]], array_index_84152[add_84043 > 32'h0000_0009 ? 4'h9 : add_84043[3:0]]);
  assign add_84159 = array_index_84153[add_84043 > 32'h0000_0009 ? 4'h9 : add_84043[3:0]] + smul_84157;
  assign array_update_84161[0] = add_84043 == 32'h0000_0000 ? add_84159 : array_index_84153[0];
  assign array_update_84161[1] = add_84043 == 32'h0000_0001 ? add_84159 : array_index_84153[1];
  assign array_update_84161[2] = add_84043 == 32'h0000_0002 ? add_84159 : array_index_84153[2];
  assign array_update_84161[3] = add_84043 == 32'h0000_0003 ? add_84159 : array_index_84153[3];
  assign array_update_84161[4] = add_84043 == 32'h0000_0004 ? add_84159 : array_index_84153[4];
  assign array_update_84161[5] = add_84043 == 32'h0000_0005 ? add_84159 : array_index_84153[5];
  assign array_update_84161[6] = add_84043 == 32'h0000_0006 ? add_84159 : array_index_84153[6];
  assign array_update_84161[7] = add_84043 == 32'h0000_0007 ? add_84159 : array_index_84153[7];
  assign array_update_84161[8] = add_84043 == 32'h0000_0008 ? add_84159 : array_index_84153[8];
  assign array_update_84161[9] = add_84043 == 32'h0000_0009 ? add_84159 : array_index_84153[9];
  assign add_84162 = add_84149 + 32'h0000_0001;
  assign array_update_84163[0] = add_82825 == 32'h0000_0000 ? array_update_84161 : array_update_84150[0];
  assign array_update_84163[1] = add_82825 == 32'h0000_0001 ? array_update_84161 : array_update_84150[1];
  assign array_update_84163[2] = add_82825 == 32'h0000_0002 ? array_update_84161 : array_update_84150[2];
  assign array_update_84163[3] = add_82825 == 32'h0000_0003 ? array_update_84161 : array_update_84150[3];
  assign array_update_84163[4] = add_82825 == 32'h0000_0004 ? array_update_84161 : array_update_84150[4];
  assign array_update_84163[5] = add_82825 == 32'h0000_0005 ? array_update_84161 : array_update_84150[5];
  assign array_update_84163[6] = add_82825 == 32'h0000_0006 ? array_update_84161 : array_update_84150[6];
  assign array_update_84163[7] = add_82825 == 32'h0000_0007 ? array_update_84161 : array_update_84150[7];
  assign array_update_84163[8] = add_82825 == 32'h0000_0008 ? array_update_84161 : array_update_84150[8];
  assign array_update_84163[9] = add_82825 == 32'h0000_0009 ? array_update_84161 : array_update_84150[9];
  assign array_index_84165 = array_update_72021[add_84162 > 32'h0000_0009 ? 4'h9 : add_84162[3:0]];
  assign array_index_84166 = array_update_84163[add_82825 > 32'h0000_0009 ? 4'h9 : add_82825[3:0]];
  assign smul_84170 = smul32b_32b_x_32b(array_index_82832[add_84162 > 32'h0000_0009 ? 4'h9 : add_84162[3:0]], array_index_84165[add_84043 > 32'h0000_0009 ? 4'h9 : add_84043[3:0]]);
  assign add_84172 = array_index_84166[add_84043 > 32'h0000_0009 ? 4'h9 : add_84043[3:0]] + smul_84170;
  assign array_update_84173[0] = add_84043 == 32'h0000_0000 ? add_84172 : array_index_84166[0];
  assign array_update_84173[1] = add_84043 == 32'h0000_0001 ? add_84172 : array_index_84166[1];
  assign array_update_84173[2] = add_84043 == 32'h0000_0002 ? add_84172 : array_index_84166[2];
  assign array_update_84173[3] = add_84043 == 32'h0000_0003 ? add_84172 : array_index_84166[3];
  assign array_update_84173[4] = add_84043 == 32'h0000_0004 ? add_84172 : array_index_84166[4];
  assign array_update_84173[5] = add_84043 == 32'h0000_0005 ? add_84172 : array_index_84166[5];
  assign array_update_84173[6] = add_84043 == 32'h0000_0006 ? add_84172 : array_index_84166[6];
  assign array_update_84173[7] = add_84043 == 32'h0000_0007 ? add_84172 : array_index_84166[7];
  assign array_update_84173[8] = add_84043 == 32'h0000_0008 ? add_84172 : array_index_84166[8];
  assign array_update_84173[9] = add_84043 == 32'h0000_0009 ? add_84172 : array_index_84166[9];
  assign array_update_84175[0] = add_82825 == 32'h0000_0000 ? array_update_84173 : array_update_84163[0];
  assign array_update_84175[1] = add_82825 == 32'h0000_0001 ? array_update_84173 : array_update_84163[1];
  assign array_update_84175[2] = add_82825 == 32'h0000_0002 ? array_update_84173 : array_update_84163[2];
  assign array_update_84175[3] = add_82825 == 32'h0000_0003 ? array_update_84173 : array_update_84163[3];
  assign array_update_84175[4] = add_82825 == 32'h0000_0004 ? array_update_84173 : array_update_84163[4];
  assign array_update_84175[5] = add_82825 == 32'h0000_0005 ? array_update_84173 : array_update_84163[5];
  assign array_update_84175[6] = add_82825 == 32'h0000_0006 ? array_update_84173 : array_update_84163[6];
  assign array_update_84175[7] = add_82825 == 32'h0000_0007 ? array_update_84173 : array_update_84163[7];
  assign array_update_84175[8] = add_82825 == 32'h0000_0008 ? array_update_84173 : array_update_84163[8];
  assign array_update_84175[9] = add_82825 == 32'h0000_0009 ? array_update_84173 : array_update_84163[9];
  assign add_84176 = add_82825 + 32'h0000_0001;
  assign array_index_84177 = array_update_84175[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign literal_84179 = 32'h0000_0000;
  assign array_update_84180[0] = literal_84179 == 32'h0000_0000 ? 32'h0000_0000 : array_index_84177[0];
  assign array_update_84180[1] = literal_84179 == 32'h0000_0001 ? 32'h0000_0000 : array_index_84177[1];
  assign array_update_84180[2] = literal_84179 == 32'h0000_0002 ? 32'h0000_0000 : array_index_84177[2];
  assign array_update_84180[3] = literal_84179 == 32'h0000_0003 ? 32'h0000_0000 : array_index_84177[3];
  assign array_update_84180[4] = literal_84179 == 32'h0000_0004 ? 32'h0000_0000 : array_index_84177[4];
  assign array_update_84180[5] = literal_84179 == 32'h0000_0005 ? 32'h0000_0000 : array_index_84177[5];
  assign array_update_84180[6] = literal_84179 == 32'h0000_0006 ? 32'h0000_0000 : array_index_84177[6];
  assign array_update_84180[7] = literal_84179 == 32'h0000_0007 ? 32'h0000_0000 : array_index_84177[7];
  assign array_update_84180[8] = literal_84179 == 32'h0000_0008 ? 32'h0000_0000 : array_index_84177[8];
  assign array_update_84180[9] = literal_84179 == 32'h0000_0009 ? 32'h0000_0000 : array_index_84177[9];
  assign literal_84181 = 32'h0000_0000;
  assign array_update_84182[0] = add_84176 == 32'h0000_0000 ? array_update_84180 : array_update_84175[0];
  assign array_update_84182[1] = add_84176 == 32'h0000_0001 ? array_update_84180 : array_update_84175[1];
  assign array_update_84182[2] = add_84176 == 32'h0000_0002 ? array_update_84180 : array_update_84175[2];
  assign array_update_84182[3] = add_84176 == 32'h0000_0003 ? array_update_84180 : array_update_84175[3];
  assign array_update_84182[4] = add_84176 == 32'h0000_0004 ? array_update_84180 : array_update_84175[4];
  assign array_update_84182[5] = add_84176 == 32'h0000_0005 ? array_update_84180 : array_update_84175[5];
  assign array_update_84182[6] = add_84176 == 32'h0000_0006 ? array_update_84180 : array_update_84175[6];
  assign array_update_84182[7] = add_84176 == 32'h0000_0007 ? array_update_84180 : array_update_84175[7];
  assign array_update_84182[8] = add_84176 == 32'h0000_0008 ? array_update_84180 : array_update_84175[8];
  assign array_update_84182[9] = add_84176 == 32'h0000_0009 ? array_update_84180 : array_update_84175[9];
  assign array_index_84183 = array_update_72020[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign array_index_84184 = array_update_72021[literal_84181 > 32'h0000_0009 ? 4'h9 : literal_84181[3:0]];
  assign array_index_84185 = array_update_84182[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_84189 = smul32b_32b_x_32b(array_index_84183[literal_84181 > 32'h0000_0009 ? 4'h9 : literal_84181[3:0]], array_index_84184[literal_84179 > 32'h0000_0009 ? 4'h9 : literal_84179[3:0]]);
  assign add_84191 = array_index_84185[literal_84179 > 32'h0000_0009 ? 4'h9 : literal_84179[3:0]] + smul_84189;
  assign array_update_84193[0] = literal_84179 == 32'h0000_0000 ? add_84191 : array_index_84185[0];
  assign array_update_84193[1] = literal_84179 == 32'h0000_0001 ? add_84191 : array_index_84185[1];
  assign array_update_84193[2] = literal_84179 == 32'h0000_0002 ? add_84191 : array_index_84185[2];
  assign array_update_84193[3] = literal_84179 == 32'h0000_0003 ? add_84191 : array_index_84185[3];
  assign array_update_84193[4] = literal_84179 == 32'h0000_0004 ? add_84191 : array_index_84185[4];
  assign array_update_84193[5] = literal_84179 == 32'h0000_0005 ? add_84191 : array_index_84185[5];
  assign array_update_84193[6] = literal_84179 == 32'h0000_0006 ? add_84191 : array_index_84185[6];
  assign array_update_84193[7] = literal_84179 == 32'h0000_0007 ? add_84191 : array_index_84185[7];
  assign array_update_84193[8] = literal_84179 == 32'h0000_0008 ? add_84191 : array_index_84185[8];
  assign array_update_84193[9] = literal_84179 == 32'h0000_0009 ? add_84191 : array_index_84185[9];
  assign add_84194 = literal_84181 + 32'h0000_0001;
  assign array_update_84195[0] = add_84176 == 32'h0000_0000 ? array_update_84193 : array_update_84182[0];
  assign array_update_84195[1] = add_84176 == 32'h0000_0001 ? array_update_84193 : array_update_84182[1];
  assign array_update_84195[2] = add_84176 == 32'h0000_0002 ? array_update_84193 : array_update_84182[2];
  assign array_update_84195[3] = add_84176 == 32'h0000_0003 ? array_update_84193 : array_update_84182[3];
  assign array_update_84195[4] = add_84176 == 32'h0000_0004 ? array_update_84193 : array_update_84182[4];
  assign array_update_84195[5] = add_84176 == 32'h0000_0005 ? array_update_84193 : array_update_84182[5];
  assign array_update_84195[6] = add_84176 == 32'h0000_0006 ? array_update_84193 : array_update_84182[6];
  assign array_update_84195[7] = add_84176 == 32'h0000_0007 ? array_update_84193 : array_update_84182[7];
  assign array_update_84195[8] = add_84176 == 32'h0000_0008 ? array_update_84193 : array_update_84182[8];
  assign array_update_84195[9] = add_84176 == 32'h0000_0009 ? array_update_84193 : array_update_84182[9];
  assign array_index_84197 = array_update_72021[add_84194 > 32'h0000_0009 ? 4'h9 : add_84194[3:0]];
  assign array_index_84198 = array_update_84195[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_84202 = smul32b_32b_x_32b(array_index_84183[add_84194 > 32'h0000_0009 ? 4'h9 : add_84194[3:0]], array_index_84197[literal_84179 > 32'h0000_0009 ? 4'h9 : literal_84179[3:0]]);
  assign add_84204 = array_index_84198[literal_84179 > 32'h0000_0009 ? 4'h9 : literal_84179[3:0]] + smul_84202;
  assign array_update_84206[0] = literal_84179 == 32'h0000_0000 ? add_84204 : array_index_84198[0];
  assign array_update_84206[1] = literal_84179 == 32'h0000_0001 ? add_84204 : array_index_84198[1];
  assign array_update_84206[2] = literal_84179 == 32'h0000_0002 ? add_84204 : array_index_84198[2];
  assign array_update_84206[3] = literal_84179 == 32'h0000_0003 ? add_84204 : array_index_84198[3];
  assign array_update_84206[4] = literal_84179 == 32'h0000_0004 ? add_84204 : array_index_84198[4];
  assign array_update_84206[5] = literal_84179 == 32'h0000_0005 ? add_84204 : array_index_84198[5];
  assign array_update_84206[6] = literal_84179 == 32'h0000_0006 ? add_84204 : array_index_84198[6];
  assign array_update_84206[7] = literal_84179 == 32'h0000_0007 ? add_84204 : array_index_84198[7];
  assign array_update_84206[8] = literal_84179 == 32'h0000_0008 ? add_84204 : array_index_84198[8];
  assign array_update_84206[9] = literal_84179 == 32'h0000_0009 ? add_84204 : array_index_84198[9];
  assign add_84207 = add_84194 + 32'h0000_0001;
  assign array_update_84208[0] = add_84176 == 32'h0000_0000 ? array_update_84206 : array_update_84195[0];
  assign array_update_84208[1] = add_84176 == 32'h0000_0001 ? array_update_84206 : array_update_84195[1];
  assign array_update_84208[2] = add_84176 == 32'h0000_0002 ? array_update_84206 : array_update_84195[2];
  assign array_update_84208[3] = add_84176 == 32'h0000_0003 ? array_update_84206 : array_update_84195[3];
  assign array_update_84208[4] = add_84176 == 32'h0000_0004 ? array_update_84206 : array_update_84195[4];
  assign array_update_84208[5] = add_84176 == 32'h0000_0005 ? array_update_84206 : array_update_84195[5];
  assign array_update_84208[6] = add_84176 == 32'h0000_0006 ? array_update_84206 : array_update_84195[6];
  assign array_update_84208[7] = add_84176 == 32'h0000_0007 ? array_update_84206 : array_update_84195[7];
  assign array_update_84208[8] = add_84176 == 32'h0000_0008 ? array_update_84206 : array_update_84195[8];
  assign array_update_84208[9] = add_84176 == 32'h0000_0009 ? array_update_84206 : array_update_84195[9];
  assign array_index_84210 = array_update_72021[add_84207 > 32'h0000_0009 ? 4'h9 : add_84207[3:0]];
  assign array_index_84211 = array_update_84208[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_84215 = smul32b_32b_x_32b(array_index_84183[add_84207 > 32'h0000_0009 ? 4'h9 : add_84207[3:0]], array_index_84210[literal_84179 > 32'h0000_0009 ? 4'h9 : literal_84179[3:0]]);
  assign add_84217 = array_index_84211[literal_84179 > 32'h0000_0009 ? 4'h9 : literal_84179[3:0]] + smul_84215;
  assign array_update_84219[0] = literal_84179 == 32'h0000_0000 ? add_84217 : array_index_84211[0];
  assign array_update_84219[1] = literal_84179 == 32'h0000_0001 ? add_84217 : array_index_84211[1];
  assign array_update_84219[2] = literal_84179 == 32'h0000_0002 ? add_84217 : array_index_84211[2];
  assign array_update_84219[3] = literal_84179 == 32'h0000_0003 ? add_84217 : array_index_84211[3];
  assign array_update_84219[4] = literal_84179 == 32'h0000_0004 ? add_84217 : array_index_84211[4];
  assign array_update_84219[5] = literal_84179 == 32'h0000_0005 ? add_84217 : array_index_84211[5];
  assign array_update_84219[6] = literal_84179 == 32'h0000_0006 ? add_84217 : array_index_84211[6];
  assign array_update_84219[7] = literal_84179 == 32'h0000_0007 ? add_84217 : array_index_84211[7];
  assign array_update_84219[8] = literal_84179 == 32'h0000_0008 ? add_84217 : array_index_84211[8];
  assign array_update_84219[9] = literal_84179 == 32'h0000_0009 ? add_84217 : array_index_84211[9];
  assign add_84220 = add_84207 + 32'h0000_0001;
  assign array_update_84221[0] = add_84176 == 32'h0000_0000 ? array_update_84219 : array_update_84208[0];
  assign array_update_84221[1] = add_84176 == 32'h0000_0001 ? array_update_84219 : array_update_84208[1];
  assign array_update_84221[2] = add_84176 == 32'h0000_0002 ? array_update_84219 : array_update_84208[2];
  assign array_update_84221[3] = add_84176 == 32'h0000_0003 ? array_update_84219 : array_update_84208[3];
  assign array_update_84221[4] = add_84176 == 32'h0000_0004 ? array_update_84219 : array_update_84208[4];
  assign array_update_84221[5] = add_84176 == 32'h0000_0005 ? array_update_84219 : array_update_84208[5];
  assign array_update_84221[6] = add_84176 == 32'h0000_0006 ? array_update_84219 : array_update_84208[6];
  assign array_update_84221[7] = add_84176 == 32'h0000_0007 ? array_update_84219 : array_update_84208[7];
  assign array_update_84221[8] = add_84176 == 32'h0000_0008 ? array_update_84219 : array_update_84208[8];
  assign array_update_84221[9] = add_84176 == 32'h0000_0009 ? array_update_84219 : array_update_84208[9];
  assign array_index_84223 = array_update_72021[add_84220 > 32'h0000_0009 ? 4'h9 : add_84220[3:0]];
  assign array_index_84224 = array_update_84221[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_84228 = smul32b_32b_x_32b(array_index_84183[add_84220 > 32'h0000_0009 ? 4'h9 : add_84220[3:0]], array_index_84223[literal_84179 > 32'h0000_0009 ? 4'h9 : literal_84179[3:0]]);
  assign add_84230 = array_index_84224[literal_84179 > 32'h0000_0009 ? 4'h9 : literal_84179[3:0]] + smul_84228;
  assign array_update_84232[0] = literal_84179 == 32'h0000_0000 ? add_84230 : array_index_84224[0];
  assign array_update_84232[1] = literal_84179 == 32'h0000_0001 ? add_84230 : array_index_84224[1];
  assign array_update_84232[2] = literal_84179 == 32'h0000_0002 ? add_84230 : array_index_84224[2];
  assign array_update_84232[3] = literal_84179 == 32'h0000_0003 ? add_84230 : array_index_84224[3];
  assign array_update_84232[4] = literal_84179 == 32'h0000_0004 ? add_84230 : array_index_84224[4];
  assign array_update_84232[5] = literal_84179 == 32'h0000_0005 ? add_84230 : array_index_84224[5];
  assign array_update_84232[6] = literal_84179 == 32'h0000_0006 ? add_84230 : array_index_84224[6];
  assign array_update_84232[7] = literal_84179 == 32'h0000_0007 ? add_84230 : array_index_84224[7];
  assign array_update_84232[8] = literal_84179 == 32'h0000_0008 ? add_84230 : array_index_84224[8];
  assign array_update_84232[9] = literal_84179 == 32'h0000_0009 ? add_84230 : array_index_84224[9];
  assign add_84233 = add_84220 + 32'h0000_0001;
  assign array_update_84234[0] = add_84176 == 32'h0000_0000 ? array_update_84232 : array_update_84221[0];
  assign array_update_84234[1] = add_84176 == 32'h0000_0001 ? array_update_84232 : array_update_84221[1];
  assign array_update_84234[2] = add_84176 == 32'h0000_0002 ? array_update_84232 : array_update_84221[2];
  assign array_update_84234[3] = add_84176 == 32'h0000_0003 ? array_update_84232 : array_update_84221[3];
  assign array_update_84234[4] = add_84176 == 32'h0000_0004 ? array_update_84232 : array_update_84221[4];
  assign array_update_84234[5] = add_84176 == 32'h0000_0005 ? array_update_84232 : array_update_84221[5];
  assign array_update_84234[6] = add_84176 == 32'h0000_0006 ? array_update_84232 : array_update_84221[6];
  assign array_update_84234[7] = add_84176 == 32'h0000_0007 ? array_update_84232 : array_update_84221[7];
  assign array_update_84234[8] = add_84176 == 32'h0000_0008 ? array_update_84232 : array_update_84221[8];
  assign array_update_84234[9] = add_84176 == 32'h0000_0009 ? array_update_84232 : array_update_84221[9];
  assign array_index_84236 = array_update_72021[add_84233 > 32'h0000_0009 ? 4'h9 : add_84233[3:0]];
  assign array_index_84237 = array_update_84234[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_84241 = smul32b_32b_x_32b(array_index_84183[add_84233 > 32'h0000_0009 ? 4'h9 : add_84233[3:0]], array_index_84236[literal_84179 > 32'h0000_0009 ? 4'h9 : literal_84179[3:0]]);
  assign add_84243 = array_index_84237[literal_84179 > 32'h0000_0009 ? 4'h9 : literal_84179[3:0]] + smul_84241;
  assign array_update_84245[0] = literal_84179 == 32'h0000_0000 ? add_84243 : array_index_84237[0];
  assign array_update_84245[1] = literal_84179 == 32'h0000_0001 ? add_84243 : array_index_84237[1];
  assign array_update_84245[2] = literal_84179 == 32'h0000_0002 ? add_84243 : array_index_84237[2];
  assign array_update_84245[3] = literal_84179 == 32'h0000_0003 ? add_84243 : array_index_84237[3];
  assign array_update_84245[4] = literal_84179 == 32'h0000_0004 ? add_84243 : array_index_84237[4];
  assign array_update_84245[5] = literal_84179 == 32'h0000_0005 ? add_84243 : array_index_84237[5];
  assign array_update_84245[6] = literal_84179 == 32'h0000_0006 ? add_84243 : array_index_84237[6];
  assign array_update_84245[7] = literal_84179 == 32'h0000_0007 ? add_84243 : array_index_84237[7];
  assign array_update_84245[8] = literal_84179 == 32'h0000_0008 ? add_84243 : array_index_84237[8];
  assign array_update_84245[9] = literal_84179 == 32'h0000_0009 ? add_84243 : array_index_84237[9];
  assign add_84246 = add_84233 + 32'h0000_0001;
  assign array_update_84247[0] = add_84176 == 32'h0000_0000 ? array_update_84245 : array_update_84234[0];
  assign array_update_84247[1] = add_84176 == 32'h0000_0001 ? array_update_84245 : array_update_84234[1];
  assign array_update_84247[2] = add_84176 == 32'h0000_0002 ? array_update_84245 : array_update_84234[2];
  assign array_update_84247[3] = add_84176 == 32'h0000_0003 ? array_update_84245 : array_update_84234[3];
  assign array_update_84247[4] = add_84176 == 32'h0000_0004 ? array_update_84245 : array_update_84234[4];
  assign array_update_84247[5] = add_84176 == 32'h0000_0005 ? array_update_84245 : array_update_84234[5];
  assign array_update_84247[6] = add_84176 == 32'h0000_0006 ? array_update_84245 : array_update_84234[6];
  assign array_update_84247[7] = add_84176 == 32'h0000_0007 ? array_update_84245 : array_update_84234[7];
  assign array_update_84247[8] = add_84176 == 32'h0000_0008 ? array_update_84245 : array_update_84234[8];
  assign array_update_84247[9] = add_84176 == 32'h0000_0009 ? array_update_84245 : array_update_84234[9];
  assign array_index_84249 = array_update_72021[add_84246 > 32'h0000_0009 ? 4'h9 : add_84246[3:0]];
  assign array_index_84250 = array_update_84247[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_84254 = smul32b_32b_x_32b(array_index_84183[add_84246 > 32'h0000_0009 ? 4'h9 : add_84246[3:0]], array_index_84249[literal_84179 > 32'h0000_0009 ? 4'h9 : literal_84179[3:0]]);
  assign add_84256 = array_index_84250[literal_84179 > 32'h0000_0009 ? 4'h9 : literal_84179[3:0]] + smul_84254;
  assign array_update_84258[0] = literal_84179 == 32'h0000_0000 ? add_84256 : array_index_84250[0];
  assign array_update_84258[1] = literal_84179 == 32'h0000_0001 ? add_84256 : array_index_84250[1];
  assign array_update_84258[2] = literal_84179 == 32'h0000_0002 ? add_84256 : array_index_84250[2];
  assign array_update_84258[3] = literal_84179 == 32'h0000_0003 ? add_84256 : array_index_84250[3];
  assign array_update_84258[4] = literal_84179 == 32'h0000_0004 ? add_84256 : array_index_84250[4];
  assign array_update_84258[5] = literal_84179 == 32'h0000_0005 ? add_84256 : array_index_84250[5];
  assign array_update_84258[6] = literal_84179 == 32'h0000_0006 ? add_84256 : array_index_84250[6];
  assign array_update_84258[7] = literal_84179 == 32'h0000_0007 ? add_84256 : array_index_84250[7];
  assign array_update_84258[8] = literal_84179 == 32'h0000_0008 ? add_84256 : array_index_84250[8];
  assign array_update_84258[9] = literal_84179 == 32'h0000_0009 ? add_84256 : array_index_84250[9];
  assign add_84259 = add_84246 + 32'h0000_0001;
  assign array_update_84260[0] = add_84176 == 32'h0000_0000 ? array_update_84258 : array_update_84247[0];
  assign array_update_84260[1] = add_84176 == 32'h0000_0001 ? array_update_84258 : array_update_84247[1];
  assign array_update_84260[2] = add_84176 == 32'h0000_0002 ? array_update_84258 : array_update_84247[2];
  assign array_update_84260[3] = add_84176 == 32'h0000_0003 ? array_update_84258 : array_update_84247[3];
  assign array_update_84260[4] = add_84176 == 32'h0000_0004 ? array_update_84258 : array_update_84247[4];
  assign array_update_84260[5] = add_84176 == 32'h0000_0005 ? array_update_84258 : array_update_84247[5];
  assign array_update_84260[6] = add_84176 == 32'h0000_0006 ? array_update_84258 : array_update_84247[6];
  assign array_update_84260[7] = add_84176 == 32'h0000_0007 ? array_update_84258 : array_update_84247[7];
  assign array_update_84260[8] = add_84176 == 32'h0000_0008 ? array_update_84258 : array_update_84247[8];
  assign array_update_84260[9] = add_84176 == 32'h0000_0009 ? array_update_84258 : array_update_84247[9];
  assign array_index_84262 = array_update_72021[add_84259 > 32'h0000_0009 ? 4'h9 : add_84259[3:0]];
  assign array_index_84263 = array_update_84260[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_84267 = smul32b_32b_x_32b(array_index_84183[add_84259 > 32'h0000_0009 ? 4'h9 : add_84259[3:0]], array_index_84262[literal_84179 > 32'h0000_0009 ? 4'h9 : literal_84179[3:0]]);
  assign add_84269 = array_index_84263[literal_84179 > 32'h0000_0009 ? 4'h9 : literal_84179[3:0]] + smul_84267;
  assign array_update_84271[0] = literal_84179 == 32'h0000_0000 ? add_84269 : array_index_84263[0];
  assign array_update_84271[1] = literal_84179 == 32'h0000_0001 ? add_84269 : array_index_84263[1];
  assign array_update_84271[2] = literal_84179 == 32'h0000_0002 ? add_84269 : array_index_84263[2];
  assign array_update_84271[3] = literal_84179 == 32'h0000_0003 ? add_84269 : array_index_84263[3];
  assign array_update_84271[4] = literal_84179 == 32'h0000_0004 ? add_84269 : array_index_84263[4];
  assign array_update_84271[5] = literal_84179 == 32'h0000_0005 ? add_84269 : array_index_84263[5];
  assign array_update_84271[6] = literal_84179 == 32'h0000_0006 ? add_84269 : array_index_84263[6];
  assign array_update_84271[7] = literal_84179 == 32'h0000_0007 ? add_84269 : array_index_84263[7];
  assign array_update_84271[8] = literal_84179 == 32'h0000_0008 ? add_84269 : array_index_84263[8];
  assign array_update_84271[9] = literal_84179 == 32'h0000_0009 ? add_84269 : array_index_84263[9];
  assign add_84272 = add_84259 + 32'h0000_0001;
  assign array_update_84273[0] = add_84176 == 32'h0000_0000 ? array_update_84271 : array_update_84260[0];
  assign array_update_84273[1] = add_84176 == 32'h0000_0001 ? array_update_84271 : array_update_84260[1];
  assign array_update_84273[2] = add_84176 == 32'h0000_0002 ? array_update_84271 : array_update_84260[2];
  assign array_update_84273[3] = add_84176 == 32'h0000_0003 ? array_update_84271 : array_update_84260[3];
  assign array_update_84273[4] = add_84176 == 32'h0000_0004 ? array_update_84271 : array_update_84260[4];
  assign array_update_84273[5] = add_84176 == 32'h0000_0005 ? array_update_84271 : array_update_84260[5];
  assign array_update_84273[6] = add_84176 == 32'h0000_0006 ? array_update_84271 : array_update_84260[6];
  assign array_update_84273[7] = add_84176 == 32'h0000_0007 ? array_update_84271 : array_update_84260[7];
  assign array_update_84273[8] = add_84176 == 32'h0000_0008 ? array_update_84271 : array_update_84260[8];
  assign array_update_84273[9] = add_84176 == 32'h0000_0009 ? array_update_84271 : array_update_84260[9];
  assign array_index_84275 = array_update_72021[add_84272 > 32'h0000_0009 ? 4'h9 : add_84272[3:0]];
  assign array_index_84276 = array_update_84273[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_84280 = smul32b_32b_x_32b(array_index_84183[add_84272 > 32'h0000_0009 ? 4'h9 : add_84272[3:0]], array_index_84275[literal_84179 > 32'h0000_0009 ? 4'h9 : literal_84179[3:0]]);
  assign add_84282 = array_index_84276[literal_84179 > 32'h0000_0009 ? 4'h9 : literal_84179[3:0]] + smul_84280;
  assign array_update_84284[0] = literal_84179 == 32'h0000_0000 ? add_84282 : array_index_84276[0];
  assign array_update_84284[1] = literal_84179 == 32'h0000_0001 ? add_84282 : array_index_84276[1];
  assign array_update_84284[2] = literal_84179 == 32'h0000_0002 ? add_84282 : array_index_84276[2];
  assign array_update_84284[3] = literal_84179 == 32'h0000_0003 ? add_84282 : array_index_84276[3];
  assign array_update_84284[4] = literal_84179 == 32'h0000_0004 ? add_84282 : array_index_84276[4];
  assign array_update_84284[5] = literal_84179 == 32'h0000_0005 ? add_84282 : array_index_84276[5];
  assign array_update_84284[6] = literal_84179 == 32'h0000_0006 ? add_84282 : array_index_84276[6];
  assign array_update_84284[7] = literal_84179 == 32'h0000_0007 ? add_84282 : array_index_84276[7];
  assign array_update_84284[8] = literal_84179 == 32'h0000_0008 ? add_84282 : array_index_84276[8];
  assign array_update_84284[9] = literal_84179 == 32'h0000_0009 ? add_84282 : array_index_84276[9];
  assign add_84285 = add_84272 + 32'h0000_0001;
  assign array_update_84286[0] = add_84176 == 32'h0000_0000 ? array_update_84284 : array_update_84273[0];
  assign array_update_84286[1] = add_84176 == 32'h0000_0001 ? array_update_84284 : array_update_84273[1];
  assign array_update_84286[2] = add_84176 == 32'h0000_0002 ? array_update_84284 : array_update_84273[2];
  assign array_update_84286[3] = add_84176 == 32'h0000_0003 ? array_update_84284 : array_update_84273[3];
  assign array_update_84286[4] = add_84176 == 32'h0000_0004 ? array_update_84284 : array_update_84273[4];
  assign array_update_84286[5] = add_84176 == 32'h0000_0005 ? array_update_84284 : array_update_84273[5];
  assign array_update_84286[6] = add_84176 == 32'h0000_0006 ? array_update_84284 : array_update_84273[6];
  assign array_update_84286[7] = add_84176 == 32'h0000_0007 ? array_update_84284 : array_update_84273[7];
  assign array_update_84286[8] = add_84176 == 32'h0000_0008 ? array_update_84284 : array_update_84273[8];
  assign array_update_84286[9] = add_84176 == 32'h0000_0009 ? array_update_84284 : array_update_84273[9];
  assign array_index_84288 = array_update_72021[add_84285 > 32'h0000_0009 ? 4'h9 : add_84285[3:0]];
  assign array_index_84289 = array_update_84286[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_84293 = smul32b_32b_x_32b(array_index_84183[add_84285 > 32'h0000_0009 ? 4'h9 : add_84285[3:0]], array_index_84288[literal_84179 > 32'h0000_0009 ? 4'h9 : literal_84179[3:0]]);
  assign add_84295 = array_index_84289[literal_84179 > 32'h0000_0009 ? 4'h9 : literal_84179[3:0]] + smul_84293;
  assign array_update_84297[0] = literal_84179 == 32'h0000_0000 ? add_84295 : array_index_84289[0];
  assign array_update_84297[1] = literal_84179 == 32'h0000_0001 ? add_84295 : array_index_84289[1];
  assign array_update_84297[2] = literal_84179 == 32'h0000_0002 ? add_84295 : array_index_84289[2];
  assign array_update_84297[3] = literal_84179 == 32'h0000_0003 ? add_84295 : array_index_84289[3];
  assign array_update_84297[4] = literal_84179 == 32'h0000_0004 ? add_84295 : array_index_84289[4];
  assign array_update_84297[5] = literal_84179 == 32'h0000_0005 ? add_84295 : array_index_84289[5];
  assign array_update_84297[6] = literal_84179 == 32'h0000_0006 ? add_84295 : array_index_84289[6];
  assign array_update_84297[7] = literal_84179 == 32'h0000_0007 ? add_84295 : array_index_84289[7];
  assign array_update_84297[8] = literal_84179 == 32'h0000_0008 ? add_84295 : array_index_84289[8];
  assign array_update_84297[9] = literal_84179 == 32'h0000_0009 ? add_84295 : array_index_84289[9];
  assign add_84298 = add_84285 + 32'h0000_0001;
  assign array_update_84299[0] = add_84176 == 32'h0000_0000 ? array_update_84297 : array_update_84286[0];
  assign array_update_84299[1] = add_84176 == 32'h0000_0001 ? array_update_84297 : array_update_84286[1];
  assign array_update_84299[2] = add_84176 == 32'h0000_0002 ? array_update_84297 : array_update_84286[2];
  assign array_update_84299[3] = add_84176 == 32'h0000_0003 ? array_update_84297 : array_update_84286[3];
  assign array_update_84299[4] = add_84176 == 32'h0000_0004 ? array_update_84297 : array_update_84286[4];
  assign array_update_84299[5] = add_84176 == 32'h0000_0005 ? array_update_84297 : array_update_84286[5];
  assign array_update_84299[6] = add_84176 == 32'h0000_0006 ? array_update_84297 : array_update_84286[6];
  assign array_update_84299[7] = add_84176 == 32'h0000_0007 ? array_update_84297 : array_update_84286[7];
  assign array_update_84299[8] = add_84176 == 32'h0000_0008 ? array_update_84297 : array_update_84286[8];
  assign array_update_84299[9] = add_84176 == 32'h0000_0009 ? array_update_84297 : array_update_84286[9];
  assign array_index_84301 = array_update_72021[add_84298 > 32'h0000_0009 ? 4'h9 : add_84298[3:0]];
  assign array_index_84302 = array_update_84299[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_84306 = smul32b_32b_x_32b(array_index_84183[add_84298 > 32'h0000_0009 ? 4'h9 : add_84298[3:0]], array_index_84301[literal_84179 > 32'h0000_0009 ? 4'h9 : literal_84179[3:0]]);
  assign add_84308 = array_index_84302[literal_84179 > 32'h0000_0009 ? 4'h9 : literal_84179[3:0]] + smul_84306;
  assign array_update_84309[0] = literal_84179 == 32'h0000_0000 ? add_84308 : array_index_84302[0];
  assign array_update_84309[1] = literal_84179 == 32'h0000_0001 ? add_84308 : array_index_84302[1];
  assign array_update_84309[2] = literal_84179 == 32'h0000_0002 ? add_84308 : array_index_84302[2];
  assign array_update_84309[3] = literal_84179 == 32'h0000_0003 ? add_84308 : array_index_84302[3];
  assign array_update_84309[4] = literal_84179 == 32'h0000_0004 ? add_84308 : array_index_84302[4];
  assign array_update_84309[5] = literal_84179 == 32'h0000_0005 ? add_84308 : array_index_84302[5];
  assign array_update_84309[6] = literal_84179 == 32'h0000_0006 ? add_84308 : array_index_84302[6];
  assign array_update_84309[7] = literal_84179 == 32'h0000_0007 ? add_84308 : array_index_84302[7];
  assign array_update_84309[8] = literal_84179 == 32'h0000_0008 ? add_84308 : array_index_84302[8];
  assign array_update_84309[9] = literal_84179 == 32'h0000_0009 ? add_84308 : array_index_84302[9];
  assign array_update_84310[0] = add_84176 == 32'h0000_0000 ? array_update_84309 : array_update_84299[0];
  assign array_update_84310[1] = add_84176 == 32'h0000_0001 ? array_update_84309 : array_update_84299[1];
  assign array_update_84310[2] = add_84176 == 32'h0000_0002 ? array_update_84309 : array_update_84299[2];
  assign array_update_84310[3] = add_84176 == 32'h0000_0003 ? array_update_84309 : array_update_84299[3];
  assign array_update_84310[4] = add_84176 == 32'h0000_0004 ? array_update_84309 : array_update_84299[4];
  assign array_update_84310[5] = add_84176 == 32'h0000_0005 ? array_update_84309 : array_update_84299[5];
  assign array_update_84310[6] = add_84176 == 32'h0000_0006 ? array_update_84309 : array_update_84299[6];
  assign array_update_84310[7] = add_84176 == 32'h0000_0007 ? array_update_84309 : array_update_84299[7];
  assign array_update_84310[8] = add_84176 == 32'h0000_0008 ? array_update_84309 : array_update_84299[8];
  assign array_update_84310[9] = add_84176 == 32'h0000_0009 ? array_update_84309 : array_update_84299[9];
  assign array_index_84312 = array_update_84310[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign add_84314 = literal_84179 + 32'h0000_0001;
  assign array_update_84315[0] = add_84314 == 32'h0000_0000 ? 32'h0000_0000 : array_index_84312[0];
  assign array_update_84315[1] = add_84314 == 32'h0000_0001 ? 32'h0000_0000 : array_index_84312[1];
  assign array_update_84315[2] = add_84314 == 32'h0000_0002 ? 32'h0000_0000 : array_index_84312[2];
  assign array_update_84315[3] = add_84314 == 32'h0000_0003 ? 32'h0000_0000 : array_index_84312[3];
  assign array_update_84315[4] = add_84314 == 32'h0000_0004 ? 32'h0000_0000 : array_index_84312[4];
  assign array_update_84315[5] = add_84314 == 32'h0000_0005 ? 32'h0000_0000 : array_index_84312[5];
  assign array_update_84315[6] = add_84314 == 32'h0000_0006 ? 32'h0000_0000 : array_index_84312[6];
  assign array_update_84315[7] = add_84314 == 32'h0000_0007 ? 32'h0000_0000 : array_index_84312[7];
  assign array_update_84315[8] = add_84314 == 32'h0000_0008 ? 32'h0000_0000 : array_index_84312[8];
  assign array_update_84315[9] = add_84314 == 32'h0000_0009 ? 32'h0000_0000 : array_index_84312[9];
  assign literal_84316 = 32'h0000_0000;
  assign array_update_84317[0] = add_84176 == 32'h0000_0000 ? array_update_84315 : array_update_84310[0];
  assign array_update_84317[1] = add_84176 == 32'h0000_0001 ? array_update_84315 : array_update_84310[1];
  assign array_update_84317[2] = add_84176 == 32'h0000_0002 ? array_update_84315 : array_update_84310[2];
  assign array_update_84317[3] = add_84176 == 32'h0000_0003 ? array_update_84315 : array_update_84310[3];
  assign array_update_84317[4] = add_84176 == 32'h0000_0004 ? array_update_84315 : array_update_84310[4];
  assign array_update_84317[5] = add_84176 == 32'h0000_0005 ? array_update_84315 : array_update_84310[5];
  assign array_update_84317[6] = add_84176 == 32'h0000_0006 ? array_update_84315 : array_update_84310[6];
  assign array_update_84317[7] = add_84176 == 32'h0000_0007 ? array_update_84315 : array_update_84310[7];
  assign array_update_84317[8] = add_84176 == 32'h0000_0008 ? array_update_84315 : array_update_84310[8];
  assign array_update_84317[9] = add_84176 == 32'h0000_0009 ? array_update_84315 : array_update_84310[9];
  assign array_index_84319 = array_update_72021[literal_84316 > 32'h0000_0009 ? 4'h9 : literal_84316[3:0]];
  assign array_index_84320 = array_update_84317[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_84324 = smul32b_32b_x_32b(array_index_84183[literal_84316 > 32'h0000_0009 ? 4'h9 : literal_84316[3:0]], array_index_84319[add_84314 > 32'h0000_0009 ? 4'h9 : add_84314[3:0]]);
  assign add_84326 = array_index_84320[add_84314 > 32'h0000_0009 ? 4'h9 : add_84314[3:0]] + smul_84324;
  assign array_update_84328[0] = add_84314 == 32'h0000_0000 ? add_84326 : array_index_84320[0];
  assign array_update_84328[1] = add_84314 == 32'h0000_0001 ? add_84326 : array_index_84320[1];
  assign array_update_84328[2] = add_84314 == 32'h0000_0002 ? add_84326 : array_index_84320[2];
  assign array_update_84328[3] = add_84314 == 32'h0000_0003 ? add_84326 : array_index_84320[3];
  assign array_update_84328[4] = add_84314 == 32'h0000_0004 ? add_84326 : array_index_84320[4];
  assign array_update_84328[5] = add_84314 == 32'h0000_0005 ? add_84326 : array_index_84320[5];
  assign array_update_84328[6] = add_84314 == 32'h0000_0006 ? add_84326 : array_index_84320[6];
  assign array_update_84328[7] = add_84314 == 32'h0000_0007 ? add_84326 : array_index_84320[7];
  assign array_update_84328[8] = add_84314 == 32'h0000_0008 ? add_84326 : array_index_84320[8];
  assign array_update_84328[9] = add_84314 == 32'h0000_0009 ? add_84326 : array_index_84320[9];
  assign add_84329 = literal_84316 + 32'h0000_0001;
  assign array_update_84330[0] = add_84176 == 32'h0000_0000 ? array_update_84328 : array_update_84317[0];
  assign array_update_84330[1] = add_84176 == 32'h0000_0001 ? array_update_84328 : array_update_84317[1];
  assign array_update_84330[2] = add_84176 == 32'h0000_0002 ? array_update_84328 : array_update_84317[2];
  assign array_update_84330[3] = add_84176 == 32'h0000_0003 ? array_update_84328 : array_update_84317[3];
  assign array_update_84330[4] = add_84176 == 32'h0000_0004 ? array_update_84328 : array_update_84317[4];
  assign array_update_84330[5] = add_84176 == 32'h0000_0005 ? array_update_84328 : array_update_84317[5];
  assign array_update_84330[6] = add_84176 == 32'h0000_0006 ? array_update_84328 : array_update_84317[6];
  assign array_update_84330[7] = add_84176 == 32'h0000_0007 ? array_update_84328 : array_update_84317[7];
  assign array_update_84330[8] = add_84176 == 32'h0000_0008 ? array_update_84328 : array_update_84317[8];
  assign array_update_84330[9] = add_84176 == 32'h0000_0009 ? array_update_84328 : array_update_84317[9];
  assign array_index_84332 = array_update_72021[add_84329 > 32'h0000_0009 ? 4'h9 : add_84329[3:0]];
  assign array_index_84333 = array_update_84330[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_84337 = smul32b_32b_x_32b(array_index_84183[add_84329 > 32'h0000_0009 ? 4'h9 : add_84329[3:0]], array_index_84332[add_84314 > 32'h0000_0009 ? 4'h9 : add_84314[3:0]]);
  assign add_84339 = array_index_84333[add_84314 > 32'h0000_0009 ? 4'h9 : add_84314[3:0]] + smul_84337;
  assign array_update_84341[0] = add_84314 == 32'h0000_0000 ? add_84339 : array_index_84333[0];
  assign array_update_84341[1] = add_84314 == 32'h0000_0001 ? add_84339 : array_index_84333[1];
  assign array_update_84341[2] = add_84314 == 32'h0000_0002 ? add_84339 : array_index_84333[2];
  assign array_update_84341[3] = add_84314 == 32'h0000_0003 ? add_84339 : array_index_84333[3];
  assign array_update_84341[4] = add_84314 == 32'h0000_0004 ? add_84339 : array_index_84333[4];
  assign array_update_84341[5] = add_84314 == 32'h0000_0005 ? add_84339 : array_index_84333[5];
  assign array_update_84341[6] = add_84314 == 32'h0000_0006 ? add_84339 : array_index_84333[6];
  assign array_update_84341[7] = add_84314 == 32'h0000_0007 ? add_84339 : array_index_84333[7];
  assign array_update_84341[8] = add_84314 == 32'h0000_0008 ? add_84339 : array_index_84333[8];
  assign array_update_84341[9] = add_84314 == 32'h0000_0009 ? add_84339 : array_index_84333[9];
  assign add_84342 = add_84329 + 32'h0000_0001;
  assign array_update_84343[0] = add_84176 == 32'h0000_0000 ? array_update_84341 : array_update_84330[0];
  assign array_update_84343[1] = add_84176 == 32'h0000_0001 ? array_update_84341 : array_update_84330[1];
  assign array_update_84343[2] = add_84176 == 32'h0000_0002 ? array_update_84341 : array_update_84330[2];
  assign array_update_84343[3] = add_84176 == 32'h0000_0003 ? array_update_84341 : array_update_84330[3];
  assign array_update_84343[4] = add_84176 == 32'h0000_0004 ? array_update_84341 : array_update_84330[4];
  assign array_update_84343[5] = add_84176 == 32'h0000_0005 ? array_update_84341 : array_update_84330[5];
  assign array_update_84343[6] = add_84176 == 32'h0000_0006 ? array_update_84341 : array_update_84330[6];
  assign array_update_84343[7] = add_84176 == 32'h0000_0007 ? array_update_84341 : array_update_84330[7];
  assign array_update_84343[8] = add_84176 == 32'h0000_0008 ? array_update_84341 : array_update_84330[8];
  assign array_update_84343[9] = add_84176 == 32'h0000_0009 ? array_update_84341 : array_update_84330[9];
  assign array_index_84345 = array_update_72021[add_84342 > 32'h0000_0009 ? 4'h9 : add_84342[3:0]];
  assign array_index_84346 = array_update_84343[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_84350 = smul32b_32b_x_32b(array_index_84183[add_84342 > 32'h0000_0009 ? 4'h9 : add_84342[3:0]], array_index_84345[add_84314 > 32'h0000_0009 ? 4'h9 : add_84314[3:0]]);
  assign add_84352 = array_index_84346[add_84314 > 32'h0000_0009 ? 4'h9 : add_84314[3:0]] + smul_84350;
  assign array_update_84354[0] = add_84314 == 32'h0000_0000 ? add_84352 : array_index_84346[0];
  assign array_update_84354[1] = add_84314 == 32'h0000_0001 ? add_84352 : array_index_84346[1];
  assign array_update_84354[2] = add_84314 == 32'h0000_0002 ? add_84352 : array_index_84346[2];
  assign array_update_84354[3] = add_84314 == 32'h0000_0003 ? add_84352 : array_index_84346[3];
  assign array_update_84354[4] = add_84314 == 32'h0000_0004 ? add_84352 : array_index_84346[4];
  assign array_update_84354[5] = add_84314 == 32'h0000_0005 ? add_84352 : array_index_84346[5];
  assign array_update_84354[6] = add_84314 == 32'h0000_0006 ? add_84352 : array_index_84346[6];
  assign array_update_84354[7] = add_84314 == 32'h0000_0007 ? add_84352 : array_index_84346[7];
  assign array_update_84354[8] = add_84314 == 32'h0000_0008 ? add_84352 : array_index_84346[8];
  assign array_update_84354[9] = add_84314 == 32'h0000_0009 ? add_84352 : array_index_84346[9];
  assign add_84355 = add_84342 + 32'h0000_0001;
  assign array_update_84356[0] = add_84176 == 32'h0000_0000 ? array_update_84354 : array_update_84343[0];
  assign array_update_84356[1] = add_84176 == 32'h0000_0001 ? array_update_84354 : array_update_84343[1];
  assign array_update_84356[2] = add_84176 == 32'h0000_0002 ? array_update_84354 : array_update_84343[2];
  assign array_update_84356[3] = add_84176 == 32'h0000_0003 ? array_update_84354 : array_update_84343[3];
  assign array_update_84356[4] = add_84176 == 32'h0000_0004 ? array_update_84354 : array_update_84343[4];
  assign array_update_84356[5] = add_84176 == 32'h0000_0005 ? array_update_84354 : array_update_84343[5];
  assign array_update_84356[6] = add_84176 == 32'h0000_0006 ? array_update_84354 : array_update_84343[6];
  assign array_update_84356[7] = add_84176 == 32'h0000_0007 ? array_update_84354 : array_update_84343[7];
  assign array_update_84356[8] = add_84176 == 32'h0000_0008 ? array_update_84354 : array_update_84343[8];
  assign array_update_84356[9] = add_84176 == 32'h0000_0009 ? array_update_84354 : array_update_84343[9];
  assign array_index_84358 = array_update_72021[add_84355 > 32'h0000_0009 ? 4'h9 : add_84355[3:0]];
  assign array_index_84359 = array_update_84356[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_84363 = smul32b_32b_x_32b(array_index_84183[add_84355 > 32'h0000_0009 ? 4'h9 : add_84355[3:0]], array_index_84358[add_84314 > 32'h0000_0009 ? 4'h9 : add_84314[3:0]]);
  assign add_84365 = array_index_84359[add_84314 > 32'h0000_0009 ? 4'h9 : add_84314[3:0]] + smul_84363;
  assign array_update_84367[0] = add_84314 == 32'h0000_0000 ? add_84365 : array_index_84359[0];
  assign array_update_84367[1] = add_84314 == 32'h0000_0001 ? add_84365 : array_index_84359[1];
  assign array_update_84367[2] = add_84314 == 32'h0000_0002 ? add_84365 : array_index_84359[2];
  assign array_update_84367[3] = add_84314 == 32'h0000_0003 ? add_84365 : array_index_84359[3];
  assign array_update_84367[4] = add_84314 == 32'h0000_0004 ? add_84365 : array_index_84359[4];
  assign array_update_84367[5] = add_84314 == 32'h0000_0005 ? add_84365 : array_index_84359[5];
  assign array_update_84367[6] = add_84314 == 32'h0000_0006 ? add_84365 : array_index_84359[6];
  assign array_update_84367[7] = add_84314 == 32'h0000_0007 ? add_84365 : array_index_84359[7];
  assign array_update_84367[8] = add_84314 == 32'h0000_0008 ? add_84365 : array_index_84359[8];
  assign array_update_84367[9] = add_84314 == 32'h0000_0009 ? add_84365 : array_index_84359[9];
  assign add_84368 = add_84355 + 32'h0000_0001;
  assign array_update_84369[0] = add_84176 == 32'h0000_0000 ? array_update_84367 : array_update_84356[0];
  assign array_update_84369[1] = add_84176 == 32'h0000_0001 ? array_update_84367 : array_update_84356[1];
  assign array_update_84369[2] = add_84176 == 32'h0000_0002 ? array_update_84367 : array_update_84356[2];
  assign array_update_84369[3] = add_84176 == 32'h0000_0003 ? array_update_84367 : array_update_84356[3];
  assign array_update_84369[4] = add_84176 == 32'h0000_0004 ? array_update_84367 : array_update_84356[4];
  assign array_update_84369[5] = add_84176 == 32'h0000_0005 ? array_update_84367 : array_update_84356[5];
  assign array_update_84369[6] = add_84176 == 32'h0000_0006 ? array_update_84367 : array_update_84356[6];
  assign array_update_84369[7] = add_84176 == 32'h0000_0007 ? array_update_84367 : array_update_84356[7];
  assign array_update_84369[8] = add_84176 == 32'h0000_0008 ? array_update_84367 : array_update_84356[8];
  assign array_update_84369[9] = add_84176 == 32'h0000_0009 ? array_update_84367 : array_update_84356[9];
  assign array_index_84371 = array_update_72021[add_84368 > 32'h0000_0009 ? 4'h9 : add_84368[3:0]];
  assign array_index_84372 = array_update_84369[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_84376 = smul32b_32b_x_32b(array_index_84183[add_84368 > 32'h0000_0009 ? 4'h9 : add_84368[3:0]], array_index_84371[add_84314 > 32'h0000_0009 ? 4'h9 : add_84314[3:0]]);
  assign add_84378 = array_index_84372[add_84314 > 32'h0000_0009 ? 4'h9 : add_84314[3:0]] + smul_84376;
  assign array_update_84380[0] = add_84314 == 32'h0000_0000 ? add_84378 : array_index_84372[0];
  assign array_update_84380[1] = add_84314 == 32'h0000_0001 ? add_84378 : array_index_84372[1];
  assign array_update_84380[2] = add_84314 == 32'h0000_0002 ? add_84378 : array_index_84372[2];
  assign array_update_84380[3] = add_84314 == 32'h0000_0003 ? add_84378 : array_index_84372[3];
  assign array_update_84380[4] = add_84314 == 32'h0000_0004 ? add_84378 : array_index_84372[4];
  assign array_update_84380[5] = add_84314 == 32'h0000_0005 ? add_84378 : array_index_84372[5];
  assign array_update_84380[6] = add_84314 == 32'h0000_0006 ? add_84378 : array_index_84372[6];
  assign array_update_84380[7] = add_84314 == 32'h0000_0007 ? add_84378 : array_index_84372[7];
  assign array_update_84380[8] = add_84314 == 32'h0000_0008 ? add_84378 : array_index_84372[8];
  assign array_update_84380[9] = add_84314 == 32'h0000_0009 ? add_84378 : array_index_84372[9];
  assign add_84381 = add_84368 + 32'h0000_0001;
  assign array_update_84382[0] = add_84176 == 32'h0000_0000 ? array_update_84380 : array_update_84369[0];
  assign array_update_84382[1] = add_84176 == 32'h0000_0001 ? array_update_84380 : array_update_84369[1];
  assign array_update_84382[2] = add_84176 == 32'h0000_0002 ? array_update_84380 : array_update_84369[2];
  assign array_update_84382[3] = add_84176 == 32'h0000_0003 ? array_update_84380 : array_update_84369[3];
  assign array_update_84382[4] = add_84176 == 32'h0000_0004 ? array_update_84380 : array_update_84369[4];
  assign array_update_84382[5] = add_84176 == 32'h0000_0005 ? array_update_84380 : array_update_84369[5];
  assign array_update_84382[6] = add_84176 == 32'h0000_0006 ? array_update_84380 : array_update_84369[6];
  assign array_update_84382[7] = add_84176 == 32'h0000_0007 ? array_update_84380 : array_update_84369[7];
  assign array_update_84382[8] = add_84176 == 32'h0000_0008 ? array_update_84380 : array_update_84369[8];
  assign array_update_84382[9] = add_84176 == 32'h0000_0009 ? array_update_84380 : array_update_84369[9];
  assign array_index_84384 = array_update_72021[add_84381 > 32'h0000_0009 ? 4'h9 : add_84381[3:0]];
  assign array_index_84385 = array_update_84382[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_84389 = smul32b_32b_x_32b(array_index_84183[add_84381 > 32'h0000_0009 ? 4'h9 : add_84381[3:0]], array_index_84384[add_84314 > 32'h0000_0009 ? 4'h9 : add_84314[3:0]]);
  assign add_84391 = array_index_84385[add_84314 > 32'h0000_0009 ? 4'h9 : add_84314[3:0]] + smul_84389;
  assign array_update_84393[0] = add_84314 == 32'h0000_0000 ? add_84391 : array_index_84385[0];
  assign array_update_84393[1] = add_84314 == 32'h0000_0001 ? add_84391 : array_index_84385[1];
  assign array_update_84393[2] = add_84314 == 32'h0000_0002 ? add_84391 : array_index_84385[2];
  assign array_update_84393[3] = add_84314 == 32'h0000_0003 ? add_84391 : array_index_84385[3];
  assign array_update_84393[4] = add_84314 == 32'h0000_0004 ? add_84391 : array_index_84385[4];
  assign array_update_84393[5] = add_84314 == 32'h0000_0005 ? add_84391 : array_index_84385[5];
  assign array_update_84393[6] = add_84314 == 32'h0000_0006 ? add_84391 : array_index_84385[6];
  assign array_update_84393[7] = add_84314 == 32'h0000_0007 ? add_84391 : array_index_84385[7];
  assign array_update_84393[8] = add_84314 == 32'h0000_0008 ? add_84391 : array_index_84385[8];
  assign array_update_84393[9] = add_84314 == 32'h0000_0009 ? add_84391 : array_index_84385[9];
  assign add_84394 = add_84381 + 32'h0000_0001;
  assign array_update_84395[0] = add_84176 == 32'h0000_0000 ? array_update_84393 : array_update_84382[0];
  assign array_update_84395[1] = add_84176 == 32'h0000_0001 ? array_update_84393 : array_update_84382[1];
  assign array_update_84395[2] = add_84176 == 32'h0000_0002 ? array_update_84393 : array_update_84382[2];
  assign array_update_84395[3] = add_84176 == 32'h0000_0003 ? array_update_84393 : array_update_84382[3];
  assign array_update_84395[4] = add_84176 == 32'h0000_0004 ? array_update_84393 : array_update_84382[4];
  assign array_update_84395[5] = add_84176 == 32'h0000_0005 ? array_update_84393 : array_update_84382[5];
  assign array_update_84395[6] = add_84176 == 32'h0000_0006 ? array_update_84393 : array_update_84382[6];
  assign array_update_84395[7] = add_84176 == 32'h0000_0007 ? array_update_84393 : array_update_84382[7];
  assign array_update_84395[8] = add_84176 == 32'h0000_0008 ? array_update_84393 : array_update_84382[8];
  assign array_update_84395[9] = add_84176 == 32'h0000_0009 ? array_update_84393 : array_update_84382[9];
  assign array_index_84397 = array_update_72021[add_84394 > 32'h0000_0009 ? 4'h9 : add_84394[3:0]];
  assign array_index_84398 = array_update_84395[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_84402 = smul32b_32b_x_32b(array_index_84183[add_84394 > 32'h0000_0009 ? 4'h9 : add_84394[3:0]], array_index_84397[add_84314 > 32'h0000_0009 ? 4'h9 : add_84314[3:0]]);
  assign add_84404 = array_index_84398[add_84314 > 32'h0000_0009 ? 4'h9 : add_84314[3:0]] + smul_84402;
  assign array_update_84406[0] = add_84314 == 32'h0000_0000 ? add_84404 : array_index_84398[0];
  assign array_update_84406[1] = add_84314 == 32'h0000_0001 ? add_84404 : array_index_84398[1];
  assign array_update_84406[2] = add_84314 == 32'h0000_0002 ? add_84404 : array_index_84398[2];
  assign array_update_84406[3] = add_84314 == 32'h0000_0003 ? add_84404 : array_index_84398[3];
  assign array_update_84406[4] = add_84314 == 32'h0000_0004 ? add_84404 : array_index_84398[4];
  assign array_update_84406[5] = add_84314 == 32'h0000_0005 ? add_84404 : array_index_84398[5];
  assign array_update_84406[6] = add_84314 == 32'h0000_0006 ? add_84404 : array_index_84398[6];
  assign array_update_84406[7] = add_84314 == 32'h0000_0007 ? add_84404 : array_index_84398[7];
  assign array_update_84406[8] = add_84314 == 32'h0000_0008 ? add_84404 : array_index_84398[8];
  assign array_update_84406[9] = add_84314 == 32'h0000_0009 ? add_84404 : array_index_84398[9];
  assign add_84407 = add_84394 + 32'h0000_0001;
  assign array_update_84408[0] = add_84176 == 32'h0000_0000 ? array_update_84406 : array_update_84395[0];
  assign array_update_84408[1] = add_84176 == 32'h0000_0001 ? array_update_84406 : array_update_84395[1];
  assign array_update_84408[2] = add_84176 == 32'h0000_0002 ? array_update_84406 : array_update_84395[2];
  assign array_update_84408[3] = add_84176 == 32'h0000_0003 ? array_update_84406 : array_update_84395[3];
  assign array_update_84408[4] = add_84176 == 32'h0000_0004 ? array_update_84406 : array_update_84395[4];
  assign array_update_84408[5] = add_84176 == 32'h0000_0005 ? array_update_84406 : array_update_84395[5];
  assign array_update_84408[6] = add_84176 == 32'h0000_0006 ? array_update_84406 : array_update_84395[6];
  assign array_update_84408[7] = add_84176 == 32'h0000_0007 ? array_update_84406 : array_update_84395[7];
  assign array_update_84408[8] = add_84176 == 32'h0000_0008 ? array_update_84406 : array_update_84395[8];
  assign array_update_84408[9] = add_84176 == 32'h0000_0009 ? array_update_84406 : array_update_84395[9];
  assign array_index_84410 = array_update_72021[add_84407 > 32'h0000_0009 ? 4'h9 : add_84407[3:0]];
  assign array_index_84411 = array_update_84408[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_84415 = smul32b_32b_x_32b(array_index_84183[add_84407 > 32'h0000_0009 ? 4'h9 : add_84407[3:0]], array_index_84410[add_84314 > 32'h0000_0009 ? 4'h9 : add_84314[3:0]]);
  assign add_84417 = array_index_84411[add_84314 > 32'h0000_0009 ? 4'h9 : add_84314[3:0]] + smul_84415;
  assign array_update_84419[0] = add_84314 == 32'h0000_0000 ? add_84417 : array_index_84411[0];
  assign array_update_84419[1] = add_84314 == 32'h0000_0001 ? add_84417 : array_index_84411[1];
  assign array_update_84419[2] = add_84314 == 32'h0000_0002 ? add_84417 : array_index_84411[2];
  assign array_update_84419[3] = add_84314 == 32'h0000_0003 ? add_84417 : array_index_84411[3];
  assign array_update_84419[4] = add_84314 == 32'h0000_0004 ? add_84417 : array_index_84411[4];
  assign array_update_84419[5] = add_84314 == 32'h0000_0005 ? add_84417 : array_index_84411[5];
  assign array_update_84419[6] = add_84314 == 32'h0000_0006 ? add_84417 : array_index_84411[6];
  assign array_update_84419[7] = add_84314 == 32'h0000_0007 ? add_84417 : array_index_84411[7];
  assign array_update_84419[8] = add_84314 == 32'h0000_0008 ? add_84417 : array_index_84411[8];
  assign array_update_84419[9] = add_84314 == 32'h0000_0009 ? add_84417 : array_index_84411[9];
  assign add_84420 = add_84407 + 32'h0000_0001;
  assign array_update_84421[0] = add_84176 == 32'h0000_0000 ? array_update_84419 : array_update_84408[0];
  assign array_update_84421[1] = add_84176 == 32'h0000_0001 ? array_update_84419 : array_update_84408[1];
  assign array_update_84421[2] = add_84176 == 32'h0000_0002 ? array_update_84419 : array_update_84408[2];
  assign array_update_84421[3] = add_84176 == 32'h0000_0003 ? array_update_84419 : array_update_84408[3];
  assign array_update_84421[4] = add_84176 == 32'h0000_0004 ? array_update_84419 : array_update_84408[4];
  assign array_update_84421[5] = add_84176 == 32'h0000_0005 ? array_update_84419 : array_update_84408[5];
  assign array_update_84421[6] = add_84176 == 32'h0000_0006 ? array_update_84419 : array_update_84408[6];
  assign array_update_84421[7] = add_84176 == 32'h0000_0007 ? array_update_84419 : array_update_84408[7];
  assign array_update_84421[8] = add_84176 == 32'h0000_0008 ? array_update_84419 : array_update_84408[8];
  assign array_update_84421[9] = add_84176 == 32'h0000_0009 ? array_update_84419 : array_update_84408[9];
  assign array_index_84423 = array_update_72021[add_84420 > 32'h0000_0009 ? 4'h9 : add_84420[3:0]];
  assign array_index_84424 = array_update_84421[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_84428 = smul32b_32b_x_32b(array_index_84183[add_84420 > 32'h0000_0009 ? 4'h9 : add_84420[3:0]], array_index_84423[add_84314 > 32'h0000_0009 ? 4'h9 : add_84314[3:0]]);
  assign add_84430 = array_index_84424[add_84314 > 32'h0000_0009 ? 4'h9 : add_84314[3:0]] + smul_84428;
  assign array_update_84432[0] = add_84314 == 32'h0000_0000 ? add_84430 : array_index_84424[0];
  assign array_update_84432[1] = add_84314 == 32'h0000_0001 ? add_84430 : array_index_84424[1];
  assign array_update_84432[2] = add_84314 == 32'h0000_0002 ? add_84430 : array_index_84424[2];
  assign array_update_84432[3] = add_84314 == 32'h0000_0003 ? add_84430 : array_index_84424[3];
  assign array_update_84432[4] = add_84314 == 32'h0000_0004 ? add_84430 : array_index_84424[4];
  assign array_update_84432[5] = add_84314 == 32'h0000_0005 ? add_84430 : array_index_84424[5];
  assign array_update_84432[6] = add_84314 == 32'h0000_0006 ? add_84430 : array_index_84424[6];
  assign array_update_84432[7] = add_84314 == 32'h0000_0007 ? add_84430 : array_index_84424[7];
  assign array_update_84432[8] = add_84314 == 32'h0000_0008 ? add_84430 : array_index_84424[8];
  assign array_update_84432[9] = add_84314 == 32'h0000_0009 ? add_84430 : array_index_84424[9];
  assign add_84433 = add_84420 + 32'h0000_0001;
  assign array_update_84434[0] = add_84176 == 32'h0000_0000 ? array_update_84432 : array_update_84421[0];
  assign array_update_84434[1] = add_84176 == 32'h0000_0001 ? array_update_84432 : array_update_84421[1];
  assign array_update_84434[2] = add_84176 == 32'h0000_0002 ? array_update_84432 : array_update_84421[2];
  assign array_update_84434[3] = add_84176 == 32'h0000_0003 ? array_update_84432 : array_update_84421[3];
  assign array_update_84434[4] = add_84176 == 32'h0000_0004 ? array_update_84432 : array_update_84421[4];
  assign array_update_84434[5] = add_84176 == 32'h0000_0005 ? array_update_84432 : array_update_84421[5];
  assign array_update_84434[6] = add_84176 == 32'h0000_0006 ? array_update_84432 : array_update_84421[6];
  assign array_update_84434[7] = add_84176 == 32'h0000_0007 ? array_update_84432 : array_update_84421[7];
  assign array_update_84434[8] = add_84176 == 32'h0000_0008 ? array_update_84432 : array_update_84421[8];
  assign array_update_84434[9] = add_84176 == 32'h0000_0009 ? array_update_84432 : array_update_84421[9];
  assign array_index_84436 = array_update_72021[add_84433 > 32'h0000_0009 ? 4'h9 : add_84433[3:0]];
  assign array_index_84437 = array_update_84434[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_84441 = smul32b_32b_x_32b(array_index_84183[add_84433 > 32'h0000_0009 ? 4'h9 : add_84433[3:0]], array_index_84436[add_84314 > 32'h0000_0009 ? 4'h9 : add_84314[3:0]]);
  assign add_84443 = array_index_84437[add_84314 > 32'h0000_0009 ? 4'h9 : add_84314[3:0]] + smul_84441;
  assign array_update_84444[0] = add_84314 == 32'h0000_0000 ? add_84443 : array_index_84437[0];
  assign array_update_84444[1] = add_84314 == 32'h0000_0001 ? add_84443 : array_index_84437[1];
  assign array_update_84444[2] = add_84314 == 32'h0000_0002 ? add_84443 : array_index_84437[2];
  assign array_update_84444[3] = add_84314 == 32'h0000_0003 ? add_84443 : array_index_84437[3];
  assign array_update_84444[4] = add_84314 == 32'h0000_0004 ? add_84443 : array_index_84437[4];
  assign array_update_84444[5] = add_84314 == 32'h0000_0005 ? add_84443 : array_index_84437[5];
  assign array_update_84444[6] = add_84314 == 32'h0000_0006 ? add_84443 : array_index_84437[6];
  assign array_update_84444[7] = add_84314 == 32'h0000_0007 ? add_84443 : array_index_84437[7];
  assign array_update_84444[8] = add_84314 == 32'h0000_0008 ? add_84443 : array_index_84437[8];
  assign array_update_84444[9] = add_84314 == 32'h0000_0009 ? add_84443 : array_index_84437[9];
  assign array_update_84445[0] = add_84176 == 32'h0000_0000 ? array_update_84444 : array_update_84434[0];
  assign array_update_84445[1] = add_84176 == 32'h0000_0001 ? array_update_84444 : array_update_84434[1];
  assign array_update_84445[2] = add_84176 == 32'h0000_0002 ? array_update_84444 : array_update_84434[2];
  assign array_update_84445[3] = add_84176 == 32'h0000_0003 ? array_update_84444 : array_update_84434[3];
  assign array_update_84445[4] = add_84176 == 32'h0000_0004 ? array_update_84444 : array_update_84434[4];
  assign array_update_84445[5] = add_84176 == 32'h0000_0005 ? array_update_84444 : array_update_84434[5];
  assign array_update_84445[6] = add_84176 == 32'h0000_0006 ? array_update_84444 : array_update_84434[6];
  assign array_update_84445[7] = add_84176 == 32'h0000_0007 ? array_update_84444 : array_update_84434[7];
  assign array_update_84445[8] = add_84176 == 32'h0000_0008 ? array_update_84444 : array_update_84434[8];
  assign array_update_84445[9] = add_84176 == 32'h0000_0009 ? array_update_84444 : array_update_84434[9];
  assign array_index_84447 = array_update_84445[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign add_84449 = add_84314 + 32'h0000_0001;
  assign array_update_84450[0] = add_84449 == 32'h0000_0000 ? 32'h0000_0000 : array_index_84447[0];
  assign array_update_84450[1] = add_84449 == 32'h0000_0001 ? 32'h0000_0000 : array_index_84447[1];
  assign array_update_84450[2] = add_84449 == 32'h0000_0002 ? 32'h0000_0000 : array_index_84447[2];
  assign array_update_84450[3] = add_84449 == 32'h0000_0003 ? 32'h0000_0000 : array_index_84447[3];
  assign array_update_84450[4] = add_84449 == 32'h0000_0004 ? 32'h0000_0000 : array_index_84447[4];
  assign array_update_84450[5] = add_84449 == 32'h0000_0005 ? 32'h0000_0000 : array_index_84447[5];
  assign array_update_84450[6] = add_84449 == 32'h0000_0006 ? 32'h0000_0000 : array_index_84447[6];
  assign array_update_84450[7] = add_84449 == 32'h0000_0007 ? 32'h0000_0000 : array_index_84447[7];
  assign array_update_84450[8] = add_84449 == 32'h0000_0008 ? 32'h0000_0000 : array_index_84447[8];
  assign array_update_84450[9] = add_84449 == 32'h0000_0009 ? 32'h0000_0000 : array_index_84447[9];
  assign literal_84451 = 32'h0000_0000;
  assign array_update_84452[0] = add_84176 == 32'h0000_0000 ? array_update_84450 : array_update_84445[0];
  assign array_update_84452[1] = add_84176 == 32'h0000_0001 ? array_update_84450 : array_update_84445[1];
  assign array_update_84452[2] = add_84176 == 32'h0000_0002 ? array_update_84450 : array_update_84445[2];
  assign array_update_84452[3] = add_84176 == 32'h0000_0003 ? array_update_84450 : array_update_84445[3];
  assign array_update_84452[4] = add_84176 == 32'h0000_0004 ? array_update_84450 : array_update_84445[4];
  assign array_update_84452[5] = add_84176 == 32'h0000_0005 ? array_update_84450 : array_update_84445[5];
  assign array_update_84452[6] = add_84176 == 32'h0000_0006 ? array_update_84450 : array_update_84445[6];
  assign array_update_84452[7] = add_84176 == 32'h0000_0007 ? array_update_84450 : array_update_84445[7];
  assign array_update_84452[8] = add_84176 == 32'h0000_0008 ? array_update_84450 : array_update_84445[8];
  assign array_update_84452[9] = add_84176 == 32'h0000_0009 ? array_update_84450 : array_update_84445[9];
  assign array_index_84454 = array_update_72021[literal_84451 > 32'h0000_0009 ? 4'h9 : literal_84451[3:0]];
  assign array_index_84455 = array_update_84452[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_84459 = smul32b_32b_x_32b(array_index_84183[literal_84451 > 32'h0000_0009 ? 4'h9 : literal_84451[3:0]], array_index_84454[add_84449 > 32'h0000_0009 ? 4'h9 : add_84449[3:0]]);
  assign add_84461 = array_index_84455[add_84449 > 32'h0000_0009 ? 4'h9 : add_84449[3:0]] + smul_84459;
  assign array_update_84463[0] = add_84449 == 32'h0000_0000 ? add_84461 : array_index_84455[0];
  assign array_update_84463[1] = add_84449 == 32'h0000_0001 ? add_84461 : array_index_84455[1];
  assign array_update_84463[2] = add_84449 == 32'h0000_0002 ? add_84461 : array_index_84455[2];
  assign array_update_84463[3] = add_84449 == 32'h0000_0003 ? add_84461 : array_index_84455[3];
  assign array_update_84463[4] = add_84449 == 32'h0000_0004 ? add_84461 : array_index_84455[4];
  assign array_update_84463[5] = add_84449 == 32'h0000_0005 ? add_84461 : array_index_84455[5];
  assign array_update_84463[6] = add_84449 == 32'h0000_0006 ? add_84461 : array_index_84455[6];
  assign array_update_84463[7] = add_84449 == 32'h0000_0007 ? add_84461 : array_index_84455[7];
  assign array_update_84463[8] = add_84449 == 32'h0000_0008 ? add_84461 : array_index_84455[8];
  assign array_update_84463[9] = add_84449 == 32'h0000_0009 ? add_84461 : array_index_84455[9];
  assign add_84464 = literal_84451 + 32'h0000_0001;
  assign array_update_84465[0] = add_84176 == 32'h0000_0000 ? array_update_84463 : array_update_84452[0];
  assign array_update_84465[1] = add_84176 == 32'h0000_0001 ? array_update_84463 : array_update_84452[1];
  assign array_update_84465[2] = add_84176 == 32'h0000_0002 ? array_update_84463 : array_update_84452[2];
  assign array_update_84465[3] = add_84176 == 32'h0000_0003 ? array_update_84463 : array_update_84452[3];
  assign array_update_84465[4] = add_84176 == 32'h0000_0004 ? array_update_84463 : array_update_84452[4];
  assign array_update_84465[5] = add_84176 == 32'h0000_0005 ? array_update_84463 : array_update_84452[5];
  assign array_update_84465[6] = add_84176 == 32'h0000_0006 ? array_update_84463 : array_update_84452[6];
  assign array_update_84465[7] = add_84176 == 32'h0000_0007 ? array_update_84463 : array_update_84452[7];
  assign array_update_84465[8] = add_84176 == 32'h0000_0008 ? array_update_84463 : array_update_84452[8];
  assign array_update_84465[9] = add_84176 == 32'h0000_0009 ? array_update_84463 : array_update_84452[9];
  assign array_index_84467 = array_update_72021[add_84464 > 32'h0000_0009 ? 4'h9 : add_84464[3:0]];
  assign array_index_84468 = array_update_84465[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_84472 = smul32b_32b_x_32b(array_index_84183[add_84464 > 32'h0000_0009 ? 4'h9 : add_84464[3:0]], array_index_84467[add_84449 > 32'h0000_0009 ? 4'h9 : add_84449[3:0]]);
  assign add_84474 = array_index_84468[add_84449 > 32'h0000_0009 ? 4'h9 : add_84449[3:0]] + smul_84472;
  assign array_update_84476[0] = add_84449 == 32'h0000_0000 ? add_84474 : array_index_84468[0];
  assign array_update_84476[1] = add_84449 == 32'h0000_0001 ? add_84474 : array_index_84468[1];
  assign array_update_84476[2] = add_84449 == 32'h0000_0002 ? add_84474 : array_index_84468[2];
  assign array_update_84476[3] = add_84449 == 32'h0000_0003 ? add_84474 : array_index_84468[3];
  assign array_update_84476[4] = add_84449 == 32'h0000_0004 ? add_84474 : array_index_84468[4];
  assign array_update_84476[5] = add_84449 == 32'h0000_0005 ? add_84474 : array_index_84468[5];
  assign array_update_84476[6] = add_84449 == 32'h0000_0006 ? add_84474 : array_index_84468[6];
  assign array_update_84476[7] = add_84449 == 32'h0000_0007 ? add_84474 : array_index_84468[7];
  assign array_update_84476[8] = add_84449 == 32'h0000_0008 ? add_84474 : array_index_84468[8];
  assign array_update_84476[9] = add_84449 == 32'h0000_0009 ? add_84474 : array_index_84468[9];
  assign add_84477 = add_84464 + 32'h0000_0001;
  assign array_update_84478[0] = add_84176 == 32'h0000_0000 ? array_update_84476 : array_update_84465[0];
  assign array_update_84478[1] = add_84176 == 32'h0000_0001 ? array_update_84476 : array_update_84465[1];
  assign array_update_84478[2] = add_84176 == 32'h0000_0002 ? array_update_84476 : array_update_84465[2];
  assign array_update_84478[3] = add_84176 == 32'h0000_0003 ? array_update_84476 : array_update_84465[3];
  assign array_update_84478[4] = add_84176 == 32'h0000_0004 ? array_update_84476 : array_update_84465[4];
  assign array_update_84478[5] = add_84176 == 32'h0000_0005 ? array_update_84476 : array_update_84465[5];
  assign array_update_84478[6] = add_84176 == 32'h0000_0006 ? array_update_84476 : array_update_84465[6];
  assign array_update_84478[7] = add_84176 == 32'h0000_0007 ? array_update_84476 : array_update_84465[7];
  assign array_update_84478[8] = add_84176 == 32'h0000_0008 ? array_update_84476 : array_update_84465[8];
  assign array_update_84478[9] = add_84176 == 32'h0000_0009 ? array_update_84476 : array_update_84465[9];
  assign array_index_84480 = array_update_72021[add_84477 > 32'h0000_0009 ? 4'h9 : add_84477[3:0]];
  assign array_index_84481 = array_update_84478[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_84485 = smul32b_32b_x_32b(array_index_84183[add_84477 > 32'h0000_0009 ? 4'h9 : add_84477[3:0]], array_index_84480[add_84449 > 32'h0000_0009 ? 4'h9 : add_84449[3:0]]);
  assign add_84487 = array_index_84481[add_84449 > 32'h0000_0009 ? 4'h9 : add_84449[3:0]] + smul_84485;
  assign array_update_84489[0] = add_84449 == 32'h0000_0000 ? add_84487 : array_index_84481[0];
  assign array_update_84489[1] = add_84449 == 32'h0000_0001 ? add_84487 : array_index_84481[1];
  assign array_update_84489[2] = add_84449 == 32'h0000_0002 ? add_84487 : array_index_84481[2];
  assign array_update_84489[3] = add_84449 == 32'h0000_0003 ? add_84487 : array_index_84481[3];
  assign array_update_84489[4] = add_84449 == 32'h0000_0004 ? add_84487 : array_index_84481[4];
  assign array_update_84489[5] = add_84449 == 32'h0000_0005 ? add_84487 : array_index_84481[5];
  assign array_update_84489[6] = add_84449 == 32'h0000_0006 ? add_84487 : array_index_84481[6];
  assign array_update_84489[7] = add_84449 == 32'h0000_0007 ? add_84487 : array_index_84481[7];
  assign array_update_84489[8] = add_84449 == 32'h0000_0008 ? add_84487 : array_index_84481[8];
  assign array_update_84489[9] = add_84449 == 32'h0000_0009 ? add_84487 : array_index_84481[9];
  assign add_84490 = add_84477 + 32'h0000_0001;
  assign array_update_84491[0] = add_84176 == 32'h0000_0000 ? array_update_84489 : array_update_84478[0];
  assign array_update_84491[1] = add_84176 == 32'h0000_0001 ? array_update_84489 : array_update_84478[1];
  assign array_update_84491[2] = add_84176 == 32'h0000_0002 ? array_update_84489 : array_update_84478[2];
  assign array_update_84491[3] = add_84176 == 32'h0000_0003 ? array_update_84489 : array_update_84478[3];
  assign array_update_84491[4] = add_84176 == 32'h0000_0004 ? array_update_84489 : array_update_84478[4];
  assign array_update_84491[5] = add_84176 == 32'h0000_0005 ? array_update_84489 : array_update_84478[5];
  assign array_update_84491[6] = add_84176 == 32'h0000_0006 ? array_update_84489 : array_update_84478[6];
  assign array_update_84491[7] = add_84176 == 32'h0000_0007 ? array_update_84489 : array_update_84478[7];
  assign array_update_84491[8] = add_84176 == 32'h0000_0008 ? array_update_84489 : array_update_84478[8];
  assign array_update_84491[9] = add_84176 == 32'h0000_0009 ? array_update_84489 : array_update_84478[9];
  assign array_index_84493 = array_update_72021[add_84490 > 32'h0000_0009 ? 4'h9 : add_84490[3:0]];
  assign array_index_84494 = array_update_84491[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_84498 = smul32b_32b_x_32b(array_index_84183[add_84490 > 32'h0000_0009 ? 4'h9 : add_84490[3:0]], array_index_84493[add_84449 > 32'h0000_0009 ? 4'h9 : add_84449[3:0]]);
  assign add_84500 = array_index_84494[add_84449 > 32'h0000_0009 ? 4'h9 : add_84449[3:0]] + smul_84498;
  assign array_update_84502[0] = add_84449 == 32'h0000_0000 ? add_84500 : array_index_84494[0];
  assign array_update_84502[1] = add_84449 == 32'h0000_0001 ? add_84500 : array_index_84494[1];
  assign array_update_84502[2] = add_84449 == 32'h0000_0002 ? add_84500 : array_index_84494[2];
  assign array_update_84502[3] = add_84449 == 32'h0000_0003 ? add_84500 : array_index_84494[3];
  assign array_update_84502[4] = add_84449 == 32'h0000_0004 ? add_84500 : array_index_84494[4];
  assign array_update_84502[5] = add_84449 == 32'h0000_0005 ? add_84500 : array_index_84494[5];
  assign array_update_84502[6] = add_84449 == 32'h0000_0006 ? add_84500 : array_index_84494[6];
  assign array_update_84502[7] = add_84449 == 32'h0000_0007 ? add_84500 : array_index_84494[7];
  assign array_update_84502[8] = add_84449 == 32'h0000_0008 ? add_84500 : array_index_84494[8];
  assign array_update_84502[9] = add_84449 == 32'h0000_0009 ? add_84500 : array_index_84494[9];
  assign add_84503 = add_84490 + 32'h0000_0001;
  assign array_update_84504[0] = add_84176 == 32'h0000_0000 ? array_update_84502 : array_update_84491[0];
  assign array_update_84504[1] = add_84176 == 32'h0000_0001 ? array_update_84502 : array_update_84491[1];
  assign array_update_84504[2] = add_84176 == 32'h0000_0002 ? array_update_84502 : array_update_84491[2];
  assign array_update_84504[3] = add_84176 == 32'h0000_0003 ? array_update_84502 : array_update_84491[3];
  assign array_update_84504[4] = add_84176 == 32'h0000_0004 ? array_update_84502 : array_update_84491[4];
  assign array_update_84504[5] = add_84176 == 32'h0000_0005 ? array_update_84502 : array_update_84491[5];
  assign array_update_84504[6] = add_84176 == 32'h0000_0006 ? array_update_84502 : array_update_84491[6];
  assign array_update_84504[7] = add_84176 == 32'h0000_0007 ? array_update_84502 : array_update_84491[7];
  assign array_update_84504[8] = add_84176 == 32'h0000_0008 ? array_update_84502 : array_update_84491[8];
  assign array_update_84504[9] = add_84176 == 32'h0000_0009 ? array_update_84502 : array_update_84491[9];
  assign array_index_84506 = array_update_72021[add_84503 > 32'h0000_0009 ? 4'h9 : add_84503[3:0]];
  assign array_index_84507 = array_update_84504[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_84511 = smul32b_32b_x_32b(array_index_84183[add_84503 > 32'h0000_0009 ? 4'h9 : add_84503[3:0]], array_index_84506[add_84449 > 32'h0000_0009 ? 4'h9 : add_84449[3:0]]);
  assign add_84513 = array_index_84507[add_84449 > 32'h0000_0009 ? 4'h9 : add_84449[3:0]] + smul_84511;
  assign array_update_84515[0] = add_84449 == 32'h0000_0000 ? add_84513 : array_index_84507[0];
  assign array_update_84515[1] = add_84449 == 32'h0000_0001 ? add_84513 : array_index_84507[1];
  assign array_update_84515[2] = add_84449 == 32'h0000_0002 ? add_84513 : array_index_84507[2];
  assign array_update_84515[3] = add_84449 == 32'h0000_0003 ? add_84513 : array_index_84507[3];
  assign array_update_84515[4] = add_84449 == 32'h0000_0004 ? add_84513 : array_index_84507[4];
  assign array_update_84515[5] = add_84449 == 32'h0000_0005 ? add_84513 : array_index_84507[5];
  assign array_update_84515[6] = add_84449 == 32'h0000_0006 ? add_84513 : array_index_84507[6];
  assign array_update_84515[7] = add_84449 == 32'h0000_0007 ? add_84513 : array_index_84507[7];
  assign array_update_84515[8] = add_84449 == 32'h0000_0008 ? add_84513 : array_index_84507[8];
  assign array_update_84515[9] = add_84449 == 32'h0000_0009 ? add_84513 : array_index_84507[9];
  assign add_84516 = add_84503 + 32'h0000_0001;
  assign array_update_84517[0] = add_84176 == 32'h0000_0000 ? array_update_84515 : array_update_84504[0];
  assign array_update_84517[1] = add_84176 == 32'h0000_0001 ? array_update_84515 : array_update_84504[1];
  assign array_update_84517[2] = add_84176 == 32'h0000_0002 ? array_update_84515 : array_update_84504[2];
  assign array_update_84517[3] = add_84176 == 32'h0000_0003 ? array_update_84515 : array_update_84504[3];
  assign array_update_84517[4] = add_84176 == 32'h0000_0004 ? array_update_84515 : array_update_84504[4];
  assign array_update_84517[5] = add_84176 == 32'h0000_0005 ? array_update_84515 : array_update_84504[5];
  assign array_update_84517[6] = add_84176 == 32'h0000_0006 ? array_update_84515 : array_update_84504[6];
  assign array_update_84517[7] = add_84176 == 32'h0000_0007 ? array_update_84515 : array_update_84504[7];
  assign array_update_84517[8] = add_84176 == 32'h0000_0008 ? array_update_84515 : array_update_84504[8];
  assign array_update_84517[9] = add_84176 == 32'h0000_0009 ? array_update_84515 : array_update_84504[9];
  assign array_index_84519 = array_update_72021[add_84516 > 32'h0000_0009 ? 4'h9 : add_84516[3:0]];
  assign array_index_84520 = array_update_84517[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_84524 = smul32b_32b_x_32b(array_index_84183[add_84516 > 32'h0000_0009 ? 4'h9 : add_84516[3:0]], array_index_84519[add_84449 > 32'h0000_0009 ? 4'h9 : add_84449[3:0]]);
  assign add_84526 = array_index_84520[add_84449 > 32'h0000_0009 ? 4'h9 : add_84449[3:0]] + smul_84524;
  assign array_update_84528[0] = add_84449 == 32'h0000_0000 ? add_84526 : array_index_84520[0];
  assign array_update_84528[1] = add_84449 == 32'h0000_0001 ? add_84526 : array_index_84520[1];
  assign array_update_84528[2] = add_84449 == 32'h0000_0002 ? add_84526 : array_index_84520[2];
  assign array_update_84528[3] = add_84449 == 32'h0000_0003 ? add_84526 : array_index_84520[3];
  assign array_update_84528[4] = add_84449 == 32'h0000_0004 ? add_84526 : array_index_84520[4];
  assign array_update_84528[5] = add_84449 == 32'h0000_0005 ? add_84526 : array_index_84520[5];
  assign array_update_84528[6] = add_84449 == 32'h0000_0006 ? add_84526 : array_index_84520[6];
  assign array_update_84528[7] = add_84449 == 32'h0000_0007 ? add_84526 : array_index_84520[7];
  assign array_update_84528[8] = add_84449 == 32'h0000_0008 ? add_84526 : array_index_84520[8];
  assign array_update_84528[9] = add_84449 == 32'h0000_0009 ? add_84526 : array_index_84520[9];
  assign add_84529 = add_84516 + 32'h0000_0001;
  assign array_update_84530[0] = add_84176 == 32'h0000_0000 ? array_update_84528 : array_update_84517[0];
  assign array_update_84530[1] = add_84176 == 32'h0000_0001 ? array_update_84528 : array_update_84517[1];
  assign array_update_84530[2] = add_84176 == 32'h0000_0002 ? array_update_84528 : array_update_84517[2];
  assign array_update_84530[3] = add_84176 == 32'h0000_0003 ? array_update_84528 : array_update_84517[3];
  assign array_update_84530[4] = add_84176 == 32'h0000_0004 ? array_update_84528 : array_update_84517[4];
  assign array_update_84530[5] = add_84176 == 32'h0000_0005 ? array_update_84528 : array_update_84517[5];
  assign array_update_84530[6] = add_84176 == 32'h0000_0006 ? array_update_84528 : array_update_84517[6];
  assign array_update_84530[7] = add_84176 == 32'h0000_0007 ? array_update_84528 : array_update_84517[7];
  assign array_update_84530[8] = add_84176 == 32'h0000_0008 ? array_update_84528 : array_update_84517[8];
  assign array_update_84530[9] = add_84176 == 32'h0000_0009 ? array_update_84528 : array_update_84517[9];
  assign array_index_84532 = array_update_72021[add_84529 > 32'h0000_0009 ? 4'h9 : add_84529[3:0]];
  assign array_index_84533 = array_update_84530[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_84537 = smul32b_32b_x_32b(array_index_84183[add_84529 > 32'h0000_0009 ? 4'h9 : add_84529[3:0]], array_index_84532[add_84449 > 32'h0000_0009 ? 4'h9 : add_84449[3:0]]);
  assign add_84539 = array_index_84533[add_84449 > 32'h0000_0009 ? 4'h9 : add_84449[3:0]] + smul_84537;
  assign array_update_84541[0] = add_84449 == 32'h0000_0000 ? add_84539 : array_index_84533[0];
  assign array_update_84541[1] = add_84449 == 32'h0000_0001 ? add_84539 : array_index_84533[1];
  assign array_update_84541[2] = add_84449 == 32'h0000_0002 ? add_84539 : array_index_84533[2];
  assign array_update_84541[3] = add_84449 == 32'h0000_0003 ? add_84539 : array_index_84533[3];
  assign array_update_84541[4] = add_84449 == 32'h0000_0004 ? add_84539 : array_index_84533[4];
  assign array_update_84541[5] = add_84449 == 32'h0000_0005 ? add_84539 : array_index_84533[5];
  assign array_update_84541[6] = add_84449 == 32'h0000_0006 ? add_84539 : array_index_84533[6];
  assign array_update_84541[7] = add_84449 == 32'h0000_0007 ? add_84539 : array_index_84533[7];
  assign array_update_84541[8] = add_84449 == 32'h0000_0008 ? add_84539 : array_index_84533[8];
  assign array_update_84541[9] = add_84449 == 32'h0000_0009 ? add_84539 : array_index_84533[9];
  assign add_84542 = add_84529 + 32'h0000_0001;
  assign array_update_84543[0] = add_84176 == 32'h0000_0000 ? array_update_84541 : array_update_84530[0];
  assign array_update_84543[1] = add_84176 == 32'h0000_0001 ? array_update_84541 : array_update_84530[1];
  assign array_update_84543[2] = add_84176 == 32'h0000_0002 ? array_update_84541 : array_update_84530[2];
  assign array_update_84543[3] = add_84176 == 32'h0000_0003 ? array_update_84541 : array_update_84530[3];
  assign array_update_84543[4] = add_84176 == 32'h0000_0004 ? array_update_84541 : array_update_84530[4];
  assign array_update_84543[5] = add_84176 == 32'h0000_0005 ? array_update_84541 : array_update_84530[5];
  assign array_update_84543[6] = add_84176 == 32'h0000_0006 ? array_update_84541 : array_update_84530[6];
  assign array_update_84543[7] = add_84176 == 32'h0000_0007 ? array_update_84541 : array_update_84530[7];
  assign array_update_84543[8] = add_84176 == 32'h0000_0008 ? array_update_84541 : array_update_84530[8];
  assign array_update_84543[9] = add_84176 == 32'h0000_0009 ? array_update_84541 : array_update_84530[9];
  assign array_index_84545 = array_update_72021[add_84542 > 32'h0000_0009 ? 4'h9 : add_84542[3:0]];
  assign array_index_84546 = array_update_84543[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_84550 = smul32b_32b_x_32b(array_index_84183[add_84542 > 32'h0000_0009 ? 4'h9 : add_84542[3:0]], array_index_84545[add_84449 > 32'h0000_0009 ? 4'h9 : add_84449[3:0]]);
  assign add_84552 = array_index_84546[add_84449 > 32'h0000_0009 ? 4'h9 : add_84449[3:0]] + smul_84550;
  assign array_update_84554[0] = add_84449 == 32'h0000_0000 ? add_84552 : array_index_84546[0];
  assign array_update_84554[1] = add_84449 == 32'h0000_0001 ? add_84552 : array_index_84546[1];
  assign array_update_84554[2] = add_84449 == 32'h0000_0002 ? add_84552 : array_index_84546[2];
  assign array_update_84554[3] = add_84449 == 32'h0000_0003 ? add_84552 : array_index_84546[3];
  assign array_update_84554[4] = add_84449 == 32'h0000_0004 ? add_84552 : array_index_84546[4];
  assign array_update_84554[5] = add_84449 == 32'h0000_0005 ? add_84552 : array_index_84546[5];
  assign array_update_84554[6] = add_84449 == 32'h0000_0006 ? add_84552 : array_index_84546[6];
  assign array_update_84554[7] = add_84449 == 32'h0000_0007 ? add_84552 : array_index_84546[7];
  assign array_update_84554[8] = add_84449 == 32'h0000_0008 ? add_84552 : array_index_84546[8];
  assign array_update_84554[9] = add_84449 == 32'h0000_0009 ? add_84552 : array_index_84546[9];
  assign add_84555 = add_84542 + 32'h0000_0001;
  assign array_update_84556[0] = add_84176 == 32'h0000_0000 ? array_update_84554 : array_update_84543[0];
  assign array_update_84556[1] = add_84176 == 32'h0000_0001 ? array_update_84554 : array_update_84543[1];
  assign array_update_84556[2] = add_84176 == 32'h0000_0002 ? array_update_84554 : array_update_84543[2];
  assign array_update_84556[3] = add_84176 == 32'h0000_0003 ? array_update_84554 : array_update_84543[3];
  assign array_update_84556[4] = add_84176 == 32'h0000_0004 ? array_update_84554 : array_update_84543[4];
  assign array_update_84556[5] = add_84176 == 32'h0000_0005 ? array_update_84554 : array_update_84543[5];
  assign array_update_84556[6] = add_84176 == 32'h0000_0006 ? array_update_84554 : array_update_84543[6];
  assign array_update_84556[7] = add_84176 == 32'h0000_0007 ? array_update_84554 : array_update_84543[7];
  assign array_update_84556[8] = add_84176 == 32'h0000_0008 ? array_update_84554 : array_update_84543[8];
  assign array_update_84556[9] = add_84176 == 32'h0000_0009 ? array_update_84554 : array_update_84543[9];
  assign array_index_84558 = array_update_72021[add_84555 > 32'h0000_0009 ? 4'h9 : add_84555[3:0]];
  assign array_index_84559 = array_update_84556[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_84563 = smul32b_32b_x_32b(array_index_84183[add_84555 > 32'h0000_0009 ? 4'h9 : add_84555[3:0]], array_index_84558[add_84449 > 32'h0000_0009 ? 4'h9 : add_84449[3:0]]);
  assign add_84565 = array_index_84559[add_84449 > 32'h0000_0009 ? 4'h9 : add_84449[3:0]] + smul_84563;
  assign array_update_84567[0] = add_84449 == 32'h0000_0000 ? add_84565 : array_index_84559[0];
  assign array_update_84567[1] = add_84449 == 32'h0000_0001 ? add_84565 : array_index_84559[1];
  assign array_update_84567[2] = add_84449 == 32'h0000_0002 ? add_84565 : array_index_84559[2];
  assign array_update_84567[3] = add_84449 == 32'h0000_0003 ? add_84565 : array_index_84559[3];
  assign array_update_84567[4] = add_84449 == 32'h0000_0004 ? add_84565 : array_index_84559[4];
  assign array_update_84567[5] = add_84449 == 32'h0000_0005 ? add_84565 : array_index_84559[5];
  assign array_update_84567[6] = add_84449 == 32'h0000_0006 ? add_84565 : array_index_84559[6];
  assign array_update_84567[7] = add_84449 == 32'h0000_0007 ? add_84565 : array_index_84559[7];
  assign array_update_84567[8] = add_84449 == 32'h0000_0008 ? add_84565 : array_index_84559[8];
  assign array_update_84567[9] = add_84449 == 32'h0000_0009 ? add_84565 : array_index_84559[9];
  assign add_84568 = add_84555 + 32'h0000_0001;
  assign array_update_84569[0] = add_84176 == 32'h0000_0000 ? array_update_84567 : array_update_84556[0];
  assign array_update_84569[1] = add_84176 == 32'h0000_0001 ? array_update_84567 : array_update_84556[1];
  assign array_update_84569[2] = add_84176 == 32'h0000_0002 ? array_update_84567 : array_update_84556[2];
  assign array_update_84569[3] = add_84176 == 32'h0000_0003 ? array_update_84567 : array_update_84556[3];
  assign array_update_84569[4] = add_84176 == 32'h0000_0004 ? array_update_84567 : array_update_84556[4];
  assign array_update_84569[5] = add_84176 == 32'h0000_0005 ? array_update_84567 : array_update_84556[5];
  assign array_update_84569[6] = add_84176 == 32'h0000_0006 ? array_update_84567 : array_update_84556[6];
  assign array_update_84569[7] = add_84176 == 32'h0000_0007 ? array_update_84567 : array_update_84556[7];
  assign array_update_84569[8] = add_84176 == 32'h0000_0008 ? array_update_84567 : array_update_84556[8];
  assign array_update_84569[9] = add_84176 == 32'h0000_0009 ? array_update_84567 : array_update_84556[9];
  assign array_index_84571 = array_update_72021[add_84568 > 32'h0000_0009 ? 4'h9 : add_84568[3:0]];
  assign array_index_84572 = array_update_84569[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_84576 = smul32b_32b_x_32b(array_index_84183[add_84568 > 32'h0000_0009 ? 4'h9 : add_84568[3:0]], array_index_84571[add_84449 > 32'h0000_0009 ? 4'h9 : add_84449[3:0]]);
  assign add_84578 = array_index_84572[add_84449 > 32'h0000_0009 ? 4'h9 : add_84449[3:0]] + smul_84576;
  assign array_update_84579[0] = add_84449 == 32'h0000_0000 ? add_84578 : array_index_84572[0];
  assign array_update_84579[1] = add_84449 == 32'h0000_0001 ? add_84578 : array_index_84572[1];
  assign array_update_84579[2] = add_84449 == 32'h0000_0002 ? add_84578 : array_index_84572[2];
  assign array_update_84579[3] = add_84449 == 32'h0000_0003 ? add_84578 : array_index_84572[3];
  assign array_update_84579[4] = add_84449 == 32'h0000_0004 ? add_84578 : array_index_84572[4];
  assign array_update_84579[5] = add_84449 == 32'h0000_0005 ? add_84578 : array_index_84572[5];
  assign array_update_84579[6] = add_84449 == 32'h0000_0006 ? add_84578 : array_index_84572[6];
  assign array_update_84579[7] = add_84449 == 32'h0000_0007 ? add_84578 : array_index_84572[7];
  assign array_update_84579[8] = add_84449 == 32'h0000_0008 ? add_84578 : array_index_84572[8];
  assign array_update_84579[9] = add_84449 == 32'h0000_0009 ? add_84578 : array_index_84572[9];
  assign array_update_84580[0] = add_84176 == 32'h0000_0000 ? array_update_84579 : array_update_84569[0];
  assign array_update_84580[1] = add_84176 == 32'h0000_0001 ? array_update_84579 : array_update_84569[1];
  assign array_update_84580[2] = add_84176 == 32'h0000_0002 ? array_update_84579 : array_update_84569[2];
  assign array_update_84580[3] = add_84176 == 32'h0000_0003 ? array_update_84579 : array_update_84569[3];
  assign array_update_84580[4] = add_84176 == 32'h0000_0004 ? array_update_84579 : array_update_84569[4];
  assign array_update_84580[5] = add_84176 == 32'h0000_0005 ? array_update_84579 : array_update_84569[5];
  assign array_update_84580[6] = add_84176 == 32'h0000_0006 ? array_update_84579 : array_update_84569[6];
  assign array_update_84580[7] = add_84176 == 32'h0000_0007 ? array_update_84579 : array_update_84569[7];
  assign array_update_84580[8] = add_84176 == 32'h0000_0008 ? array_update_84579 : array_update_84569[8];
  assign array_update_84580[9] = add_84176 == 32'h0000_0009 ? array_update_84579 : array_update_84569[9];
  assign array_index_84582 = array_update_84580[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign add_84584 = add_84449 + 32'h0000_0001;
  assign array_update_84585[0] = add_84584 == 32'h0000_0000 ? 32'h0000_0000 : array_index_84582[0];
  assign array_update_84585[1] = add_84584 == 32'h0000_0001 ? 32'h0000_0000 : array_index_84582[1];
  assign array_update_84585[2] = add_84584 == 32'h0000_0002 ? 32'h0000_0000 : array_index_84582[2];
  assign array_update_84585[3] = add_84584 == 32'h0000_0003 ? 32'h0000_0000 : array_index_84582[3];
  assign array_update_84585[4] = add_84584 == 32'h0000_0004 ? 32'h0000_0000 : array_index_84582[4];
  assign array_update_84585[5] = add_84584 == 32'h0000_0005 ? 32'h0000_0000 : array_index_84582[5];
  assign array_update_84585[6] = add_84584 == 32'h0000_0006 ? 32'h0000_0000 : array_index_84582[6];
  assign array_update_84585[7] = add_84584 == 32'h0000_0007 ? 32'h0000_0000 : array_index_84582[7];
  assign array_update_84585[8] = add_84584 == 32'h0000_0008 ? 32'h0000_0000 : array_index_84582[8];
  assign array_update_84585[9] = add_84584 == 32'h0000_0009 ? 32'h0000_0000 : array_index_84582[9];
  assign literal_84586 = 32'h0000_0000;
  assign array_update_84587[0] = add_84176 == 32'h0000_0000 ? array_update_84585 : array_update_84580[0];
  assign array_update_84587[1] = add_84176 == 32'h0000_0001 ? array_update_84585 : array_update_84580[1];
  assign array_update_84587[2] = add_84176 == 32'h0000_0002 ? array_update_84585 : array_update_84580[2];
  assign array_update_84587[3] = add_84176 == 32'h0000_0003 ? array_update_84585 : array_update_84580[3];
  assign array_update_84587[4] = add_84176 == 32'h0000_0004 ? array_update_84585 : array_update_84580[4];
  assign array_update_84587[5] = add_84176 == 32'h0000_0005 ? array_update_84585 : array_update_84580[5];
  assign array_update_84587[6] = add_84176 == 32'h0000_0006 ? array_update_84585 : array_update_84580[6];
  assign array_update_84587[7] = add_84176 == 32'h0000_0007 ? array_update_84585 : array_update_84580[7];
  assign array_update_84587[8] = add_84176 == 32'h0000_0008 ? array_update_84585 : array_update_84580[8];
  assign array_update_84587[9] = add_84176 == 32'h0000_0009 ? array_update_84585 : array_update_84580[9];
  assign array_index_84589 = array_update_72021[literal_84586 > 32'h0000_0009 ? 4'h9 : literal_84586[3:0]];
  assign array_index_84590 = array_update_84587[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_84594 = smul32b_32b_x_32b(array_index_84183[literal_84586 > 32'h0000_0009 ? 4'h9 : literal_84586[3:0]], array_index_84589[add_84584 > 32'h0000_0009 ? 4'h9 : add_84584[3:0]]);
  assign add_84596 = array_index_84590[add_84584 > 32'h0000_0009 ? 4'h9 : add_84584[3:0]] + smul_84594;
  assign array_update_84598[0] = add_84584 == 32'h0000_0000 ? add_84596 : array_index_84590[0];
  assign array_update_84598[1] = add_84584 == 32'h0000_0001 ? add_84596 : array_index_84590[1];
  assign array_update_84598[2] = add_84584 == 32'h0000_0002 ? add_84596 : array_index_84590[2];
  assign array_update_84598[3] = add_84584 == 32'h0000_0003 ? add_84596 : array_index_84590[3];
  assign array_update_84598[4] = add_84584 == 32'h0000_0004 ? add_84596 : array_index_84590[4];
  assign array_update_84598[5] = add_84584 == 32'h0000_0005 ? add_84596 : array_index_84590[5];
  assign array_update_84598[6] = add_84584 == 32'h0000_0006 ? add_84596 : array_index_84590[6];
  assign array_update_84598[7] = add_84584 == 32'h0000_0007 ? add_84596 : array_index_84590[7];
  assign array_update_84598[8] = add_84584 == 32'h0000_0008 ? add_84596 : array_index_84590[8];
  assign array_update_84598[9] = add_84584 == 32'h0000_0009 ? add_84596 : array_index_84590[9];
  assign add_84599 = literal_84586 + 32'h0000_0001;
  assign array_update_84600[0] = add_84176 == 32'h0000_0000 ? array_update_84598 : array_update_84587[0];
  assign array_update_84600[1] = add_84176 == 32'h0000_0001 ? array_update_84598 : array_update_84587[1];
  assign array_update_84600[2] = add_84176 == 32'h0000_0002 ? array_update_84598 : array_update_84587[2];
  assign array_update_84600[3] = add_84176 == 32'h0000_0003 ? array_update_84598 : array_update_84587[3];
  assign array_update_84600[4] = add_84176 == 32'h0000_0004 ? array_update_84598 : array_update_84587[4];
  assign array_update_84600[5] = add_84176 == 32'h0000_0005 ? array_update_84598 : array_update_84587[5];
  assign array_update_84600[6] = add_84176 == 32'h0000_0006 ? array_update_84598 : array_update_84587[6];
  assign array_update_84600[7] = add_84176 == 32'h0000_0007 ? array_update_84598 : array_update_84587[7];
  assign array_update_84600[8] = add_84176 == 32'h0000_0008 ? array_update_84598 : array_update_84587[8];
  assign array_update_84600[9] = add_84176 == 32'h0000_0009 ? array_update_84598 : array_update_84587[9];
  assign array_index_84602 = array_update_72021[add_84599 > 32'h0000_0009 ? 4'h9 : add_84599[3:0]];
  assign array_index_84603 = array_update_84600[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_84607 = smul32b_32b_x_32b(array_index_84183[add_84599 > 32'h0000_0009 ? 4'h9 : add_84599[3:0]], array_index_84602[add_84584 > 32'h0000_0009 ? 4'h9 : add_84584[3:0]]);
  assign add_84609 = array_index_84603[add_84584 > 32'h0000_0009 ? 4'h9 : add_84584[3:0]] + smul_84607;
  assign array_update_84611[0] = add_84584 == 32'h0000_0000 ? add_84609 : array_index_84603[0];
  assign array_update_84611[1] = add_84584 == 32'h0000_0001 ? add_84609 : array_index_84603[1];
  assign array_update_84611[2] = add_84584 == 32'h0000_0002 ? add_84609 : array_index_84603[2];
  assign array_update_84611[3] = add_84584 == 32'h0000_0003 ? add_84609 : array_index_84603[3];
  assign array_update_84611[4] = add_84584 == 32'h0000_0004 ? add_84609 : array_index_84603[4];
  assign array_update_84611[5] = add_84584 == 32'h0000_0005 ? add_84609 : array_index_84603[5];
  assign array_update_84611[6] = add_84584 == 32'h0000_0006 ? add_84609 : array_index_84603[6];
  assign array_update_84611[7] = add_84584 == 32'h0000_0007 ? add_84609 : array_index_84603[7];
  assign array_update_84611[8] = add_84584 == 32'h0000_0008 ? add_84609 : array_index_84603[8];
  assign array_update_84611[9] = add_84584 == 32'h0000_0009 ? add_84609 : array_index_84603[9];
  assign add_84612 = add_84599 + 32'h0000_0001;
  assign array_update_84613[0] = add_84176 == 32'h0000_0000 ? array_update_84611 : array_update_84600[0];
  assign array_update_84613[1] = add_84176 == 32'h0000_0001 ? array_update_84611 : array_update_84600[1];
  assign array_update_84613[2] = add_84176 == 32'h0000_0002 ? array_update_84611 : array_update_84600[2];
  assign array_update_84613[3] = add_84176 == 32'h0000_0003 ? array_update_84611 : array_update_84600[3];
  assign array_update_84613[4] = add_84176 == 32'h0000_0004 ? array_update_84611 : array_update_84600[4];
  assign array_update_84613[5] = add_84176 == 32'h0000_0005 ? array_update_84611 : array_update_84600[5];
  assign array_update_84613[6] = add_84176 == 32'h0000_0006 ? array_update_84611 : array_update_84600[6];
  assign array_update_84613[7] = add_84176 == 32'h0000_0007 ? array_update_84611 : array_update_84600[7];
  assign array_update_84613[8] = add_84176 == 32'h0000_0008 ? array_update_84611 : array_update_84600[8];
  assign array_update_84613[9] = add_84176 == 32'h0000_0009 ? array_update_84611 : array_update_84600[9];
  assign array_index_84615 = array_update_72021[add_84612 > 32'h0000_0009 ? 4'h9 : add_84612[3:0]];
  assign array_index_84616 = array_update_84613[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_84620 = smul32b_32b_x_32b(array_index_84183[add_84612 > 32'h0000_0009 ? 4'h9 : add_84612[3:0]], array_index_84615[add_84584 > 32'h0000_0009 ? 4'h9 : add_84584[3:0]]);
  assign add_84622 = array_index_84616[add_84584 > 32'h0000_0009 ? 4'h9 : add_84584[3:0]] + smul_84620;
  assign array_update_84624[0] = add_84584 == 32'h0000_0000 ? add_84622 : array_index_84616[0];
  assign array_update_84624[1] = add_84584 == 32'h0000_0001 ? add_84622 : array_index_84616[1];
  assign array_update_84624[2] = add_84584 == 32'h0000_0002 ? add_84622 : array_index_84616[2];
  assign array_update_84624[3] = add_84584 == 32'h0000_0003 ? add_84622 : array_index_84616[3];
  assign array_update_84624[4] = add_84584 == 32'h0000_0004 ? add_84622 : array_index_84616[4];
  assign array_update_84624[5] = add_84584 == 32'h0000_0005 ? add_84622 : array_index_84616[5];
  assign array_update_84624[6] = add_84584 == 32'h0000_0006 ? add_84622 : array_index_84616[6];
  assign array_update_84624[7] = add_84584 == 32'h0000_0007 ? add_84622 : array_index_84616[7];
  assign array_update_84624[8] = add_84584 == 32'h0000_0008 ? add_84622 : array_index_84616[8];
  assign array_update_84624[9] = add_84584 == 32'h0000_0009 ? add_84622 : array_index_84616[9];
  assign add_84625 = add_84612 + 32'h0000_0001;
  assign array_update_84626[0] = add_84176 == 32'h0000_0000 ? array_update_84624 : array_update_84613[0];
  assign array_update_84626[1] = add_84176 == 32'h0000_0001 ? array_update_84624 : array_update_84613[1];
  assign array_update_84626[2] = add_84176 == 32'h0000_0002 ? array_update_84624 : array_update_84613[2];
  assign array_update_84626[3] = add_84176 == 32'h0000_0003 ? array_update_84624 : array_update_84613[3];
  assign array_update_84626[4] = add_84176 == 32'h0000_0004 ? array_update_84624 : array_update_84613[4];
  assign array_update_84626[5] = add_84176 == 32'h0000_0005 ? array_update_84624 : array_update_84613[5];
  assign array_update_84626[6] = add_84176 == 32'h0000_0006 ? array_update_84624 : array_update_84613[6];
  assign array_update_84626[7] = add_84176 == 32'h0000_0007 ? array_update_84624 : array_update_84613[7];
  assign array_update_84626[8] = add_84176 == 32'h0000_0008 ? array_update_84624 : array_update_84613[8];
  assign array_update_84626[9] = add_84176 == 32'h0000_0009 ? array_update_84624 : array_update_84613[9];
  assign array_index_84628 = array_update_72021[add_84625 > 32'h0000_0009 ? 4'h9 : add_84625[3:0]];
  assign array_index_84629 = array_update_84626[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_84633 = smul32b_32b_x_32b(array_index_84183[add_84625 > 32'h0000_0009 ? 4'h9 : add_84625[3:0]], array_index_84628[add_84584 > 32'h0000_0009 ? 4'h9 : add_84584[3:0]]);
  assign add_84635 = array_index_84629[add_84584 > 32'h0000_0009 ? 4'h9 : add_84584[3:0]] + smul_84633;
  assign array_update_84637[0] = add_84584 == 32'h0000_0000 ? add_84635 : array_index_84629[0];
  assign array_update_84637[1] = add_84584 == 32'h0000_0001 ? add_84635 : array_index_84629[1];
  assign array_update_84637[2] = add_84584 == 32'h0000_0002 ? add_84635 : array_index_84629[2];
  assign array_update_84637[3] = add_84584 == 32'h0000_0003 ? add_84635 : array_index_84629[3];
  assign array_update_84637[4] = add_84584 == 32'h0000_0004 ? add_84635 : array_index_84629[4];
  assign array_update_84637[5] = add_84584 == 32'h0000_0005 ? add_84635 : array_index_84629[5];
  assign array_update_84637[6] = add_84584 == 32'h0000_0006 ? add_84635 : array_index_84629[6];
  assign array_update_84637[7] = add_84584 == 32'h0000_0007 ? add_84635 : array_index_84629[7];
  assign array_update_84637[8] = add_84584 == 32'h0000_0008 ? add_84635 : array_index_84629[8];
  assign array_update_84637[9] = add_84584 == 32'h0000_0009 ? add_84635 : array_index_84629[9];
  assign add_84638 = add_84625 + 32'h0000_0001;
  assign array_update_84639[0] = add_84176 == 32'h0000_0000 ? array_update_84637 : array_update_84626[0];
  assign array_update_84639[1] = add_84176 == 32'h0000_0001 ? array_update_84637 : array_update_84626[1];
  assign array_update_84639[2] = add_84176 == 32'h0000_0002 ? array_update_84637 : array_update_84626[2];
  assign array_update_84639[3] = add_84176 == 32'h0000_0003 ? array_update_84637 : array_update_84626[3];
  assign array_update_84639[4] = add_84176 == 32'h0000_0004 ? array_update_84637 : array_update_84626[4];
  assign array_update_84639[5] = add_84176 == 32'h0000_0005 ? array_update_84637 : array_update_84626[5];
  assign array_update_84639[6] = add_84176 == 32'h0000_0006 ? array_update_84637 : array_update_84626[6];
  assign array_update_84639[7] = add_84176 == 32'h0000_0007 ? array_update_84637 : array_update_84626[7];
  assign array_update_84639[8] = add_84176 == 32'h0000_0008 ? array_update_84637 : array_update_84626[8];
  assign array_update_84639[9] = add_84176 == 32'h0000_0009 ? array_update_84637 : array_update_84626[9];
  assign array_index_84641 = array_update_72021[add_84638 > 32'h0000_0009 ? 4'h9 : add_84638[3:0]];
  assign array_index_84642 = array_update_84639[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_84646 = smul32b_32b_x_32b(array_index_84183[add_84638 > 32'h0000_0009 ? 4'h9 : add_84638[3:0]], array_index_84641[add_84584 > 32'h0000_0009 ? 4'h9 : add_84584[3:0]]);
  assign add_84648 = array_index_84642[add_84584 > 32'h0000_0009 ? 4'h9 : add_84584[3:0]] + smul_84646;
  assign array_update_84650[0] = add_84584 == 32'h0000_0000 ? add_84648 : array_index_84642[0];
  assign array_update_84650[1] = add_84584 == 32'h0000_0001 ? add_84648 : array_index_84642[1];
  assign array_update_84650[2] = add_84584 == 32'h0000_0002 ? add_84648 : array_index_84642[2];
  assign array_update_84650[3] = add_84584 == 32'h0000_0003 ? add_84648 : array_index_84642[3];
  assign array_update_84650[4] = add_84584 == 32'h0000_0004 ? add_84648 : array_index_84642[4];
  assign array_update_84650[5] = add_84584 == 32'h0000_0005 ? add_84648 : array_index_84642[5];
  assign array_update_84650[6] = add_84584 == 32'h0000_0006 ? add_84648 : array_index_84642[6];
  assign array_update_84650[7] = add_84584 == 32'h0000_0007 ? add_84648 : array_index_84642[7];
  assign array_update_84650[8] = add_84584 == 32'h0000_0008 ? add_84648 : array_index_84642[8];
  assign array_update_84650[9] = add_84584 == 32'h0000_0009 ? add_84648 : array_index_84642[9];
  assign add_84651 = add_84638 + 32'h0000_0001;
  assign array_update_84652[0] = add_84176 == 32'h0000_0000 ? array_update_84650 : array_update_84639[0];
  assign array_update_84652[1] = add_84176 == 32'h0000_0001 ? array_update_84650 : array_update_84639[1];
  assign array_update_84652[2] = add_84176 == 32'h0000_0002 ? array_update_84650 : array_update_84639[2];
  assign array_update_84652[3] = add_84176 == 32'h0000_0003 ? array_update_84650 : array_update_84639[3];
  assign array_update_84652[4] = add_84176 == 32'h0000_0004 ? array_update_84650 : array_update_84639[4];
  assign array_update_84652[5] = add_84176 == 32'h0000_0005 ? array_update_84650 : array_update_84639[5];
  assign array_update_84652[6] = add_84176 == 32'h0000_0006 ? array_update_84650 : array_update_84639[6];
  assign array_update_84652[7] = add_84176 == 32'h0000_0007 ? array_update_84650 : array_update_84639[7];
  assign array_update_84652[8] = add_84176 == 32'h0000_0008 ? array_update_84650 : array_update_84639[8];
  assign array_update_84652[9] = add_84176 == 32'h0000_0009 ? array_update_84650 : array_update_84639[9];
  assign array_index_84654 = array_update_72021[add_84651 > 32'h0000_0009 ? 4'h9 : add_84651[3:0]];
  assign array_index_84655 = array_update_84652[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_84659 = smul32b_32b_x_32b(array_index_84183[add_84651 > 32'h0000_0009 ? 4'h9 : add_84651[3:0]], array_index_84654[add_84584 > 32'h0000_0009 ? 4'h9 : add_84584[3:0]]);
  assign add_84661 = array_index_84655[add_84584 > 32'h0000_0009 ? 4'h9 : add_84584[3:0]] + smul_84659;
  assign array_update_84663[0] = add_84584 == 32'h0000_0000 ? add_84661 : array_index_84655[0];
  assign array_update_84663[1] = add_84584 == 32'h0000_0001 ? add_84661 : array_index_84655[1];
  assign array_update_84663[2] = add_84584 == 32'h0000_0002 ? add_84661 : array_index_84655[2];
  assign array_update_84663[3] = add_84584 == 32'h0000_0003 ? add_84661 : array_index_84655[3];
  assign array_update_84663[4] = add_84584 == 32'h0000_0004 ? add_84661 : array_index_84655[4];
  assign array_update_84663[5] = add_84584 == 32'h0000_0005 ? add_84661 : array_index_84655[5];
  assign array_update_84663[6] = add_84584 == 32'h0000_0006 ? add_84661 : array_index_84655[6];
  assign array_update_84663[7] = add_84584 == 32'h0000_0007 ? add_84661 : array_index_84655[7];
  assign array_update_84663[8] = add_84584 == 32'h0000_0008 ? add_84661 : array_index_84655[8];
  assign array_update_84663[9] = add_84584 == 32'h0000_0009 ? add_84661 : array_index_84655[9];
  assign add_84664 = add_84651 + 32'h0000_0001;
  assign array_update_84665[0] = add_84176 == 32'h0000_0000 ? array_update_84663 : array_update_84652[0];
  assign array_update_84665[1] = add_84176 == 32'h0000_0001 ? array_update_84663 : array_update_84652[1];
  assign array_update_84665[2] = add_84176 == 32'h0000_0002 ? array_update_84663 : array_update_84652[2];
  assign array_update_84665[3] = add_84176 == 32'h0000_0003 ? array_update_84663 : array_update_84652[3];
  assign array_update_84665[4] = add_84176 == 32'h0000_0004 ? array_update_84663 : array_update_84652[4];
  assign array_update_84665[5] = add_84176 == 32'h0000_0005 ? array_update_84663 : array_update_84652[5];
  assign array_update_84665[6] = add_84176 == 32'h0000_0006 ? array_update_84663 : array_update_84652[6];
  assign array_update_84665[7] = add_84176 == 32'h0000_0007 ? array_update_84663 : array_update_84652[7];
  assign array_update_84665[8] = add_84176 == 32'h0000_0008 ? array_update_84663 : array_update_84652[8];
  assign array_update_84665[9] = add_84176 == 32'h0000_0009 ? array_update_84663 : array_update_84652[9];
  assign array_index_84667 = array_update_72021[add_84664 > 32'h0000_0009 ? 4'h9 : add_84664[3:0]];
  assign array_index_84668 = array_update_84665[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_84672 = smul32b_32b_x_32b(array_index_84183[add_84664 > 32'h0000_0009 ? 4'h9 : add_84664[3:0]], array_index_84667[add_84584 > 32'h0000_0009 ? 4'h9 : add_84584[3:0]]);
  assign add_84674 = array_index_84668[add_84584 > 32'h0000_0009 ? 4'h9 : add_84584[3:0]] + smul_84672;
  assign array_update_84676[0] = add_84584 == 32'h0000_0000 ? add_84674 : array_index_84668[0];
  assign array_update_84676[1] = add_84584 == 32'h0000_0001 ? add_84674 : array_index_84668[1];
  assign array_update_84676[2] = add_84584 == 32'h0000_0002 ? add_84674 : array_index_84668[2];
  assign array_update_84676[3] = add_84584 == 32'h0000_0003 ? add_84674 : array_index_84668[3];
  assign array_update_84676[4] = add_84584 == 32'h0000_0004 ? add_84674 : array_index_84668[4];
  assign array_update_84676[5] = add_84584 == 32'h0000_0005 ? add_84674 : array_index_84668[5];
  assign array_update_84676[6] = add_84584 == 32'h0000_0006 ? add_84674 : array_index_84668[6];
  assign array_update_84676[7] = add_84584 == 32'h0000_0007 ? add_84674 : array_index_84668[7];
  assign array_update_84676[8] = add_84584 == 32'h0000_0008 ? add_84674 : array_index_84668[8];
  assign array_update_84676[9] = add_84584 == 32'h0000_0009 ? add_84674 : array_index_84668[9];
  assign add_84677 = add_84664 + 32'h0000_0001;
  assign array_update_84678[0] = add_84176 == 32'h0000_0000 ? array_update_84676 : array_update_84665[0];
  assign array_update_84678[1] = add_84176 == 32'h0000_0001 ? array_update_84676 : array_update_84665[1];
  assign array_update_84678[2] = add_84176 == 32'h0000_0002 ? array_update_84676 : array_update_84665[2];
  assign array_update_84678[3] = add_84176 == 32'h0000_0003 ? array_update_84676 : array_update_84665[3];
  assign array_update_84678[4] = add_84176 == 32'h0000_0004 ? array_update_84676 : array_update_84665[4];
  assign array_update_84678[5] = add_84176 == 32'h0000_0005 ? array_update_84676 : array_update_84665[5];
  assign array_update_84678[6] = add_84176 == 32'h0000_0006 ? array_update_84676 : array_update_84665[6];
  assign array_update_84678[7] = add_84176 == 32'h0000_0007 ? array_update_84676 : array_update_84665[7];
  assign array_update_84678[8] = add_84176 == 32'h0000_0008 ? array_update_84676 : array_update_84665[8];
  assign array_update_84678[9] = add_84176 == 32'h0000_0009 ? array_update_84676 : array_update_84665[9];
  assign array_index_84680 = array_update_72021[add_84677 > 32'h0000_0009 ? 4'h9 : add_84677[3:0]];
  assign array_index_84681 = array_update_84678[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_84685 = smul32b_32b_x_32b(array_index_84183[add_84677 > 32'h0000_0009 ? 4'h9 : add_84677[3:0]], array_index_84680[add_84584 > 32'h0000_0009 ? 4'h9 : add_84584[3:0]]);
  assign add_84687 = array_index_84681[add_84584 > 32'h0000_0009 ? 4'h9 : add_84584[3:0]] + smul_84685;
  assign array_update_84689[0] = add_84584 == 32'h0000_0000 ? add_84687 : array_index_84681[0];
  assign array_update_84689[1] = add_84584 == 32'h0000_0001 ? add_84687 : array_index_84681[1];
  assign array_update_84689[2] = add_84584 == 32'h0000_0002 ? add_84687 : array_index_84681[2];
  assign array_update_84689[3] = add_84584 == 32'h0000_0003 ? add_84687 : array_index_84681[3];
  assign array_update_84689[4] = add_84584 == 32'h0000_0004 ? add_84687 : array_index_84681[4];
  assign array_update_84689[5] = add_84584 == 32'h0000_0005 ? add_84687 : array_index_84681[5];
  assign array_update_84689[6] = add_84584 == 32'h0000_0006 ? add_84687 : array_index_84681[6];
  assign array_update_84689[7] = add_84584 == 32'h0000_0007 ? add_84687 : array_index_84681[7];
  assign array_update_84689[8] = add_84584 == 32'h0000_0008 ? add_84687 : array_index_84681[8];
  assign array_update_84689[9] = add_84584 == 32'h0000_0009 ? add_84687 : array_index_84681[9];
  assign add_84690 = add_84677 + 32'h0000_0001;
  assign array_update_84691[0] = add_84176 == 32'h0000_0000 ? array_update_84689 : array_update_84678[0];
  assign array_update_84691[1] = add_84176 == 32'h0000_0001 ? array_update_84689 : array_update_84678[1];
  assign array_update_84691[2] = add_84176 == 32'h0000_0002 ? array_update_84689 : array_update_84678[2];
  assign array_update_84691[3] = add_84176 == 32'h0000_0003 ? array_update_84689 : array_update_84678[3];
  assign array_update_84691[4] = add_84176 == 32'h0000_0004 ? array_update_84689 : array_update_84678[4];
  assign array_update_84691[5] = add_84176 == 32'h0000_0005 ? array_update_84689 : array_update_84678[5];
  assign array_update_84691[6] = add_84176 == 32'h0000_0006 ? array_update_84689 : array_update_84678[6];
  assign array_update_84691[7] = add_84176 == 32'h0000_0007 ? array_update_84689 : array_update_84678[7];
  assign array_update_84691[8] = add_84176 == 32'h0000_0008 ? array_update_84689 : array_update_84678[8];
  assign array_update_84691[9] = add_84176 == 32'h0000_0009 ? array_update_84689 : array_update_84678[9];
  assign array_index_84693 = array_update_72021[add_84690 > 32'h0000_0009 ? 4'h9 : add_84690[3:0]];
  assign array_index_84694 = array_update_84691[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_84698 = smul32b_32b_x_32b(array_index_84183[add_84690 > 32'h0000_0009 ? 4'h9 : add_84690[3:0]], array_index_84693[add_84584 > 32'h0000_0009 ? 4'h9 : add_84584[3:0]]);
  assign add_84700 = array_index_84694[add_84584 > 32'h0000_0009 ? 4'h9 : add_84584[3:0]] + smul_84698;
  assign array_update_84702[0] = add_84584 == 32'h0000_0000 ? add_84700 : array_index_84694[0];
  assign array_update_84702[1] = add_84584 == 32'h0000_0001 ? add_84700 : array_index_84694[1];
  assign array_update_84702[2] = add_84584 == 32'h0000_0002 ? add_84700 : array_index_84694[2];
  assign array_update_84702[3] = add_84584 == 32'h0000_0003 ? add_84700 : array_index_84694[3];
  assign array_update_84702[4] = add_84584 == 32'h0000_0004 ? add_84700 : array_index_84694[4];
  assign array_update_84702[5] = add_84584 == 32'h0000_0005 ? add_84700 : array_index_84694[5];
  assign array_update_84702[6] = add_84584 == 32'h0000_0006 ? add_84700 : array_index_84694[6];
  assign array_update_84702[7] = add_84584 == 32'h0000_0007 ? add_84700 : array_index_84694[7];
  assign array_update_84702[8] = add_84584 == 32'h0000_0008 ? add_84700 : array_index_84694[8];
  assign array_update_84702[9] = add_84584 == 32'h0000_0009 ? add_84700 : array_index_84694[9];
  assign add_84703 = add_84690 + 32'h0000_0001;
  assign array_update_84704[0] = add_84176 == 32'h0000_0000 ? array_update_84702 : array_update_84691[0];
  assign array_update_84704[1] = add_84176 == 32'h0000_0001 ? array_update_84702 : array_update_84691[1];
  assign array_update_84704[2] = add_84176 == 32'h0000_0002 ? array_update_84702 : array_update_84691[2];
  assign array_update_84704[3] = add_84176 == 32'h0000_0003 ? array_update_84702 : array_update_84691[3];
  assign array_update_84704[4] = add_84176 == 32'h0000_0004 ? array_update_84702 : array_update_84691[4];
  assign array_update_84704[5] = add_84176 == 32'h0000_0005 ? array_update_84702 : array_update_84691[5];
  assign array_update_84704[6] = add_84176 == 32'h0000_0006 ? array_update_84702 : array_update_84691[6];
  assign array_update_84704[7] = add_84176 == 32'h0000_0007 ? array_update_84702 : array_update_84691[7];
  assign array_update_84704[8] = add_84176 == 32'h0000_0008 ? array_update_84702 : array_update_84691[8];
  assign array_update_84704[9] = add_84176 == 32'h0000_0009 ? array_update_84702 : array_update_84691[9];
  assign array_index_84706 = array_update_72021[add_84703 > 32'h0000_0009 ? 4'h9 : add_84703[3:0]];
  assign array_index_84707 = array_update_84704[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_84711 = smul32b_32b_x_32b(array_index_84183[add_84703 > 32'h0000_0009 ? 4'h9 : add_84703[3:0]], array_index_84706[add_84584 > 32'h0000_0009 ? 4'h9 : add_84584[3:0]]);
  assign add_84713 = array_index_84707[add_84584 > 32'h0000_0009 ? 4'h9 : add_84584[3:0]] + smul_84711;
  assign array_update_84714[0] = add_84584 == 32'h0000_0000 ? add_84713 : array_index_84707[0];
  assign array_update_84714[1] = add_84584 == 32'h0000_0001 ? add_84713 : array_index_84707[1];
  assign array_update_84714[2] = add_84584 == 32'h0000_0002 ? add_84713 : array_index_84707[2];
  assign array_update_84714[3] = add_84584 == 32'h0000_0003 ? add_84713 : array_index_84707[3];
  assign array_update_84714[4] = add_84584 == 32'h0000_0004 ? add_84713 : array_index_84707[4];
  assign array_update_84714[5] = add_84584 == 32'h0000_0005 ? add_84713 : array_index_84707[5];
  assign array_update_84714[6] = add_84584 == 32'h0000_0006 ? add_84713 : array_index_84707[6];
  assign array_update_84714[7] = add_84584 == 32'h0000_0007 ? add_84713 : array_index_84707[7];
  assign array_update_84714[8] = add_84584 == 32'h0000_0008 ? add_84713 : array_index_84707[8];
  assign array_update_84714[9] = add_84584 == 32'h0000_0009 ? add_84713 : array_index_84707[9];
  assign array_update_84715[0] = add_84176 == 32'h0000_0000 ? array_update_84714 : array_update_84704[0];
  assign array_update_84715[1] = add_84176 == 32'h0000_0001 ? array_update_84714 : array_update_84704[1];
  assign array_update_84715[2] = add_84176 == 32'h0000_0002 ? array_update_84714 : array_update_84704[2];
  assign array_update_84715[3] = add_84176 == 32'h0000_0003 ? array_update_84714 : array_update_84704[3];
  assign array_update_84715[4] = add_84176 == 32'h0000_0004 ? array_update_84714 : array_update_84704[4];
  assign array_update_84715[5] = add_84176 == 32'h0000_0005 ? array_update_84714 : array_update_84704[5];
  assign array_update_84715[6] = add_84176 == 32'h0000_0006 ? array_update_84714 : array_update_84704[6];
  assign array_update_84715[7] = add_84176 == 32'h0000_0007 ? array_update_84714 : array_update_84704[7];
  assign array_update_84715[8] = add_84176 == 32'h0000_0008 ? array_update_84714 : array_update_84704[8];
  assign array_update_84715[9] = add_84176 == 32'h0000_0009 ? array_update_84714 : array_update_84704[9];
  assign array_index_84717 = array_update_84715[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign add_84719 = add_84584 + 32'h0000_0001;
  assign array_update_84720[0] = add_84719 == 32'h0000_0000 ? 32'h0000_0000 : array_index_84717[0];
  assign array_update_84720[1] = add_84719 == 32'h0000_0001 ? 32'h0000_0000 : array_index_84717[1];
  assign array_update_84720[2] = add_84719 == 32'h0000_0002 ? 32'h0000_0000 : array_index_84717[2];
  assign array_update_84720[3] = add_84719 == 32'h0000_0003 ? 32'h0000_0000 : array_index_84717[3];
  assign array_update_84720[4] = add_84719 == 32'h0000_0004 ? 32'h0000_0000 : array_index_84717[4];
  assign array_update_84720[5] = add_84719 == 32'h0000_0005 ? 32'h0000_0000 : array_index_84717[5];
  assign array_update_84720[6] = add_84719 == 32'h0000_0006 ? 32'h0000_0000 : array_index_84717[6];
  assign array_update_84720[7] = add_84719 == 32'h0000_0007 ? 32'h0000_0000 : array_index_84717[7];
  assign array_update_84720[8] = add_84719 == 32'h0000_0008 ? 32'h0000_0000 : array_index_84717[8];
  assign array_update_84720[9] = add_84719 == 32'h0000_0009 ? 32'h0000_0000 : array_index_84717[9];
  assign literal_84721 = 32'h0000_0000;
  assign array_update_84722[0] = add_84176 == 32'h0000_0000 ? array_update_84720 : array_update_84715[0];
  assign array_update_84722[1] = add_84176 == 32'h0000_0001 ? array_update_84720 : array_update_84715[1];
  assign array_update_84722[2] = add_84176 == 32'h0000_0002 ? array_update_84720 : array_update_84715[2];
  assign array_update_84722[3] = add_84176 == 32'h0000_0003 ? array_update_84720 : array_update_84715[3];
  assign array_update_84722[4] = add_84176 == 32'h0000_0004 ? array_update_84720 : array_update_84715[4];
  assign array_update_84722[5] = add_84176 == 32'h0000_0005 ? array_update_84720 : array_update_84715[5];
  assign array_update_84722[6] = add_84176 == 32'h0000_0006 ? array_update_84720 : array_update_84715[6];
  assign array_update_84722[7] = add_84176 == 32'h0000_0007 ? array_update_84720 : array_update_84715[7];
  assign array_update_84722[8] = add_84176 == 32'h0000_0008 ? array_update_84720 : array_update_84715[8];
  assign array_update_84722[9] = add_84176 == 32'h0000_0009 ? array_update_84720 : array_update_84715[9];
  assign array_index_84724 = array_update_72021[literal_84721 > 32'h0000_0009 ? 4'h9 : literal_84721[3:0]];
  assign array_index_84725 = array_update_84722[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_84729 = smul32b_32b_x_32b(array_index_84183[literal_84721 > 32'h0000_0009 ? 4'h9 : literal_84721[3:0]], array_index_84724[add_84719 > 32'h0000_0009 ? 4'h9 : add_84719[3:0]]);
  assign add_84731 = array_index_84725[add_84719 > 32'h0000_0009 ? 4'h9 : add_84719[3:0]] + smul_84729;
  assign array_update_84733[0] = add_84719 == 32'h0000_0000 ? add_84731 : array_index_84725[0];
  assign array_update_84733[1] = add_84719 == 32'h0000_0001 ? add_84731 : array_index_84725[1];
  assign array_update_84733[2] = add_84719 == 32'h0000_0002 ? add_84731 : array_index_84725[2];
  assign array_update_84733[3] = add_84719 == 32'h0000_0003 ? add_84731 : array_index_84725[3];
  assign array_update_84733[4] = add_84719 == 32'h0000_0004 ? add_84731 : array_index_84725[4];
  assign array_update_84733[5] = add_84719 == 32'h0000_0005 ? add_84731 : array_index_84725[5];
  assign array_update_84733[6] = add_84719 == 32'h0000_0006 ? add_84731 : array_index_84725[6];
  assign array_update_84733[7] = add_84719 == 32'h0000_0007 ? add_84731 : array_index_84725[7];
  assign array_update_84733[8] = add_84719 == 32'h0000_0008 ? add_84731 : array_index_84725[8];
  assign array_update_84733[9] = add_84719 == 32'h0000_0009 ? add_84731 : array_index_84725[9];
  assign add_84734 = literal_84721 + 32'h0000_0001;
  assign array_update_84735[0] = add_84176 == 32'h0000_0000 ? array_update_84733 : array_update_84722[0];
  assign array_update_84735[1] = add_84176 == 32'h0000_0001 ? array_update_84733 : array_update_84722[1];
  assign array_update_84735[2] = add_84176 == 32'h0000_0002 ? array_update_84733 : array_update_84722[2];
  assign array_update_84735[3] = add_84176 == 32'h0000_0003 ? array_update_84733 : array_update_84722[3];
  assign array_update_84735[4] = add_84176 == 32'h0000_0004 ? array_update_84733 : array_update_84722[4];
  assign array_update_84735[5] = add_84176 == 32'h0000_0005 ? array_update_84733 : array_update_84722[5];
  assign array_update_84735[6] = add_84176 == 32'h0000_0006 ? array_update_84733 : array_update_84722[6];
  assign array_update_84735[7] = add_84176 == 32'h0000_0007 ? array_update_84733 : array_update_84722[7];
  assign array_update_84735[8] = add_84176 == 32'h0000_0008 ? array_update_84733 : array_update_84722[8];
  assign array_update_84735[9] = add_84176 == 32'h0000_0009 ? array_update_84733 : array_update_84722[9];
  assign array_index_84737 = array_update_72021[add_84734 > 32'h0000_0009 ? 4'h9 : add_84734[3:0]];
  assign array_index_84738 = array_update_84735[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_84742 = smul32b_32b_x_32b(array_index_84183[add_84734 > 32'h0000_0009 ? 4'h9 : add_84734[3:0]], array_index_84737[add_84719 > 32'h0000_0009 ? 4'h9 : add_84719[3:0]]);
  assign add_84744 = array_index_84738[add_84719 > 32'h0000_0009 ? 4'h9 : add_84719[3:0]] + smul_84742;
  assign array_update_84746[0] = add_84719 == 32'h0000_0000 ? add_84744 : array_index_84738[0];
  assign array_update_84746[1] = add_84719 == 32'h0000_0001 ? add_84744 : array_index_84738[1];
  assign array_update_84746[2] = add_84719 == 32'h0000_0002 ? add_84744 : array_index_84738[2];
  assign array_update_84746[3] = add_84719 == 32'h0000_0003 ? add_84744 : array_index_84738[3];
  assign array_update_84746[4] = add_84719 == 32'h0000_0004 ? add_84744 : array_index_84738[4];
  assign array_update_84746[5] = add_84719 == 32'h0000_0005 ? add_84744 : array_index_84738[5];
  assign array_update_84746[6] = add_84719 == 32'h0000_0006 ? add_84744 : array_index_84738[6];
  assign array_update_84746[7] = add_84719 == 32'h0000_0007 ? add_84744 : array_index_84738[7];
  assign array_update_84746[8] = add_84719 == 32'h0000_0008 ? add_84744 : array_index_84738[8];
  assign array_update_84746[9] = add_84719 == 32'h0000_0009 ? add_84744 : array_index_84738[9];
  assign add_84747 = add_84734 + 32'h0000_0001;
  assign array_update_84748[0] = add_84176 == 32'h0000_0000 ? array_update_84746 : array_update_84735[0];
  assign array_update_84748[1] = add_84176 == 32'h0000_0001 ? array_update_84746 : array_update_84735[1];
  assign array_update_84748[2] = add_84176 == 32'h0000_0002 ? array_update_84746 : array_update_84735[2];
  assign array_update_84748[3] = add_84176 == 32'h0000_0003 ? array_update_84746 : array_update_84735[3];
  assign array_update_84748[4] = add_84176 == 32'h0000_0004 ? array_update_84746 : array_update_84735[4];
  assign array_update_84748[5] = add_84176 == 32'h0000_0005 ? array_update_84746 : array_update_84735[5];
  assign array_update_84748[6] = add_84176 == 32'h0000_0006 ? array_update_84746 : array_update_84735[6];
  assign array_update_84748[7] = add_84176 == 32'h0000_0007 ? array_update_84746 : array_update_84735[7];
  assign array_update_84748[8] = add_84176 == 32'h0000_0008 ? array_update_84746 : array_update_84735[8];
  assign array_update_84748[9] = add_84176 == 32'h0000_0009 ? array_update_84746 : array_update_84735[9];
  assign array_index_84750 = array_update_72021[add_84747 > 32'h0000_0009 ? 4'h9 : add_84747[3:0]];
  assign array_index_84751 = array_update_84748[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_84755 = smul32b_32b_x_32b(array_index_84183[add_84747 > 32'h0000_0009 ? 4'h9 : add_84747[3:0]], array_index_84750[add_84719 > 32'h0000_0009 ? 4'h9 : add_84719[3:0]]);
  assign add_84757 = array_index_84751[add_84719 > 32'h0000_0009 ? 4'h9 : add_84719[3:0]] + smul_84755;
  assign array_update_84759[0] = add_84719 == 32'h0000_0000 ? add_84757 : array_index_84751[0];
  assign array_update_84759[1] = add_84719 == 32'h0000_0001 ? add_84757 : array_index_84751[1];
  assign array_update_84759[2] = add_84719 == 32'h0000_0002 ? add_84757 : array_index_84751[2];
  assign array_update_84759[3] = add_84719 == 32'h0000_0003 ? add_84757 : array_index_84751[3];
  assign array_update_84759[4] = add_84719 == 32'h0000_0004 ? add_84757 : array_index_84751[4];
  assign array_update_84759[5] = add_84719 == 32'h0000_0005 ? add_84757 : array_index_84751[5];
  assign array_update_84759[6] = add_84719 == 32'h0000_0006 ? add_84757 : array_index_84751[6];
  assign array_update_84759[7] = add_84719 == 32'h0000_0007 ? add_84757 : array_index_84751[7];
  assign array_update_84759[8] = add_84719 == 32'h0000_0008 ? add_84757 : array_index_84751[8];
  assign array_update_84759[9] = add_84719 == 32'h0000_0009 ? add_84757 : array_index_84751[9];
  assign add_84760 = add_84747 + 32'h0000_0001;
  assign array_update_84761[0] = add_84176 == 32'h0000_0000 ? array_update_84759 : array_update_84748[0];
  assign array_update_84761[1] = add_84176 == 32'h0000_0001 ? array_update_84759 : array_update_84748[1];
  assign array_update_84761[2] = add_84176 == 32'h0000_0002 ? array_update_84759 : array_update_84748[2];
  assign array_update_84761[3] = add_84176 == 32'h0000_0003 ? array_update_84759 : array_update_84748[3];
  assign array_update_84761[4] = add_84176 == 32'h0000_0004 ? array_update_84759 : array_update_84748[4];
  assign array_update_84761[5] = add_84176 == 32'h0000_0005 ? array_update_84759 : array_update_84748[5];
  assign array_update_84761[6] = add_84176 == 32'h0000_0006 ? array_update_84759 : array_update_84748[6];
  assign array_update_84761[7] = add_84176 == 32'h0000_0007 ? array_update_84759 : array_update_84748[7];
  assign array_update_84761[8] = add_84176 == 32'h0000_0008 ? array_update_84759 : array_update_84748[8];
  assign array_update_84761[9] = add_84176 == 32'h0000_0009 ? array_update_84759 : array_update_84748[9];
  assign array_index_84763 = array_update_72021[add_84760 > 32'h0000_0009 ? 4'h9 : add_84760[3:0]];
  assign array_index_84764 = array_update_84761[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_84768 = smul32b_32b_x_32b(array_index_84183[add_84760 > 32'h0000_0009 ? 4'h9 : add_84760[3:0]], array_index_84763[add_84719 > 32'h0000_0009 ? 4'h9 : add_84719[3:0]]);
  assign add_84770 = array_index_84764[add_84719 > 32'h0000_0009 ? 4'h9 : add_84719[3:0]] + smul_84768;
  assign array_update_84772[0] = add_84719 == 32'h0000_0000 ? add_84770 : array_index_84764[0];
  assign array_update_84772[1] = add_84719 == 32'h0000_0001 ? add_84770 : array_index_84764[1];
  assign array_update_84772[2] = add_84719 == 32'h0000_0002 ? add_84770 : array_index_84764[2];
  assign array_update_84772[3] = add_84719 == 32'h0000_0003 ? add_84770 : array_index_84764[3];
  assign array_update_84772[4] = add_84719 == 32'h0000_0004 ? add_84770 : array_index_84764[4];
  assign array_update_84772[5] = add_84719 == 32'h0000_0005 ? add_84770 : array_index_84764[5];
  assign array_update_84772[6] = add_84719 == 32'h0000_0006 ? add_84770 : array_index_84764[6];
  assign array_update_84772[7] = add_84719 == 32'h0000_0007 ? add_84770 : array_index_84764[7];
  assign array_update_84772[8] = add_84719 == 32'h0000_0008 ? add_84770 : array_index_84764[8];
  assign array_update_84772[9] = add_84719 == 32'h0000_0009 ? add_84770 : array_index_84764[9];
  assign add_84773 = add_84760 + 32'h0000_0001;
  assign array_update_84774[0] = add_84176 == 32'h0000_0000 ? array_update_84772 : array_update_84761[0];
  assign array_update_84774[1] = add_84176 == 32'h0000_0001 ? array_update_84772 : array_update_84761[1];
  assign array_update_84774[2] = add_84176 == 32'h0000_0002 ? array_update_84772 : array_update_84761[2];
  assign array_update_84774[3] = add_84176 == 32'h0000_0003 ? array_update_84772 : array_update_84761[3];
  assign array_update_84774[4] = add_84176 == 32'h0000_0004 ? array_update_84772 : array_update_84761[4];
  assign array_update_84774[5] = add_84176 == 32'h0000_0005 ? array_update_84772 : array_update_84761[5];
  assign array_update_84774[6] = add_84176 == 32'h0000_0006 ? array_update_84772 : array_update_84761[6];
  assign array_update_84774[7] = add_84176 == 32'h0000_0007 ? array_update_84772 : array_update_84761[7];
  assign array_update_84774[8] = add_84176 == 32'h0000_0008 ? array_update_84772 : array_update_84761[8];
  assign array_update_84774[9] = add_84176 == 32'h0000_0009 ? array_update_84772 : array_update_84761[9];
  assign array_index_84776 = array_update_72021[add_84773 > 32'h0000_0009 ? 4'h9 : add_84773[3:0]];
  assign array_index_84777 = array_update_84774[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_84781 = smul32b_32b_x_32b(array_index_84183[add_84773 > 32'h0000_0009 ? 4'h9 : add_84773[3:0]], array_index_84776[add_84719 > 32'h0000_0009 ? 4'h9 : add_84719[3:0]]);
  assign add_84783 = array_index_84777[add_84719 > 32'h0000_0009 ? 4'h9 : add_84719[3:0]] + smul_84781;
  assign array_update_84785[0] = add_84719 == 32'h0000_0000 ? add_84783 : array_index_84777[0];
  assign array_update_84785[1] = add_84719 == 32'h0000_0001 ? add_84783 : array_index_84777[1];
  assign array_update_84785[2] = add_84719 == 32'h0000_0002 ? add_84783 : array_index_84777[2];
  assign array_update_84785[3] = add_84719 == 32'h0000_0003 ? add_84783 : array_index_84777[3];
  assign array_update_84785[4] = add_84719 == 32'h0000_0004 ? add_84783 : array_index_84777[4];
  assign array_update_84785[5] = add_84719 == 32'h0000_0005 ? add_84783 : array_index_84777[5];
  assign array_update_84785[6] = add_84719 == 32'h0000_0006 ? add_84783 : array_index_84777[6];
  assign array_update_84785[7] = add_84719 == 32'h0000_0007 ? add_84783 : array_index_84777[7];
  assign array_update_84785[8] = add_84719 == 32'h0000_0008 ? add_84783 : array_index_84777[8];
  assign array_update_84785[9] = add_84719 == 32'h0000_0009 ? add_84783 : array_index_84777[9];
  assign add_84786 = add_84773 + 32'h0000_0001;
  assign array_update_84787[0] = add_84176 == 32'h0000_0000 ? array_update_84785 : array_update_84774[0];
  assign array_update_84787[1] = add_84176 == 32'h0000_0001 ? array_update_84785 : array_update_84774[1];
  assign array_update_84787[2] = add_84176 == 32'h0000_0002 ? array_update_84785 : array_update_84774[2];
  assign array_update_84787[3] = add_84176 == 32'h0000_0003 ? array_update_84785 : array_update_84774[3];
  assign array_update_84787[4] = add_84176 == 32'h0000_0004 ? array_update_84785 : array_update_84774[4];
  assign array_update_84787[5] = add_84176 == 32'h0000_0005 ? array_update_84785 : array_update_84774[5];
  assign array_update_84787[6] = add_84176 == 32'h0000_0006 ? array_update_84785 : array_update_84774[6];
  assign array_update_84787[7] = add_84176 == 32'h0000_0007 ? array_update_84785 : array_update_84774[7];
  assign array_update_84787[8] = add_84176 == 32'h0000_0008 ? array_update_84785 : array_update_84774[8];
  assign array_update_84787[9] = add_84176 == 32'h0000_0009 ? array_update_84785 : array_update_84774[9];
  assign array_index_84789 = array_update_72021[add_84786 > 32'h0000_0009 ? 4'h9 : add_84786[3:0]];
  assign array_index_84790 = array_update_84787[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_84794 = smul32b_32b_x_32b(array_index_84183[add_84786 > 32'h0000_0009 ? 4'h9 : add_84786[3:0]], array_index_84789[add_84719 > 32'h0000_0009 ? 4'h9 : add_84719[3:0]]);
  assign add_84796 = array_index_84790[add_84719 > 32'h0000_0009 ? 4'h9 : add_84719[3:0]] + smul_84794;
  assign array_update_84798[0] = add_84719 == 32'h0000_0000 ? add_84796 : array_index_84790[0];
  assign array_update_84798[1] = add_84719 == 32'h0000_0001 ? add_84796 : array_index_84790[1];
  assign array_update_84798[2] = add_84719 == 32'h0000_0002 ? add_84796 : array_index_84790[2];
  assign array_update_84798[3] = add_84719 == 32'h0000_0003 ? add_84796 : array_index_84790[3];
  assign array_update_84798[4] = add_84719 == 32'h0000_0004 ? add_84796 : array_index_84790[4];
  assign array_update_84798[5] = add_84719 == 32'h0000_0005 ? add_84796 : array_index_84790[5];
  assign array_update_84798[6] = add_84719 == 32'h0000_0006 ? add_84796 : array_index_84790[6];
  assign array_update_84798[7] = add_84719 == 32'h0000_0007 ? add_84796 : array_index_84790[7];
  assign array_update_84798[8] = add_84719 == 32'h0000_0008 ? add_84796 : array_index_84790[8];
  assign array_update_84798[9] = add_84719 == 32'h0000_0009 ? add_84796 : array_index_84790[9];
  assign add_84799 = add_84786 + 32'h0000_0001;
  assign array_update_84800[0] = add_84176 == 32'h0000_0000 ? array_update_84798 : array_update_84787[0];
  assign array_update_84800[1] = add_84176 == 32'h0000_0001 ? array_update_84798 : array_update_84787[1];
  assign array_update_84800[2] = add_84176 == 32'h0000_0002 ? array_update_84798 : array_update_84787[2];
  assign array_update_84800[3] = add_84176 == 32'h0000_0003 ? array_update_84798 : array_update_84787[3];
  assign array_update_84800[4] = add_84176 == 32'h0000_0004 ? array_update_84798 : array_update_84787[4];
  assign array_update_84800[5] = add_84176 == 32'h0000_0005 ? array_update_84798 : array_update_84787[5];
  assign array_update_84800[6] = add_84176 == 32'h0000_0006 ? array_update_84798 : array_update_84787[6];
  assign array_update_84800[7] = add_84176 == 32'h0000_0007 ? array_update_84798 : array_update_84787[7];
  assign array_update_84800[8] = add_84176 == 32'h0000_0008 ? array_update_84798 : array_update_84787[8];
  assign array_update_84800[9] = add_84176 == 32'h0000_0009 ? array_update_84798 : array_update_84787[9];
  assign array_index_84802 = array_update_72021[add_84799 > 32'h0000_0009 ? 4'h9 : add_84799[3:0]];
  assign array_index_84803 = array_update_84800[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_84807 = smul32b_32b_x_32b(array_index_84183[add_84799 > 32'h0000_0009 ? 4'h9 : add_84799[3:0]], array_index_84802[add_84719 > 32'h0000_0009 ? 4'h9 : add_84719[3:0]]);
  assign add_84809 = array_index_84803[add_84719 > 32'h0000_0009 ? 4'h9 : add_84719[3:0]] + smul_84807;
  assign array_update_84811[0] = add_84719 == 32'h0000_0000 ? add_84809 : array_index_84803[0];
  assign array_update_84811[1] = add_84719 == 32'h0000_0001 ? add_84809 : array_index_84803[1];
  assign array_update_84811[2] = add_84719 == 32'h0000_0002 ? add_84809 : array_index_84803[2];
  assign array_update_84811[3] = add_84719 == 32'h0000_0003 ? add_84809 : array_index_84803[3];
  assign array_update_84811[4] = add_84719 == 32'h0000_0004 ? add_84809 : array_index_84803[4];
  assign array_update_84811[5] = add_84719 == 32'h0000_0005 ? add_84809 : array_index_84803[5];
  assign array_update_84811[6] = add_84719 == 32'h0000_0006 ? add_84809 : array_index_84803[6];
  assign array_update_84811[7] = add_84719 == 32'h0000_0007 ? add_84809 : array_index_84803[7];
  assign array_update_84811[8] = add_84719 == 32'h0000_0008 ? add_84809 : array_index_84803[8];
  assign array_update_84811[9] = add_84719 == 32'h0000_0009 ? add_84809 : array_index_84803[9];
  assign add_84812 = add_84799 + 32'h0000_0001;
  assign array_update_84813[0] = add_84176 == 32'h0000_0000 ? array_update_84811 : array_update_84800[0];
  assign array_update_84813[1] = add_84176 == 32'h0000_0001 ? array_update_84811 : array_update_84800[1];
  assign array_update_84813[2] = add_84176 == 32'h0000_0002 ? array_update_84811 : array_update_84800[2];
  assign array_update_84813[3] = add_84176 == 32'h0000_0003 ? array_update_84811 : array_update_84800[3];
  assign array_update_84813[4] = add_84176 == 32'h0000_0004 ? array_update_84811 : array_update_84800[4];
  assign array_update_84813[5] = add_84176 == 32'h0000_0005 ? array_update_84811 : array_update_84800[5];
  assign array_update_84813[6] = add_84176 == 32'h0000_0006 ? array_update_84811 : array_update_84800[6];
  assign array_update_84813[7] = add_84176 == 32'h0000_0007 ? array_update_84811 : array_update_84800[7];
  assign array_update_84813[8] = add_84176 == 32'h0000_0008 ? array_update_84811 : array_update_84800[8];
  assign array_update_84813[9] = add_84176 == 32'h0000_0009 ? array_update_84811 : array_update_84800[9];
  assign array_index_84815 = array_update_72021[add_84812 > 32'h0000_0009 ? 4'h9 : add_84812[3:0]];
  assign array_index_84816 = array_update_84813[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_84820 = smul32b_32b_x_32b(array_index_84183[add_84812 > 32'h0000_0009 ? 4'h9 : add_84812[3:0]], array_index_84815[add_84719 > 32'h0000_0009 ? 4'h9 : add_84719[3:0]]);
  assign add_84822 = array_index_84816[add_84719 > 32'h0000_0009 ? 4'h9 : add_84719[3:0]] + smul_84820;
  assign array_update_84824[0] = add_84719 == 32'h0000_0000 ? add_84822 : array_index_84816[0];
  assign array_update_84824[1] = add_84719 == 32'h0000_0001 ? add_84822 : array_index_84816[1];
  assign array_update_84824[2] = add_84719 == 32'h0000_0002 ? add_84822 : array_index_84816[2];
  assign array_update_84824[3] = add_84719 == 32'h0000_0003 ? add_84822 : array_index_84816[3];
  assign array_update_84824[4] = add_84719 == 32'h0000_0004 ? add_84822 : array_index_84816[4];
  assign array_update_84824[5] = add_84719 == 32'h0000_0005 ? add_84822 : array_index_84816[5];
  assign array_update_84824[6] = add_84719 == 32'h0000_0006 ? add_84822 : array_index_84816[6];
  assign array_update_84824[7] = add_84719 == 32'h0000_0007 ? add_84822 : array_index_84816[7];
  assign array_update_84824[8] = add_84719 == 32'h0000_0008 ? add_84822 : array_index_84816[8];
  assign array_update_84824[9] = add_84719 == 32'h0000_0009 ? add_84822 : array_index_84816[9];
  assign add_84825 = add_84812 + 32'h0000_0001;
  assign array_update_84826[0] = add_84176 == 32'h0000_0000 ? array_update_84824 : array_update_84813[0];
  assign array_update_84826[1] = add_84176 == 32'h0000_0001 ? array_update_84824 : array_update_84813[1];
  assign array_update_84826[2] = add_84176 == 32'h0000_0002 ? array_update_84824 : array_update_84813[2];
  assign array_update_84826[3] = add_84176 == 32'h0000_0003 ? array_update_84824 : array_update_84813[3];
  assign array_update_84826[4] = add_84176 == 32'h0000_0004 ? array_update_84824 : array_update_84813[4];
  assign array_update_84826[5] = add_84176 == 32'h0000_0005 ? array_update_84824 : array_update_84813[5];
  assign array_update_84826[6] = add_84176 == 32'h0000_0006 ? array_update_84824 : array_update_84813[6];
  assign array_update_84826[7] = add_84176 == 32'h0000_0007 ? array_update_84824 : array_update_84813[7];
  assign array_update_84826[8] = add_84176 == 32'h0000_0008 ? array_update_84824 : array_update_84813[8];
  assign array_update_84826[9] = add_84176 == 32'h0000_0009 ? array_update_84824 : array_update_84813[9];
  assign array_index_84828 = array_update_72021[add_84825 > 32'h0000_0009 ? 4'h9 : add_84825[3:0]];
  assign array_index_84829 = array_update_84826[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_84833 = smul32b_32b_x_32b(array_index_84183[add_84825 > 32'h0000_0009 ? 4'h9 : add_84825[3:0]], array_index_84828[add_84719 > 32'h0000_0009 ? 4'h9 : add_84719[3:0]]);
  assign add_84835 = array_index_84829[add_84719 > 32'h0000_0009 ? 4'h9 : add_84719[3:0]] + smul_84833;
  assign array_update_84837[0] = add_84719 == 32'h0000_0000 ? add_84835 : array_index_84829[0];
  assign array_update_84837[1] = add_84719 == 32'h0000_0001 ? add_84835 : array_index_84829[1];
  assign array_update_84837[2] = add_84719 == 32'h0000_0002 ? add_84835 : array_index_84829[2];
  assign array_update_84837[3] = add_84719 == 32'h0000_0003 ? add_84835 : array_index_84829[3];
  assign array_update_84837[4] = add_84719 == 32'h0000_0004 ? add_84835 : array_index_84829[4];
  assign array_update_84837[5] = add_84719 == 32'h0000_0005 ? add_84835 : array_index_84829[5];
  assign array_update_84837[6] = add_84719 == 32'h0000_0006 ? add_84835 : array_index_84829[6];
  assign array_update_84837[7] = add_84719 == 32'h0000_0007 ? add_84835 : array_index_84829[7];
  assign array_update_84837[8] = add_84719 == 32'h0000_0008 ? add_84835 : array_index_84829[8];
  assign array_update_84837[9] = add_84719 == 32'h0000_0009 ? add_84835 : array_index_84829[9];
  assign add_84838 = add_84825 + 32'h0000_0001;
  assign array_update_84839[0] = add_84176 == 32'h0000_0000 ? array_update_84837 : array_update_84826[0];
  assign array_update_84839[1] = add_84176 == 32'h0000_0001 ? array_update_84837 : array_update_84826[1];
  assign array_update_84839[2] = add_84176 == 32'h0000_0002 ? array_update_84837 : array_update_84826[2];
  assign array_update_84839[3] = add_84176 == 32'h0000_0003 ? array_update_84837 : array_update_84826[3];
  assign array_update_84839[4] = add_84176 == 32'h0000_0004 ? array_update_84837 : array_update_84826[4];
  assign array_update_84839[5] = add_84176 == 32'h0000_0005 ? array_update_84837 : array_update_84826[5];
  assign array_update_84839[6] = add_84176 == 32'h0000_0006 ? array_update_84837 : array_update_84826[6];
  assign array_update_84839[7] = add_84176 == 32'h0000_0007 ? array_update_84837 : array_update_84826[7];
  assign array_update_84839[8] = add_84176 == 32'h0000_0008 ? array_update_84837 : array_update_84826[8];
  assign array_update_84839[9] = add_84176 == 32'h0000_0009 ? array_update_84837 : array_update_84826[9];
  assign array_index_84841 = array_update_72021[add_84838 > 32'h0000_0009 ? 4'h9 : add_84838[3:0]];
  assign array_index_84842 = array_update_84839[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_84846 = smul32b_32b_x_32b(array_index_84183[add_84838 > 32'h0000_0009 ? 4'h9 : add_84838[3:0]], array_index_84841[add_84719 > 32'h0000_0009 ? 4'h9 : add_84719[3:0]]);
  assign add_84848 = array_index_84842[add_84719 > 32'h0000_0009 ? 4'h9 : add_84719[3:0]] + smul_84846;
  assign array_update_84849[0] = add_84719 == 32'h0000_0000 ? add_84848 : array_index_84842[0];
  assign array_update_84849[1] = add_84719 == 32'h0000_0001 ? add_84848 : array_index_84842[1];
  assign array_update_84849[2] = add_84719 == 32'h0000_0002 ? add_84848 : array_index_84842[2];
  assign array_update_84849[3] = add_84719 == 32'h0000_0003 ? add_84848 : array_index_84842[3];
  assign array_update_84849[4] = add_84719 == 32'h0000_0004 ? add_84848 : array_index_84842[4];
  assign array_update_84849[5] = add_84719 == 32'h0000_0005 ? add_84848 : array_index_84842[5];
  assign array_update_84849[6] = add_84719 == 32'h0000_0006 ? add_84848 : array_index_84842[6];
  assign array_update_84849[7] = add_84719 == 32'h0000_0007 ? add_84848 : array_index_84842[7];
  assign array_update_84849[8] = add_84719 == 32'h0000_0008 ? add_84848 : array_index_84842[8];
  assign array_update_84849[9] = add_84719 == 32'h0000_0009 ? add_84848 : array_index_84842[9];
  assign array_update_84850[0] = add_84176 == 32'h0000_0000 ? array_update_84849 : array_update_84839[0];
  assign array_update_84850[1] = add_84176 == 32'h0000_0001 ? array_update_84849 : array_update_84839[1];
  assign array_update_84850[2] = add_84176 == 32'h0000_0002 ? array_update_84849 : array_update_84839[2];
  assign array_update_84850[3] = add_84176 == 32'h0000_0003 ? array_update_84849 : array_update_84839[3];
  assign array_update_84850[4] = add_84176 == 32'h0000_0004 ? array_update_84849 : array_update_84839[4];
  assign array_update_84850[5] = add_84176 == 32'h0000_0005 ? array_update_84849 : array_update_84839[5];
  assign array_update_84850[6] = add_84176 == 32'h0000_0006 ? array_update_84849 : array_update_84839[6];
  assign array_update_84850[7] = add_84176 == 32'h0000_0007 ? array_update_84849 : array_update_84839[7];
  assign array_update_84850[8] = add_84176 == 32'h0000_0008 ? array_update_84849 : array_update_84839[8];
  assign array_update_84850[9] = add_84176 == 32'h0000_0009 ? array_update_84849 : array_update_84839[9];
  assign array_index_84852 = array_update_84850[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign add_84854 = add_84719 + 32'h0000_0001;
  assign array_update_84855[0] = add_84854 == 32'h0000_0000 ? 32'h0000_0000 : array_index_84852[0];
  assign array_update_84855[1] = add_84854 == 32'h0000_0001 ? 32'h0000_0000 : array_index_84852[1];
  assign array_update_84855[2] = add_84854 == 32'h0000_0002 ? 32'h0000_0000 : array_index_84852[2];
  assign array_update_84855[3] = add_84854 == 32'h0000_0003 ? 32'h0000_0000 : array_index_84852[3];
  assign array_update_84855[4] = add_84854 == 32'h0000_0004 ? 32'h0000_0000 : array_index_84852[4];
  assign array_update_84855[5] = add_84854 == 32'h0000_0005 ? 32'h0000_0000 : array_index_84852[5];
  assign array_update_84855[6] = add_84854 == 32'h0000_0006 ? 32'h0000_0000 : array_index_84852[6];
  assign array_update_84855[7] = add_84854 == 32'h0000_0007 ? 32'h0000_0000 : array_index_84852[7];
  assign array_update_84855[8] = add_84854 == 32'h0000_0008 ? 32'h0000_0000 : array_index_84852[8];
  assign array_update_84855[9] = add_84854 == 32'h0000_0009 ? 32'h0000_0000 : array_index_84852[9];
  assign literal_84856 = 32'h0000_0000;
  assign array_update_84857[0] = add_84176 == 32'h0000_0000 ? array_update_84855 : array_update_84850[0];
  assign array_update_84857[1] = add_84176 == 32'h0000_0001 ? array_update_84855 : array_update_84850[1];
  assign array_update_84857[2] = add_84176 == 32'h0000_0002 ? array_update_84855 : array_update_84850[2];
  assign array_update_84857[3] = add_84176 == 32'h0000_0003 ? array_update_84855 : array_update_84850[3];
  assign array_update_84857[4] = add_84176 == 32'h0000_0004 ? array_update_84855 : array_update_84850[4];
  assign array_update_84857[5] = add_84176 == 32'h0000_0005 ? array_update_84855 : array_update_84850[5];
  assign array_update_84857[6] = add_84176 == 32'h0000_0006 ? array_update_84855 : array_update_84850[6];
  assign array_update_84857[7] = add_84176 == 32'h0000_0007 ? array_update_84855 : array_update_84850[7];
  assign array_update_84857[8] = add_84176 == 32'h0000_0008 ? array_update_84855 : array_update_84850[8];
  assign array_update_84857[9] = add_84176 == 32'h0000_0009 ? array_update_84855 : array_update_84850[9];
  assign array_index_84859 = array_update_72021[literal_84856 > 32'h0000_0009 ? 4'h9 : literal_84856[3:0]];
  assign array_index_84860 = array_update_84857[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_84864 = smul32b_32b_x_32b(array_index_84183[literal_84856 > 32'h0000_0009 ? 4'h9 : literal_84856[3:0]], array_index_84859[add_84854 > 32'h0000_0009 ? 4'h9 : add_84854[3:0]]);
  assign add_84866 = array_index_84860[add_84854 > 32'h0000_0009 ? 4'h9 : add_84854[3:0]] + smul_84864;
  assign array_update_84868[0] = add_84854 == 32'h0000_0000 ? add_84866 : array_index_84860[0];
  assign array_update_84868[1] = add_84854 == 32'h0000_0001 ? add_84866 : array_index_84860[1];
  assign array_update_84868[2] = add_84854 == 32'h0000_0002 ? add_84866 : array_index_84860[2];
  assign array_update_84868[3] = add_84854 == 32'h0000_0003 ? add_84866 : array_index_84860[3];
  assign array_update_84868[4] = add_84854 == 32'h0000_0004 ? add_84866 : array_index_84860[4];
  assign array_update_84868[5] = add_84854 == 32'h0000_0005 ? add_84866 : array_index_84860[5];
  assign array_update_84868[6] = add_84854 == 32'h0000_0006 ? add_84866 : array_index_84860[6];
  assign array_update_84868[7] = add_84854 == 32'h0000_0007 ? add_84866 : array_index_84860[7];
  assign array_update_84868[8] = add_84854 == 32'h0000_0008 ? add_84866 : array_index_84860[8];
  assign array_update_84868[9] = add_84854 == 32'h0000_0009 ? add_84866 : array_index_84860[9];
  assign add_84869 = literal_84856 + 32'h0000_0001;
  assign array_update_84870[0] = add_84176 == 32'h0000_0000 ? array_update_84868 : array_update_84857[0];
  assign array_update_84870[1] = add_84176 == 32'h0000_0001 ? array_update_84868 : array_update_84857[1];
  assign array_update_84870[2] = add_84176 == 32'h0000_0002 ? array_update_84868 : array_update_84857[2];
  assign array_update_84870[3] = add_84176 == 32'h0000_0003 ? array_update_84868 : array_update_84857[3];
  assign array_update_84870[4] = add_84176 == 32'h0000_0004 ? array_update_84868 : array_update_84857[4];
  assign array_update_84870[5] = add_84176 == 32'h0000_0005 ? array_update_84868 : array_update_84857[5];
  assign array_update_84870[6] = add_84176 == 32'h0000_0006 ? array_update_84868 : array_update_84857[6];
  assign array_update_84870[7] = add_84176 == 32'h0000_0007 ? array_update_84868 : array_update_84857[7];
  assign array_update_84870[8] = add_84176 == 32'h0000_0008 ? array_update_84868 : array_update_84857[8];
  assign array_update_84870[9] = add_84176 == 32'h0000_0009 ? array_update_84868 : array_update_84857[9];
  assign array_index_84872 = array_update_72021[add_84869 > 32'h0000_0009 ? 4'h9 : add_84869[3:0]];
  assign array_index_84873 = array_update_84870[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_84877 = smul32b_32b_x_32b(array_index_84183[add_84869 > 32'h0000_0009 ? 4'h9 : add_84869[3:0]], array_index_84872[add_84854 > 32'h0000_0009 ? 4'h9 : add_84854[3:0]]);
  assign add_84879 = array_index_84873[add_84854 > 32'h0000_0009 ? 4'h9 : add_84854[3:0]] + smul_84877;
  assign array_update_84881[0] = add_84854 == 32'h0000_0000 ? add_84879 : array_index_84873[0];
  assign array_update_84881[1] = add_84854 == 32'h0000_0001 ? add_84879 : array_index_84873[1];
  assign array_update_84881[2] = add_84854 == 32'h0000_0002 ? add_84879 : array_index_84873[2];
  assign array_update_84881[3] = add_84854 == 32'h0000_0003 ? add_84879 : array_index_84873[3];
  assign array_update_84881[4] = add_84854 == 32'h0000_0004 ? add_84879 : array_index_84873[4];
  assign array_update_84881[5] = add_84854 == 32'h0000_0005 ? add_84879 : array_index_84873[5];
  assign array_update_84881[6] = add_84854 == 32'h0000_0006 ? add_84879 : array_index_84873[6];
  assign array_update_84881[7] = add_84854 == 32'h0000_0007 ? add_84879 : array_index_84873[7];
  assign array_update_84881[8] = add_84854 == 32'h0000_0008 ? add_84879 : array_index_84873[8];
  assign array_update_84881[9] = add_84854 == 32'h0000_0009 ? add_84879 : array_index_84873[9];
  assign add_84882 = add_84869 + 32'h0000_0001;
  assign array_update_84883[0] = add_84176 == 32'h0000_0000 ? array_update_84881 : array_update_84870[0];
  assign array_update_84883[1] = add_84176 == 32'h0000_0001 ? array_update_84881 : array_update_84870[1];
  assign array_update_84883[2] = add_84176 == 32'h0000_0002 ? array_update_84881 : array_update_84870[2];
  assign array_update_84883[3] = add_84176 == 32'h0000_0003 ? array_update_84881 : array_update_84870[3];
  assign array_update_84883[4] = add_84176 == 32'h0000_0004 ? array_update_84881 : array_update_84870[4];
  assign array_update_84883[5] = add_84176 == 32'h0000_0005 ? array_update_84881 : array_update_84870[5];
  assign array_update_84883[6] = add_84176 == 32'h0000_0006 ? array_update_84881 : array_update_84870[6];
  assign array_update_84883[7] = add_84176 == 32'h0000_0007 ? array_update_84881 : array_update_84870[7];
  assign array_update_84883[8] = add_84176 == 32'h0000_0008 ? array_update_84881 : array_update_84870[8];
  assign array_update_84883[9] = add_84176 == 32'h0000_0009 ? array_update_84881 : array_update_84870[9];
  assign array_index_84885 = array_update_72021[add_84882 > 32'h0000_0009 ? 4'h9 : add_84882[3:0]];
  assign array_index_84886 = array_update_84883[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_84890 = smul32b_32b_x_32b(array_index_84183[add_84882 > 32'h0000_0009 ? 4'h9 : add_84882[3:0]], array_index_84885[add_84854 > 32'h0000_0009 ? 4'h9 : add_84854[3:0]]);
  assign add_84892 = array_index_84886[add_84854 > 32'h0000_0009 ? 4'h9 : add_84854[3:0]] + smul_84890;
  assign array_update_84894[0] = add_84854 == 32'h0000_0000 ? add_84892 : array_index_84886[0];
  assign array_update_84894[1] = add_84854 == 32'h0000_0001 ? add_84892 : array_index_84886[1];
  assign array_update_84894[2] = add_84854 == 32'h0000_0002 ? add_84892 : array_index_84886[2];
  assign array_update_84894[3] = add_84854 == 32'h0000_0003 ? add_84892 : array_index_84886[3];
  assign array_update_84894[4] = add_84854 == 32'h0000_0004 ? add_84892 : array_index_84886[4];
  assign array_update_84894[5] = add_84854 == 32'h0000_0005 ? add_84892 : array_index_84886[5];
  assign array_update_84894[6] = add_84854 == 32'h0000_0006 ? add_84892 : array_index_84886[6];
  assign array_update_84894[7] = add_84854 == 32'h0000_0007 ? add_84892 : array_index_84886[7];
  assign array_update_84894[8] = add_84854 == 32'h0000_0008 ? add_84892 : array_index_84886[8];
  assign array_update_84894[9] = add_84854 == 32'h0000_0009 ? add_84892 : array_index_84886[9];
  assign add_84895 = add_84882 + 32'h0000_0001;
  assign array_update_84896[0] = add_84176 == 32'h0000_0000 ? array_update_84894 : array_update_84883[0];
  assign array_update_84896[1] = add_84176 == 32'h0000_0001 ? array_update_84894 : array_update_84883[1];
  assign array_update_84896[2] = add_84176 == 32'h0000_0002 ? array_update_84894 : array_update_84883[2];
  assign array_update_84896[3] = add_84176 == 32'h0000_0003 ? array_update_84894 : array_update_84883[3];
  assign array_update_84896[4] = add_84176 == 32'h0000_0004 ? array_update_84894 : array_update_84883[4];
  assign array_update_84896[5] = add_84176 == 32'h0000_0005 ? array_update_84894 : array_update_84883[5];
  assign array_update_84896[6] = add_84176 == 32'h0000_0006 ? array_update_84894 : array_update_84883[6];
  assign array_update_84896[7] = add_84176 == 32'h0000_0007 ? array_update_84894 : array_update_84883[7];
  assign array_update_84896[8] = add_84176 == 32'h0000_0008 ? array_update_84894 : array_update_84883[8];
  assign array_update_84896[9] = add_84176 == 32'h0000_0009 ? array_update_84894 : array_update_84883[9];
  assign array_index_84898 = array_update_72021[add_84895 > 32'h0000_0009 ? 4'h9 : add_84895[3:0]];
  assign array_index_84899 = array_update_84896[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_84903 = smul32b_32b_x_32b(array_index_84183[add_84895 > 32'h0000_0009 ? 4'h9 : add_84895[3:0]], array_index_84898[add_84854 > 32'h0000_0009 ? 4'h9 : add_84854[3:0]]);
  assign add_84905 = array_index_84899[add_84854 > 32'h0000_0009 ? 4'h9 : add_84854[3:0]] + smul_84903;
  assign array_update_84907[0] = add_84854 == 32'h0000_0000 ? add_84905 : array_index_84899[0];
  assign array_update_84907[1] = add_84854 == 32'h0000_0001 ? add_84905 : array_index_84899[1];
  assign array_update_84907[2] = add_84854 == 32'h0000_0002 ? add_84905 : array_index_84899[2];
  assign array_update_84907[3] = add_84854 == 32'h0000_0003 ? add_84905 : array_index_84899[3];
  assign array_update_84907[4] = add_84854 == 32'h0000_0004 ? add_84905 : array_index_84899[4];
  assign array_update_84907[5] = add_84854 == 32'h0000_0005 ? add_84905 : array_index_84899[5];
  assign array_update_84907[6] = add_84854 == 32'h0000_0006 ? add_84905 : array_index_84899[6];
  assign array_update_84907[7] = add_84854 == 32'h0000_0007 ? add_84905 : array_index_84899[7];
  assign array_update_84907[8] = add_84854 == 32'h0000_0008 ? add_84905 : array_index_84899[8];
  assign array_update_84907[9] = add_84854 == 32'h0000_0009 ? add_84905 : array_index_84899[9];
  assign add_84908 = add_84895 + 32'h0000_0001;
  assign array_update_84909[0] = add_84176 == 32'h0000_0000 ? array_update_84907 : array_update_84896[0];
  assign array_update_84909[1] = add_84176 == 32'h0000_0001 ? array_update_84907 : array_update_84896[1];
  assign array_update_84909[2] = add_84176 == 32'h0000_0002 ? array_update_84907 : array_update_84896[2];
  assign array_update_84909[3] = add_84176 == 32'h0000_0003 ? array_update_84907 : array_update_84896[3];
  assign array_update_84909[4] = add_84176 == 32'h0000_0004 ? array_update_84907 : array_update_84896[4];
  assign array_update_84909[5] = add_84176 == 32'h0000_0005 ? array_update_84907 : array_update_84896[5];
  assign array_update_84909[6] = add_84176 == 32'h0000_0006 ? array_update_84907 : array_update_84896[6];
  assign array_update_84909[7] = add_84176 == 32'h0000_0007 ? array_update_84907 : array_update_84896[7];
  assign array_update_84909[8] = add_84176 == 32'h0000_0008 ? array_update_84907 : array_update_84896[8];
  assign array_update_84909[9] = add_84176 == 32'h0000_0009 ? array_update_84907 : array_update_84896[9];
  assign array_index_84911 = array_update_72021[add_84908 > 32'h0000_0009 ? 4'h9 : add_84908[3:0]];
  assign array_index_84912 = array_update_84909[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_84916 = smul32b_32b_x_32b(array_index_84183[add_84908 > 32'h0000_0009 ? 4'h9 : add_84908[3:0]], array_index_84911[add_84854 > 32'h0000_0009 ? 4'h9 : add_84854[3:0]]);
  assign add_84918 = array_index_84912[add_84854 > 32'h0000_0009 ? 4'h9 : add_84854[3:0]] + smul_84916;
  assign array_update_84920[0] = add_84854 == 32'h0000_0000 ? add_84918 : array_index_84912[0];
  assign array_update_84920[1] = add_84854 == 32'h0000_0001 ? add_84918 : array_index_84912[1];
  assign array_update_84920[2] = add_84854 == 32'h0000_0002 ? add_84918 : array_index_84912[2];
  assign array_update_84920[3] = add_84854 == 32'h0000_0003 ? add_84918 : array_index_84912[3];
  assign array_update_84920[4] = add_84854 == 32'h0000_0004 ? add_84918 : array_index_84912[4];
  assign array_update_84920[5] = add_84854 == 32'h0000_0005 ? add_84918 : array_index_84912[5];
  assign array_update_84920[6] = add_84854 == 32'h0000_0006 ? add_84918 : array_index_84912[6];
  assign array_update_84920[7] = add_84854 == 32'h0000_0007 ? add_84918 : array_index_84912[7];
  assign array_update_84920[8] = add_84854 == 32'h0000_0008 ? add_84918 : array_index_84912[8];
  assign array_update_84920[9] = add_84854 == 32'h0000_0009 ? add_84918 : array_index_84912[9];
  assign add_84921 = add_84908 + 32'h0000_0001;
  assign array_update_84922[0] = add_84176 == 32'h0000_0000 ? array_update_84920 : array_update_84909[0];
  assign array_update_84922[1] = add_84176 == 32'h0000_0001 ? array_update_84920 : array_update_84909[1];
  assign array_update_84922[2] = add_84176 == 32'h0000_0002 ? array_update_84920 : array_update_84909[2];
  assign array_update_84922[3] = add_84176 == 32'h0000_0003 ? array_update_84920 : array_update_84909[3];
  assign array_update_84922[4] = add_84176 == 32'h0000_0004 ? array_update_84920 : array_update_84909[4];
  assign array_update_84922[5] = add_84176 == 32'h0000_0005 ? array_update_84920 : array_update_84909[5];
  assign array_update_84922[6] = add_84176 == 32'h0000_0006 ? array_update_84920 : array_update_84909[6];
  assign array_update_84922[7] = add_84176 == 32'h0000_0007 ? array_update_84920 : array_update_84909[7];
  assign array_update_84922[8] = add_84176 == 32'h0000_0008 ? array_update_84920 : array_update_84909[8];
  assign array_update_84922[9] = add_84176 == 32'h0000_0009 ? array_update_84920 : array_update_84909[9];
  assign array_index_84924 = array_update_72021[add_84921 > 32'h0000_0009 ? 4'h9 : add_84921[3:0]];
  assign array_index_84925 = array_update_84922[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_84929 = smul32b_32b_x_32b(array_index_84183[add_84921 > 32'h0000_0009 ? 4'h9 : add_84921[3:0]], array_index_84924[add_84854 > 32'h0000_0009 ? 4'h9 : add_84854[3:0]]);
  assign add_84931 = array_index_84925[add_84854 > 32'h0000_0009 ? 4'h9 : add_84854[3:0]] + smul_84929;
  assign array_update_84933[0] = add_84854 == 32'h0000_0000 ? add_84931 : array_index_84925[0];
  assign array_update_84933[1] = add_84854 == 32'h0000_0001 ? add_84931 : array_index_84925[1];
  assign array_update_84933[2] = add_84854 == 32'h0000_0002 ? add_84931 : array_index_84925[2];
  assign array_update_84933[3] = add_84854 == 32'h0000_0003 ? add_84931 : array_index_84925[3];
  assign array_update_84933[4] = add_84854 == 32'h0000_0004 ? add_84931 : array_index_84925[4];
  assign array_update_84933[5] = add_84854 == 32'h0000_0005 ? add_84931 : array_index_84925[5];
  assign array_update_84933[6] = add_84854 == 32'h0000_0006 ? add_84931 : array_index_84925[6];
  assign array_update_84933[7] = add_84854 == 32'h0000_0007 ? add_84931 : array_index_84925[7];
  assign array_update_84933[8] = add_84854 == 32'h0000_0008 ? add_84931 : array_index_84925[8];
  assign array_update_84933[9] = add_84854 == 32'h0000_0009 ? add_84931 : array_index_84925[9];
  assign add_84934 = add_84921 + 32'h0000_0001;
  assign array_update_84935[0] = add_84176 == 32'h0000_0000 ? array_update_84933 : array_update_84922[0];
  assign array_update_84935[1] = add_84176 == 32'h0000_0001 ? array_update_84933 : array_update_84922[1];
  assign array_update_84935[2] = add_84176 == 32'h0000_0002 ? array_update_84933 : array_update_84922[2];
  assign array_update_84935[3] = add_84176 == 32'h0000_0003 ? array_update_84933 : array_update_84922[3];
  assign array_update_84935[4] = add_84176 == 32'h0000_0004 ? array_update_84933 : array_update_84922[4];
  assign array_update_84935[5] = add_84176 == 32'h0000_0005 ? array_update_84933 : array_update_84922[5];
  assign array_update_84935[6] = add_84176 == 32'h0000_0006 ? array_update_84933 : array_update_84922[6];
  assign array_update_84935[7] = add_84176 == 32'h0000_0007 ? array_update_84933 : array_update_84922[7];
  assign array_update_84935[8] = add_84176 == 32'h0000_0008 ? array_update_84933 : array_update_84922[8];
  assign array_update_84935[9] = add_84176 == 32'h0000_0009 ? array_update_84933 : array_update_84922[9];
  assign array_index_84937 = array_update_72021[add_84934 > 32'h0000_0009 ? 4'h9 : add_84934[3:0]];
  assign array_index_84938 = array_update_84935[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_84942 = smul32b_32b_x_32b(array_index_84183[add_84934 > 32'h0000_0009 ? 4'h9 : add_84934[3:0]], array_index_84937[add_84854 > 32'h0000_0009 ? 4'h9 : add_84854[3:0]]);
  assign add_84944 = array_index_84938[add_84854 > 32'h0000_0009 ? 4'h9 : add_84854[3:0]] + smul_84942;
  assign array_update_84946[0] = add_84854 == 32'h0000_0000 ? add_84944 : array_index_84938[0];
  assign array_update_84946[1] = add_84854 == 32'h0000_0001 ? add_84944 : array_index_84938[1];
  assign array_update_84946[2] = add_84854 == 32'h0000_0002 ? add_84944 : array_index_84938[2];
  assign array_update_84946[3] = add_84854 == 32'h0000_0003 ? add_84944 : array_index_84938[3];
  assign array_update_84946[4] = add_84854 == 32'h0000_0004 ? add_84944 : array_index_84938[4];
  assign array_update_84946[5] = add_84854 == 32'h0000_0005 ? add_84944 : array_index_84938[5];
  assign array_update_84946[6] = add_84854 == 32'h0000_0006 ? add_84944 : array_index_84938[6];
  assign array_update_84946[7] = add_84854 == 32'h0000_0007 ? add_84944 : array_index_84938[7];
  assign array_update_84946[8] = add_84854 == 32'h0000_0008 ? add_84944 : array_index_84938[8];
  assign array_update_84946[9] = add_84854 == 32'h0000_0009 ? add_84944 : array_index_84938[9];
  assign add_84947 = add_84934 + 32'h0000_0001;
  assign array_update_84948[0] = add_84176 == 32'h0000_0000 ? array_update_84946 : array_update_84935[0];
  assign array_update_84948[1] = add_84176 == 32'h0000_0001 ? array_update_84946 : array_update_84935[1];
  assign array_update_84948[2] = add_84176 == 32'h0000_0002 ? array_update_84946 : array_update_84935[2];
  assign array_update_84948[3] = add_84176 == 32'h0000_0003 ? array_update_84946 : array_update_84935[3];
  assign array_update_84948[4] = add_84176 == 32'h0000_0004 ? array_update_84946 : array_update_84935[4];
  assign array_update_84948[5] = add_84176 == 32'h0000_0005 ? array_update_84946 : array_update_84935[5];
  assign array_update_84948[6] = add_84176 == 32'h0000_0006 ? array_update_84946 : array_update_84935[6];
  assign array_update_84948[7] = add_84176 == 32'h0000_0007 ? array_update_84946 : array_update_84935[7];
  assign array_update_84948[8] = add_84176 == 32'h0000_0008 ? array_update_84946 : array_update_84935[8];
  assign array_update_84948[9] = add_84176 == 32'h0000_0009 ? array_update_84946 : array_update_84935[9];
  assign array_index_84950 = array_update_72021[add_84947 > 32'h0000_0009 ? 4'h9 : add_84947[3:0]];
  assign array_index_84951 = array_update_84948[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_84955 = smul32b_32b_x_32b(array_index_84183[add_84947 > 32'h0000_0009 ? 4'h9 : add_84947[3:0]], array_index_84950[add_84854 > 32'h0000_0009 ? 4'h9 : add_84854[3:0]]);
  assign add_84957 = array_index_84951[add_84854 > 32'h0000_0009 ? 4'h9 : add_84854[3:0]] + smul_84955;
  assign array_update_84959[0] = add_84854 == 32'h0000_0000 ? add_84957 : array_index_84951[0];
  assign array_update_84959[1] = add_84854 == 32'h0000_0001 ? add_84957 : array_index_84951[1];
  assign array_update_84959[2] = add_84854 == 32'h0000_0002 ? add_84957 : array_index_84951[2];
  assign array_update_84959[3] = add_84854 == 32'h0000_0003 ? add_84957 : array_index_84951[3];
  assign array_update_84959[4] = add_84854 == 32'h0000_0004 ? add_84957 : array_index_84951[4];
  assign array_update_84959[5] = add_84854 == 32'h0000_0005 ? add_84957 : array_index_84951[5];
  assign array_update_84959[6] = add_84854 == 32'h0000_0006 ? add_84957 : array_index_84951[6];
  assign array_update_84959[7] = add_84854 == 32'h0000_0007 ? add_84957 : array_index_84951[7];
  assign array_update_84959[8] = add_84854 == 32'h0000_0008 ? add_84957 : array_index_84951[8];
  assign array_update_84959[9] = add_84854 == 32'h0000_0009 ? add_84957 : array_index_84951[9];
  assign add_84960 = add_84947 + 32'h0000_0001;
  assign array_update_84961[0] = add_84176 == 32'h0000_0000 ? array_update_84959 : array_update_84948[0];
  assign array_update_84961[1] = add_84176 == 32'h0000_0001 ? array_update_84959 : array_update_84948[1];
  assign array_update_84961[2] = add_84176 == 32'h0000_0002 ? array_update_84959 : array_update_84948[2];
  assign array_update_84961[3] = add_84176 == 32'h0000_0003 ? array_update_84959 : array_update_84948[3];
  assign array_update_84961[4] = add_84176 == 32'h0000_0004 ? array_update_84959 : array_update_84948[4];
  assign array_update_84961[5] = add_84176 == 32'h0000_0005 ? array_update_84959 : array_update_84948[5];
  assign array_update_84961[6] = add_84176 == 32'h0000_0006 ? array_update_84959 : array_update_84948[6];
  assign array_update_84961[7] = add_84176 == 32'h0000_0007 ? array_update_84959 : array_update_84948[7];
  assign array_update_84961[8] = add_84176 == 32'h0000_0008 ? array_update_84959 : array_update_84948[8];
  assign array_update_84961[9] = add_84176 == 32'h0000_0009 ? array_update_84959 : array_update_84948[9];
  assign array_index_84963 = array_update_72021[add_84960 > 32'h0000_0009 ? 4'h9 : add_84960[3:0]];
  assign array_index_84964 = array_update_84961[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_84968 = smul32b_32b_x_32b(array_index_84183[add_84960 > 32'h0000_0009 ? 4'h9 : add_84960[3:0]], array_index_84963[add_84854 > 32'h0000_0009 ? 4'h9 : add_84854[3:0]]);
  assign add_84970 = array_index_84964[add_84854 > 32'h0000_0009 ? 4'h9 : add_84854[3:0]] + smul_84968;
  assign array_update_84972[0] = add_84854 == 32'h0000_0000 ? add_84970 : array_index_84964[0];
  assign array_update_84972[1] = add_84854 == 32'h0000_0001 ? add_84970 : array_index_84964[1];
  assign array_update_84972[2] = add_84854 == 32'h0000_0002 ? add_84970 : array_index_84964[2];
  assign array_update_84972[3] = add_84854 == 32'h0000_0003 ? add_84970 : array_index_84964[3];
  assign array_update_84972[4] = add_84854 == 32'h0000_0004 ? add_84970 : array_index_84964[4];
  assign array_update_84972[5] = add_84854 == 32'h0000_0005 ? add_84970 : array_index_84964[5];
  assign array_update_84972[6] = add_84854 == 32'h0000_0006 ? add_84970 : array_index_84964[6];
  assign array_update_84972[7] = add_84854 == 32'h0000_0007 ? add_84970 : array_index_84964[7];
  assign array_update_84972[8] = add_84854 == 32'h0000_0008 ? add_84970 : array_index_84964[8];
  assign array_update_84972[9] = add_84854 == 32'h0000_0009 ? add_84970 : array_index_84964[9];
  assign add_84973 = add_84960 + 32'h0000_0001;
  assign array_update_84974[0] = add_84176 == 32'h0000_0000 ? array_update_84972 : array_update_84961[0];
  assign array_update_84974[1] = add_84176 == 32'h0000_0001 ? array_update_84972 : array_update_84961[1];
  assign array_update_84974[2] = add_84176 == 32'h0000_0002 ? array_update_84972 : array_update_84961[2];
  assign array_update_84974[3] = add_84176 == 32'h0000_0003 ? array_update_84972 : array_update_84961[3];
  assign array_update_84974[4] = add_84176 == 32'h0000_0004 ? array_update_84972 : array_update_84961[4];
  assign array_update_84974[5] = add_84176 == 32'h0000_0005 ? array_update_84972 : array_update_84961[5];
  assign array_update_84974[6] = add_84176 == 32'h0000_0006 ? array_update_84972 : array_update_84961[6];
  assign array_update_84974[7] = add_84176 == 32'h0000_0007 ? array_update_84972 : array_update_84961[7];
  assign array_update_84974[8] = add_84176 == 32'h0000_0008 ? array_update_84972 : array_update_84961[8];
  assign array_update_84974[9] = add_84176 == 32'h0000_0009 ? array_update_84972 : array_update_84961[9];
  assign array_index_84976 = array_update_72021[add_84973 > 32'h0000_0009 ? 4'h9 : add_84973[3:0]];
  assign array_index_84977 = array_update_84974[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_84981 = smul32b_32b_x_32b(array_index_84183[add_84973 > 32'h0000_0009 ? 4'h9 : add_84973[3:0]], array_index_84976[add_84854 > 32'h0000_0009 ? 4'h9 : add_84854[3:0]]);
  assign add_84983 = array_index_84977[add_84854 > 32'h0000_0009 ? 4'h9 : add_84854[3:0]] + smul_84981;
  assign array_update_84984[0] = add_84854 == 32'h0000_0000 ? add_84983 : array_index_84977[0];
  assign array_update_84984[1] = add_84854 == 32'h0000_0001 ? add_84983 : array_index_84977[1];
  assign array_update_84984[2] = add_84854 == 32'h0000_0002 ? add_84983 : array_index_84977[2];
  assign array_update_84984[3] = add_84854 == 32'h0000_0003 ? add_84983 : array_index_84977[3];
  assign array_update_84984[4] = add_84854 == 32'h0000_0004 ? add_84983 : array_index_84977[4];
  assign array_update_84984[5] = add_84854 == 32'h0000_0005 ? add_84983 : array_index_84977[5];
  assign array_update_84984[6] = add_84854 == 32'h0000_0006 ? add_84983 : array_index_84977[6];
  assign array_update_84984[7] = add_84854 == 32'h0000_0007 ? add_84983 : array_index_84977[7];
  assign array_update_84984[8] = add_84854 == 32'h0000_0008 ? add_84983 : array_index_84977[8];
  assign array_update_84984[9] = add_84854 == 32'h0000_0009 ? add_84983 : array_index_84977[9];
  assign array_update_84985[0] = add_84176 == 32'h0000_0000 ? array_update_84984 : array_update_84974[0];
  assign array_update_84985[1] = add_84176 == 32'h0000_0001 ? array_update_84984 : array_update_84974[1];
  assign array_update_84985[2] = add_84176 == 32'h0000_0002 ? array_update_84984 : array_update_84974[2];
  assign array_update_84985[3] = add_84176 == 32'h0000_0003 ? array_update_84984 : array_update_84974[3];
  assign array_update_84985[4] = add_84176 == 32'h0000_0004 ? array_update_84984 : array_update_84974[4];
  assign array_update_84985[5] = add_84176 == 32'h0000_0005 ? array_update_84984 : array_update_84974[5];
  assign array_update_84985[6] = add_84176 == 32'h0000_0006 ? array_update_84984 : array_update_84974[6];
  assign array_update_84985[7] = add_84176 == 32'h0000_0007 ? array_update_84984 : array_update_84974[7];
  assign array_update_84985[8] = add_84176 == 32'h0000_0008 ? array_update_84984 : array_update_84974[8];
  assign array_update_84985[9] = add_84176 == 32'h0000_0009 ? array_update_84984 : array_update_84974[9];
  assign array_index_84987 = array_update_84985[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign add_84989 = add_84854 + 32'h0000_0001;
  assign array_update_84990[0] = add_84989 == 32'h0000_0000 ? 32'h0000_0000 : array_index_84987[0];
  assign array_update_84990[1] = add_84989 == 32'h0000_0001 ? 32'h0000_0000 : array_index_84987[1];
  assign array_update_84990[2] = add_84989 == 32'h0000_0002 ? 32'h0000_0000 : array_index_84987[2];
  assign array_update_84990[3] = add_84989 == 32'h0000_0003 ? 32'h0000_0000 : array_index_84987[3];
  assign array_update_84990[4] = add_84989 == 32'h0000_0004 ? 32'h0000_0000 : array_index_84987[4];
  assign array_update_84990[5] = add_84989 == 32'h0000_0005 ? 32'h0000_0000 : array_index_84987[5];
  assign array_update_84990[6] = add_84989 == 32'h0000_0006 ? 32'h0000_0000 : array_index_84987[6];
  assign array_update_84990[7] = add_84989 == 32'h0000_0007 ? 32'h0000_0000 : array_index_84987[7];
  assign array_update_84990[8] = add_84989 == 32'h0000_0008 ? 32'h0000_0000 : array_index_84987[8];
  assign array_update_84990[9] = add_84989 == 32'h0000_0009 ? 32'h0000_0000 : array_index_84987[9];
  assign literal_84991 = 32'h0000_0000;
  assign array_update_84992[0] = add_84176 == 32'h0000_0000 ? array_update_84990 : array_update_84985[0];
  assign array_update_84992[1] = add_84176 == 32'h0000_0001 ? array_update_84990 : array_update_84985[1];
  assign array_update_84992[2] = add_84176 == 32'h0000_0002 ? array_update_84990 : array_update_84985[2];
  assign array_update_84992[3] = add_84176 == 32'h0000_0003 ? array_update_84990 : array_update_84985[3];
  assign array_update_84992[4] = add_84176 == 32'h0000_0004 ? array_update_84990 : array_update_84985[4];
  assign array_update_84992[5] = add_84176 == 32'h0000_0005 ? array_update_84990 : array_update_84985[5];
  assign array_update_84992[6] = add_84176 == 32'h0000_0006 ? array_update_84990 : array_update_84985[6];
  assign array_update_84992[7] = add_84176 == 32'h0000_0007 ? array_update_84990 : array_update_84985[7];
  assign array_update_84992[8] = add_84176 == 32'h0000_0008 ? array_update_84990 : array_update_84985[8];
  assign array_update_84992[9] = add_84176 == 32'h0000_0009 ? array_update_84990 : array_update_84985[9];
  assign array_index_84994 = array_update_72021[literal_84991 > 32'h0000_0009 ? 4'h9 : literal_84991[3:0]];
  assign array_index_84995 = array_update_84992[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_84999 = smul32b_32b_x_32b(array_index_84183[literal_84991 > 32'h0000_0009 ? 4'h9 : literal_84991[3:0]], array_index_84994[add_84989 > 32'h0000_0009 ? 4'h9 : add_84989[3:0]]);
  assign add_85001 = array_index_84995[add_84989 > 32'h0000_0009 ? 4'h9 : add_84989[3:0]] + smul_84999;
  assign array_update_85003[0] = add_84989 == 32'h0000_0000 ? add_85001 : array_index_84995[0];
  assign array_update_85003[1] = add_84989 == 32'h0000_0001 ? add_85001 : array_index_84995[1];
  assign array_update_85003[2] = add_84989 == 32'h0000_0002 ? add_85001 : array_index_84995[2];
  assign array_update_85003[3] = add_84989 == 32'h0000_0003 ? add_85001 : array_index_84995[3];
  assign array_update_85003[4] = add_84989 == 32'h0000_0004 ? add_85001 : array_index_84995[4];
  assign array_update_85003[5] = add_84989 == 32'h0000_0005 ? add_85001 : array_index_84995[5];
  assign array_update_85003[6] = add_84989 == 32'h0000_0006 ? add_85001 : array_index_84995[6];
  assign array_update_85003[7] = add_84989 == 32'h0000_0007 ? add_85001 : array_index_84995[7];
  assign array_update_85003[8] = add_84989 == 32'h0000_0008 ? add_85001 : array_index_84995[8];
  assign array_update_85003[9] = add_84989 == 32'h0000_0009 ? add_85001 : array_index_84995[9];
  assign add_85004 = literal_84991 + 32'h0000_0001;
  assign array_update_85005[0] = add_84176 == 32'h0000_0000 ? array_update_85003 : array_update_84992[0];
  assign array_update_85005[1] = add_84176 == 32'h0000_0001 ? array_update_85003 : array_update_84992[1];
  assign array_update_85005[2] = add_84176 == 32'h0000_0002 ? array_update_85003 : array_update_84992[2];
  assign array_update_85005[3] = add_84176 == 32'h0000_0003 ? array_update_85003 : array_update_84992[3];
  assign array_update_85005[4] = add_84176 == 32'h0000_0004 ? array_update_85003 : array_update_84992[4];
  assign array_update_85005[5] = add_84176 == 32'h0000_0005 ? array_update_85003 : array_update_84992[5];
  assign array_update_85005[6] = add_84176 == 32'h0000_0006 ? array_update_85003 : array_update_84992[6];
  assign array_update_85005[7] = add_84176 == 32'h0000_0007 ? array_update_85003 : array_update_84992[7];
  assign array_update_85005[8] = add_84176 == 32'h0000_0008 ? array_update_85003 : array_update_84992[8];
  assign array_update_85005[9] = add_84176 == 32'h0000_0009 ? array_update_85003 : array_update_84992[9];
  assign array_index_85007 = array_update_72021[add_85004 > 32'h0000_0009 ? 4'h9 : add_85004[3:0]];
  assign array_index_85008 = array_update_85005[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_85012 = smul32b_32b_x_32b(array_index_84183[add_85004 > 32'h0000_0009 ? 4'h9 : add_85004[3:0]], array_index_85007[add_84989 > 32'h0000_0009 ? 4'h9 : add_84989[3:0]]);
  assign add_85014 = array_index_85008[add_84989 > 32'h0000_0009 ? 4'h9 : add_84989[3:0]] + smul_85012;
  assign array_update_85016[0] = add_84989 == 32'h0000_0000 ? add_85014 : array_index_85008[0];
  assign array_update_85016[1] = add_84989 == 32'h0000_0001 ? add_85014 : array_index_85008[1];
  assign array_update_85016[2] = add_84989 == 32'h0000_0002 ? add_85014 : array_index_85008[2];
  assign array_update_85016[3] = add_84989 == 32'h0000_0003 ? add_85014 : array_index_85008[3];
  assign array_update_85016[4] = add_84989 == 32'h0000_0004 ? add_85014 : array_index_85008[4];
  assign array_update_85016[5] = add_84989 == 32'h0000_0005 ? add_85014 : array_index_85008[5];
  assign array_update_85016[6] = add_84989 == 32'h0000_0006 ? add_85014 : array_index_85008[6];
  assign array_update_85016[7] = add_84989 == 32'h0000_0007 ? add_85014 : array_index_85008[7];
  assign array_update_85016[8] = add_84989 == 32'h0000_0008 ? add_85014 : array_index_85008[8];
  assign array_update_85016[9] = add_84989 == 32'h0000_0009 ? add_85014 : array_index_85008[9];
  assign add_85017 = add_85004 + 32'h0000_0001;
  assign array_update_85018[0] = add_84176 == 32'h0000_0000 ? array_update_85016 : array_update_85005[0];
  assign array_update_85018[1] = add_84176 == 32'h0000_0001 ? array_update_85016 : array_update_85005[1];
  assign array_update_85018[2] = add_84176 == 32'h0000_0002 ? array_update_85016 : array_update_85005[2];
  assign array_update_85018[3] = add_84176 == 32'h0000_0003 ? array_update_85016 : array_update_85005[3];
  assign array_update_85018[4] = add_84176 == 32'h0000_0004 ? array_update_85016 : array_update_85005[4];
  assign array_update_85018[5] = add_84176 == 32'h0000_0005 ? array_update_85016 : array_update_85005[5];
  assign array_update_85018[6] = add_84176 == 32'h0000_0006 ? array_update_85016 : array_update_85005[6];
  assign array_update_85018[7] = add_84176 == 32'h0000_0007 ? array_update_85016 : array_update_85005[7];
  assign array_update_85018[8] = add_84176 == 32'h0000_0008 ? array_update_85016 : array_update_85005[8];
  assign array_update_85018[9] = add_84176 == 32'h0000_0009 ? array_update_85016 : array_update_85005[9];
  assign array_index_85020 = array_update_72021[add_85017 > 32'h0000_0009 ? 4'h9 : add_85017[3:0]];
  assign array_index_85021 = array_update_85018[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_85025 = smul32b_32b_x_32b(array_index_84183[add_85017 > 32'h0000_0009 ? 4'h9 : add_85017[3:0]], array_index_85020[add_84989 > 32'h0000_0009 ? 4'h9 : add_84989[3:0]]);
  assign add_85027 = array_index_85021[add_84989 > 32'h0000_0009 ? 4'h9 : add_84989[3:0]] + smul_85025;
  assign array_update_85029[0] = add_84989 == 32'h0000_0000 ? add_85027 : array_index_85021[0];
  assign array_update_85029[1] = add_84989 == 32'h0000_0001 ? add_85027 : array_index_85021[1];
  assign array_update_85029[2] = add_84989 == 32'h0000_0002 ? add_85027 : array_index_85021[2];
  assign array_update_85029[3] = add_84989 == 32'h0000_0003 ? add_85027 : array_index_85021[3];
  assign array_update_85029[4] = add_84989 == 32'h0000_0004 ? add_85027 : array_index_85021[4];
  assign array_update_85029[5] = add_84989 == 32'h0000_0005 ? add_85027 : array_index_85021[5];
  assign array_update_85029[6] = add_84989 == 32'h0000_0006 ? add_85027 : array_index_85021[6];
  assign array_update_85029[7] = add_84989 == 32'h0000_0007 ? add_85027 : array_index_85021[7];
  assign array_update_85029[8] = add_84989 == 32'h0000_0008 ? add_85027 : array_index_85021[8];
  assign array_update_85029[9] = add_84989 == 32'h0000_0009 ? add_85027 : array_index_85021[9];
  assign add_85030 = add_85017 + 32'h0000_0001;
  assign array_update_85031[0] = add_84176 == 32'h0000_0000 ? array_update_85029 : array_update_85018[0];
  assign array_update_85031[1] = add_84176 == 32'h0000_0001 ? array_update_85029 : array_update_85018[1];
  assign array_update_85031[2] = add_84176 == 32'h0000_0002 ? array_update_85029 : array_update_85018[2];
  assign array_update_85031[3] = add_84176 == 32'h0000_0003 ? array_update_85029 : array_update_85018[3];
  assign array_update_85031[4] = add_84176 == 32'h0000_0004 ? array_update_85029 : array_update_85018[4];
  assign array_update_85031[5] = add_84176 == 32'h0000_0005 ? array_update_85029 : array_update_85018[5];
  assign array_update_85031[6] = add_84176 == 32'h0000_0006 ? array_update_85029 : array_update_85018[6];
  assign array_update_85031[7] = add_84176 == 32'h0000_0007 ? array_update_85029 : array_update_85018[7];
  assign array_update_85031[8] = add_84176 == 32'h0000_0008 ? array_update_85029 : array_update_85018[8];
  assign array_update_85031[9] = add_84176 == 32'h0000_0009 ? array_update_85029 : array_update_85018[9];
  assign array_index_85033 = array_update_72021[add_85030 > 32'h0000_0009 ? 4'h9 : add_85030[3:0]];
  assign array_index_85034 = array_update_85031[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_85038 = smul32b_32b_x_32b(array_index_84183[add_85030 > 32'h0000_0009 ? 4'h9 : add_85030[3:0]], array_index_85033[add_84989 > 32'h0000_0009 ? 4'h9 : add_84989[3:0]]);
  assign add_85040 = array_index_85034[add_84989 > 32'h0000_0009 ? 4'h9 : add_84989[3:0]] + smul_85038;
  assign array_update_85042[0] = add_84989 == 32'h0000_0000 ? add_85040 : array_index_85034[0];
  assign array_update_85042[1] = add_84989 == 32'h0000_0001 ? add_85040 : array_index_85034[1];
  assign array_update_85042[2] = add_84989 == 32'h0000_0002 ? add_85040 : array_index_85034[2];
  assign array_update_85042[3] = add_84989 == 32'h0000_0003 ? add_85040 : array_index_85034[3];
  assign array_update_85042[4] = add_84989 == 32'h0000_0004 ? add_85040 : array_index_85034[4];
  assign array_update_85042[5] = add_84989 == 32'h0000_0005 ? add_85040 : array_index_85034[5];
  assign array_update_85042[6] = add_84989 == 32'h0000_0006 ? add_85040 : array_index_85034[6];
  assign array_update_85042[7] = add_84989 == 32'h0000_0007 ? add_85040 : array_index_85034[7];
  assign array_update_85042[8] = add_84989 == 32'h0000_0008 ? add_85040 : array_index_85034[8];
  assign array_update_85042[9] = add_84989 == 32'h0000_0009 ? add_85040 : array_index_85034[9];
  assign add_85043 = add_85030 + 32'h0000_0001;
  assign array_update_85044[0] = add_84176 == 32'h0000_0000 ? array_update_85042 : array_update_85031[0];
  assign array_update_85044[1] = add_84176 == 32'h0000_0001 ? array_update_85042 : array_update_85031[1];
  assign array_update_85044[2] = add_84176 == 32'h0000_0002 ? array_update_85042 : array_update_85031[2];
  assign array_update_85044[3] = add_84176 == 32'h0000_0003 ? array_update_85042 : array_update_85031[3];
  assign array_update_85044[4] = add_84176 == 32'h0000_0004 ? array_update_85042 : array_update_85031[4];
  assign array_update_85044[5] = add_84176 == 32'h0000_0005 ? array_update_85042 : array_update_85031[5];
  assign array_update_85044[6] = add_84176 == 32'h0000_0006 ? array_update_85042 : array_update_85031[6];
  assign array_update_85044[7] = add_84176 == 32'h0000_0007 ? array_update_85042 : array_update_85031[7];
  assign array_update_85044[8] = add_84176 == 32'h0000_0008 ? array_update_85042 : array_update_85031[8];
  assign array_update_85044[9] = add_84176 == 32'h0000_0009 ? array_update_85042 : array_update_85031[9];
  assign array_index_85046 = array_update_72021[add_85043 > 32'h0000_0009 ? 4'h9 : add_85043[3:0]];
  assign array_index_85047 = array_update_85044[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_85051 = smul32b_32b_x_32b(array_index_84183[add_85043 > 32'h0000_0009 ? 4'h9 : add_85043[3:0]], array_index_85046[add_84989 > 32'h0000_0009 ? 4'h9 : add_84989[3:0]]);
  assign add_85053 = array_index_85047[add_84989 > 32'h0000_0009 ? 4'h9 : add_84989[3:0]] + smul_85051;
  assign array_update_85055[0] = add_84989 == 32'h0000_0000 ? add_85053 : array_index_85047[0];
  assign array_update_85055[1] = add_84989 == 32'h0000_0001 ? add_85053 : array_index_85047[1];
  assign array_update_85055[2] = add_84989 == 32'h0000_0002 ? add_85053 : array_index_85047[2];
  assign array_update_85055[3] = add_84989 == 32'h0000_0003 ? add_85053 : array_index_85047[3];
  assign array_update_85055[4] = add_84989 == 32'h0000_0004 ? add_85053 : array_index_85047[4];
  assign array_update_85055[5] = add_84989 == 32'h0000_0005 ? add_85053 : array_index_85047[5];
  assign array_update_85055[6] = add_84989 == 32'h0000_0006 ? add_85053 : array_index_85047[6];
  assign array_update_85055[7] = add_84989 == 32'h0000_0007 ? add_85053 : array_index_85047[7];
  assign array_update_85055[8] = add_84989 == 32'h0000_0008 ? add_85053 : array_index_85047[8];
  assign array_update_85055[9] = add_84989 == 32'h0000_0009 ? add_85053 : array_index_85047[9];
  assign add_85056 = add_85043 + 32'h0000_0001;
  assign array_update_85057[0] = add_84176 == 32'h0000_0000 ? array_update_85055 : array_update_85044[0];
  assign array_update_85057[1] = add_84176 == 32'h0000_0001 ? array_update_85055 : array_update_85044[1];
  assign array_update_85057[2] = add_84176 == 32'h0000_0002 ? array_update_85055 : array_update_85044[2];
  assign array_update_85057[3] = add_84176 == 32'h0000_0003 ? array_update_85055 : array_update_85044[3];
  assign array_update_85057[4] = add_84176 == 32'h0000_0004 ? array_update_85055 : array_update_85044[4];
  assign array_update_85057[5] = add_84176 == 32'h0000_0005 ? array_update_85055 : array_update_85044[5];
  assign array_update_85057[6] = add_84176 == 32'h0000_0006 ? array_update_85055 : array_update_85044[6];
  assign array_update_85057[7] = add_84176 == 32'h0000_0007 ? array_update_85055 : array_update_85044[7];
  assign array_update_85057[8] = add_84176 == 32'h0000_0008 ? array_update_85055 : array_update_85044[8];
  assign array_update_85057[9] = add_84176 == 32'h0000_0009 ? array_update_85055 : array_update_85044[9];
  assign array_index_85059 = array_update_72021[add_85056 > 32'h0000_0009 ? 4'h9 : add_85056[3:0]];
  assign array_index_85060 = array_update_85057[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_85064 = smul32b_32b_x_32b(array_index_84183[add_85056 > 32'h0000_0009 ? 4'h9 : add_85056[3:0]], array_index_85059[add_84989 > 32'h0000_0009 ? 4'h9 : add_84989[3:0]]);
  assign add_85066 = array_index_85060[add_84989 > 32'h0000_0009 ? 4'h9 : add_84989[3:0]] + smul_85064;
  assign array_update_85068[0] = add_84989 == 32'h0000_0000 ? add_85066 : array_index_85060[0];
  assign array_update_85068[1] = add_84989 == 32'h0000_0001 ? add_85066 : array_index_85060[1];
  assign array_update_85068[2] = add_84989 == 32'h0000_0002 ? add_85066 : array_index_85060[2];
  assign array_update_85068[3] = add_84989 == 32'h0000_0003 ? add_85066 : array_index_85060[3];
  assign array_update_85068[4] = add_84989 == 32'h0000_0004 ? add_85066 : array_index_85060[4];
  assign array_update_85068[5] = add_84989 == 32'h0000_0005 ? add_85066 : array_index_85060[5];
  assign array_update_85068[6] = add_84989 == 32'h0000_0006 ? add_85066 : array_index_85060[6];
  assign array_update_85068[7] = add_84989 == 32'h0000_0007 ? add_85066 : array_index_85060[7];
  assign array_update_85068[8] = add_84989 == 32'h0000_0008 ? add_85066 : array_index_85060[8];
  assign array_update_85068[9] = add_84989 == 32'h0000_0009 ? add_85066 : array_index_85060[9];
  assign add_85069 = add_85056 + 32'h0000_0001;
  assign array_update_85070[0] = add_84176 == 32'h0000_0000 ? array_update_85068 : array_update_85057[0];
  assign array_update_85070[1] = add_84176 == 32'h0000_0001 ? array_update_85068 : array_update_85057[1];
  assign array_update_85070[2] = add_84176 == 32'h0000_0002 ? array_update_85068 : array_update_85057[2];
  assign array_update_85070[3] = add_84176 == 32'h0000_0003 ? array_update_85068 : array_update_85057[3];
  assign array_update_85070[4] = add_84176 == 32'h0000_0004 ? array_update_85068 : array_update_85057[4];
  assign array_update_85070[5] = add_84176 == 32'h0000_0005 ? array_update_85068 : array_update_85057[5];
  assign array_update_85070[6] = add_84176 == 32'h0000_0006 ? array_update_85068 : array_update_85057[6];
  assign array_update_85070[7] = add_84176 == 32'h0000_0007 ? array_update_85068 : array_update_85057[7];
  assign array_update_85070[8] = add_84176 == 32'h0000_0008 ? array_update_85068 : array_update_85057[8];
  assign array_update_85070[9] = add_84176 == 32'h0000_0009 ? array_update_85068 : array_update_85057[9];
  assign array_index_85072 = array_update_72021[add_85069 > 32'h0000_0009 ? 4'h9 : add_85069[3:0]];
  assign array_index_85073 = array_update_85070[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_85077 = smul32b_32b_x_32b(array_index_84183[add_85069 > 32'h0000_0009 ? 4'h9 : add_85069[3:0]], array_index_85072[add_84989 > 32'h0000_0009 ? 4'h9 : add_84989[3:0]]);
  assign add_85079 = array_index_85073[add_84989 > 32'h0000_0009 ? 4'h9 : add_84989[3:0]] + smul_85077;
  assign array_update_85081[0] = add_84989 == 32'h0000_0000 ? add_85079 : array_index_85073[0];
  assign array_update_85081[1] = add_84989 == 32'h0000_0001 ? add_85079 : array_index_85073[1];
  assign array_update_85081[2] = add_84989 == 32'h0000_0002 ? add_85079 : array_index_85073[2];
  assign array_update_85081[3] = add_84989 == 32'h0000_0003 ? add_85079 : array_index_85073[3];
  assign array_update_85081[4] = add_84989 == 32'h0000_0004 ? add_85079 : array_index_85073[4];
  assign array_update_85081[5] = add_84989 == 32'h0000_0005 ? add_85079 : array_index_85073[5];
  assign array_update_85081[6] = add_84989 == 32'h0000_0006 ? add_85079 : array_index_85073[6];
  assign array_update_85081[7] = add_84989 == 32'h0000_0007 ? add_85079 : array_index_85073[7];
  assign array_update_85081[8] = add_84989 == 32'h0000_0008 ? add_85079 : array_index_85073[8];
  assign array_update_85081[9] = add_84989 == 32'h0000_0009 ? add_85079 : array_index_85073[9];
  assign add_85082 = add_85069 + 32'h0000_0001;
  assign array_update_85083[0] = add_84176 == 32'h0000_0000 ? array_update_85081 : array_update_85070[0];
  assign array_update_85083[1] = add_84176 == 32'h0000_0001 ? array_update_85081 : array_update_85070[1];
  assign array_update_85083[2] = add_84176 == 32'h0000_0002 ? array_update_85081 : array_update_85070[2];
  assign array_update_85083[3] = add_84176 == 32'h0000_0003 ? array_update_85081 : array_update_85070[3];
  assign array_update_85083[4] = add_84176 == 32'h0000_0004 ? array_update_85081 : array_update_85070[4];
  assign array_update_85083[5] = add_84176 == 32'h0000_0005 ? array_update_85081 : array_update_85070[5];
  assign array_update_85083[6] = add_84176 == 32'h0000_0006 ? array_update_85081 : array_update_85070[6];
  assign array_update_85083[7] = add_84176 == 32'h0000_0007 ? array_update_85081 : array_update_85070[7];
  assign array_update_85083[8] = add_84176 == 32'h0000_0008 ? array_update_85081 : array_update_85070[8];
  assign array_update_85083[9] = add_84176 == 32'h0000_0009 ? array_update_85081 : array_update_85070[9];
  assign array_index_85085 = array_update_72021[add_85082 > 32'h0000_0009 ? 4'h9 : add_85082[3:0]];
  assign array_index_85086 = array_update_85083[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_85090 = smul32b_32b_x_32b(array_index_84183[add_85082 > 32'h0000_0009 ? 4'h9 : add_85082[3:0]], array_index_85085[add_84989 > 32'h0000_0009 ? 4'h9 : add_84989[3:0]]);
  assign add_85092 = array_index_85086[add_84989 > 32'h0000_0009 ? 4'h9 : add_84989[3:0]] + smul_85090;
  assign array_update_85094[0] = add_84989 == 32'h0000_0000 ? add_85092 : array_index_85086[0];
  assign array_update_85094[1] = add_84989 == 32'h0000_0001 ? add_85092 : array_index_85086[1];
  assign array_update_85094[2] = add_84989 == 32'h0000_0002 ? add_85092 : array_index_85086[2];
  assign array_update_85094[3] = add_84989 == 32'h0000_0003 ? add_85092 : array_index_85086[3];
  assign array_update_85094[4] = add_84989 == 32'h0000_0004 ? add_85092 : array_index_85086[4];
  assign array_update_85094[5] = add_84989 == 32'h0000_0005 ? add_85092 : array_index_85086[5];
  assign array_update_85094[6] = add_84989 == 32'h0000_0006 ? add_85092 : array_index_85086[6];
  assign array_update_85094[7] = add_84989 == 32'h0000_0007 ? add_85092 : array_index_85086[7];
  assign array_update_85094[8] = add_84989 == 32'h0000_0008 ? add_85092 : array_index_85086[8];
  assign array_update_85094[9] = add_84989 == 32'h0000_0009 ? add_85092 : array_index_85086[9];
  assign add_85095 = add_85082 + 32'h0000_0001;
  assign array_update_85096[0] = add_84176 == 32'h0000_0000 ? array_update_85094 : array_update_85083[0];
  assign array_update_85096[1] = add_84176 == 32'h0000_0001 ? array_update_85094 : array_update_85083[1];
  assign array_update_85096[2] = add_84176 == 32'h0000_0002 ? array_update_85094 : array_update_85083[2];
  assign array_update_85096[3] = add_84176 == 32'h0000_0003 ? array_update_85094 : array_update_85083[3];
  assign array_update_85096[4] = add_84176 == 32'h0000_0004 ? array_update_85094 : array_update_85083[4];
  assign array_update_85096[5] = add_84176 == 32'h0000_0005 ? array_update_85094 : array_update_85083[5];
  assign array_update_85096[6] = add_84176 == 32'h0000_0006 ? array_update_85094 : array_update_85083[6];
  assign array_update_85096[7] = add_84176 == 32'h0000_0007 ? array_update_85094 : array_update_85083[7];
  assign array_update_85096[8] = add_84176 == 32'h0000_0008 ? array_update_85094 : array_update_85083[8];
  assign array_update_85096[9] = add_84176 == 32'h0000_0009 ? array_update_85094 : array_update_85083[9];
  assign array_index_85098 = array_update_72021[add_85095 > 32'h0000_0009 ? 4'h9 : add_85095[3:0]];
  assign array_index_85099 = array_update_85096[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_85103 = smul32b_32b_x_32b(array_index_84183[add_85095 > 32'h0000_0009 ? 4'h9 : add_85095[3:0]], array_index_85098[add_84989 > 32'h0000_0009 ? 4'h9 : add_84989[3:0]]);
  assign add_85105 = array_index_85099[add_84989 > 32'h0000_0009 ? 4'h9 : add_84989[3:0]] + smul_85103;
  assign array_update_85107[0] = add_84989 == 32'h0000_0000 ? add_85105 : array_index_85099[0];
  assign array_update_85107[1] = add_84989 == 32'h0000_0001 ? add_85105 : array_index_85099[1];
  assign array_update_85107[2] = add_84989 == 32'h0000_0002 ? add_85105 : array_index_85099[2];
  assign array_update_85107[3] = add_84989 == 32'h0000_0003 ? add_85105 : array_index_85099[3];
  assign array_update_85107[4] = add_84989 == 32'h0000_0004 ? add_85105 : array_index_85099[4];
  assign array_update_85107[5] = add_84989 == 32'h0000_0005 ? add_85105 : array_index_85099[5];
  assign array_update_85107[6] = add_84989 == 32'h0000_0006 ? add_85105 : array_index_85099[6];
  assign array_update_85107[7] = add_84989 == 32'h0000_0007 ? add_85105 : array_index_85099[7];
  assign array_update_85107[8] = add_84989 == 32'h0000_0008 ? add_85105 : array_index_85099[8];
  assign array_update_85107[9] = add_84989 == 32'h0000_0009 ? add_85105 : array_index_85099[9];
  assign add_85108 = add_85095 + 32'h0000_0001;
  assign array_update_85109[0] = add_84176 == 32'h0000_0000 ? array_update_85107 : array_update_85096[0];
  assign array_update_85109[1] = add_84176 == 32'h0000_0001 ? array_update_85107 : array_update_85096[1];
  assign array_update_85109[2] = add_84176 == 32'h0000_0002 ? array_update_85107 : array_update_85096[2];
  assign array_update_85109[3] = add_84176 == 32'h0000_0003 ? array_update_85107 : array_update_85096[3];
  assign array_update_85109[4] = add_84176 == 32'h0000_0004 ? array_update_85107 : array_update_85096[4];
  assign array_update_85109[5] = add_84176 == 32'h0000_0005 ? array_update_85107 : array_update_85096[5];
  assign array_update_85109[6] = add_84176 == 32'h0000_0006 ? array_update_85107 : array_update_85096[6];
  assign array_update_85109[7] = add_84176 == 32'h0000_0007 ? array_update_85107 : array_update_85096[7];
  assign array_update_85109[8] = add_84176 == 32'h0000_0008 ? array_update_85107 : array_update_85096[8];
  assign array_update_85109[9] = add_84176 == 32'h0000_0009 ? array_update_85107 : array_update_85096[9];
  assign array_index_85111 = array_update_72021[add_85108 > 32'h0000_0009 ? 4'h9 : add_85108[3:0]];
  assign array_index_85112 = array_update_85109[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_85116 = smul32b_32b_x_32b(array_index_84183[add_85108 > 32'h0000_0009 ? 4'h9 : add_85108[3:0]], array_index_85111[add_84989 > 32'h0000_0009 ? 4'h9 : add_84989[3:0]]);
  assign add_85118 = array_index_85112[add_84989 > 32'h0000_0009 ? 4'h9 : add_84989[3:0]] + smul_85116;
  assign array_update_85119[0] = add_84989 == 32'h0000_0000 ? add_85118 : array_index_85112[0];
  assign array_update_85119[1] = add_84989 == 32'h0000_0001 ? add_85118 : array_index_85112[1];
  assign array_update_85119[2] = add_84989 == 32'h0000_0002 ? add_85118 : array_index_85112[2];
  assign array_update_85119[3] = add_84989 == 32'h0000_0003 ? add_85118 : array_index_85112[3];
  assign array_update_85119[4] = add_84989 == 32'h0000_0004 ? add_85118 : array_index_85112[4];
  assign array_update_85119[5] = add_84989 == 32'h0000_0005 ? add_85118 : array_index_85112[5];
  assign array_update_85119[6] = add_84989 == 32'h0000_0006 ? add_85118 : array_index_85112[6];
  assign array_update_85119[7] = add_84989 == 32'h0000_0007 ? add_85118 : array_index_85112[7];
  assign array_update_85119[8] = add_84989 == 32'h0000_0008 ? add_85118 : array_index_85112[8];
  assign array_update_85119[9] = add_84989 == 32'h0000_0009 ? add_85118 : array_index_85112[9];
  assign array_update_85120[0] = add_84176 == 32'h0000_0000 ? array_update_85119 : array_update_85109[0];
  assign array_update_85120[1] = add_84176 == 32'h0000_0001 ? array_update_85119 : array_update_85109[1];
  assign array_update_85120[2] = add_84176 == 32'h0000_0002 ? array_update_85119 : array_update_85109[2];
  assign array_update_85120[3] = add_84176 == 32'h0000_0003 ? array_update_85119 : array_update_85109[3];
  assign array_update_85120[4] = add_84176 == 32'h0000_0004 ? array_update_85119 : array_update_85109[4];
  assign array_update_85120[5] = add_84176 == 32'h0000_0005 ? array_update_85119 : array_update_85109[5];
  assign array_update_85120[6] = add_84176 == 32'h0000_0006 ? array_update_85119 : array_update_85109[6];
  assign array_update_85120[7] = add_84176 == 32'h0000_0007 ? array_update_85119 : array_update_85109[7];
  assign array_update_85120[8] = add_84176 == 32'h0000_0008 ? array_update_85119 : array_update_85109[8];
  assign array_update_85120[9] = add_84176 == 32'h0000_0009 ? array_update_85119 : array_update_85109[9];
  assign array_index_85122 = array_update_85120[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign add_85124 = add_84989 + 32'h0000_0001;
  assign array_update_85125[0] = add_85124 == 32'h0000_0000 ? 32'h0000_0000 : array_index_85122[0];
  assign array_update_85125[1] = add_85124 == 32'h0000_0001 ? 32'h0000_0000 : array_index_85122[1];
  assign array_update_85125[2] = add_85124 == 32'h0000_0002 ? 32'h0000_0000 : array_index_85122[2];
  assign array_update_85125[3] = add_85124 == 32'h0000_0003 ? 32'h0000_0000 : array_index_85122[3];
  assign array_update_85125[4] = add_85124 == 32'h0000_0004 ? 32'h0000_0000 : array_index_85122[4];
  assign array_update_85125[5] = add_85124 == 32'h0000_0005 ? 32'h0000_0000 : array_index_85122[5];
  assign array_update_85125[6] = add_85124 == 32'h0000_0006 ? 32'h0000_0000 : array_index_85122[6];
  assign array_update_85125[7] = add_85124 == 32'h0000_0007 ? 32'h0000_0000 : array_index_85122[7];
  assign array_update_85125[8] = add_85124 == 32'h0000_0008 ? 32'h0000_0000 : array_index_85122[8];
  assign array_update_85125[9] = add_85124 == 32'h0000_0009 ? 32'h0000_0000 : array_index_85122[9];
  assign literal_85126 = 32'h0000_0000;
  assign array_update_85127[0] = add_84176 == 32'h0000_0000 ? array_update_85125 : array_update_85120[0];
  assign array_update_85127[1] = add_84176 == 32'h0000_0001 ? array_update_85125 : array_update_85120[1];
  assign array_update_85127[2] = add_84176 == 32'h0000_0002 ? array_update_85125 : array_update_85120[2];
  assign array_update_85127[3] = add_84176 == 32'h0000_0003 ? array_update_85125 : array_update_85120[3];
  assign array_update_85127[4] = add_84176 == 32'h0000_0004 ? array_update_85125 : array_update_85120[4];
  assign array_update_85127[5] = add_84176 == 32'h0000_0005 ? array_update_85125 : array_update_85120[5];
  assign array_update_85127[6] = add_84176 == 32'h0000_0006 ? array_update_85125 : array_update_85120[6];
  assign array_update_85127[7] = add_84176 == 32'h0000_0007 ? array_update_85125 : array_update_85120[7];
  assign array_update_85127[8] = add_84176 == 32'h0000_0008 ? array_update_85125 : array_update_85120[8];
  assign array_update_85127[9] = add_84176 == 32'h0000_0009 ? array_update_85125 : array_update_85120[9];
  assign array_index_85129 = array_update_72021[literal_85126 > 32'h0000_0009 ? 4'h9 : literal_85126[3:0]];
  assign array_index_85130 = array_update_85127[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_85134 = smul32b_32b_x_32b(array_index_84183[literal_85126 > 32'h0000_0009 ? 4'h9 : literal_85126[3:0]], array_index_85129[add_85124 > 32'h0000_0009 ? 4'h9 : add_85124[3:0]]);
  assign add_85136 = array_index_85130[add_85124 > 32'h0000_0009 ? 4'h9 : add_85124[3:0]] + smul_85134;
  assign array_update_85138[0] = add_85124 == 32'h0000_0000 ? add_85136 : array_index_85130[0];
  assign array_update_85138[1] = add_85124 == 32'h0000_0001 ? add_85136 : array_index_85130[1];
  assign array_update_85138[2] = add_85124 == 32'h0000_0002 ? add_85136 : array_index_85130[2];
  assign array_update_85138[3] = add_85124 == 32'h0000_0003 ? add_85136 : array_index_85130[3];
  assign array_update_85138[4] = add_85124 == 32'h0000_0004 ? add_85136 : array_index_85130[4];
  assign array_update_85138[5] = add_85124 == 32'h0000_0005 ? add_85136 : array_index_85130[5];
  assign array_update_85138[6] = add_85124 == 32'h0000_0006 ? add_85136 : array_index_85130[6];
  assign array_update_85138[7] = add_85124 == 32'h0000_0007 ? add_85136 : array_index_85130[7];
  assign array_update_85138[8] = add_85124 == 32'h0000_0008 ? add_85136 : array_index_85130[8];
  assign array_update_85138[9] = add_85124 == 32'h0000_0009 ? add_85136 : array_index_85130[9];
  assign add_85139 = literal_85126 + 32'h0000_0001;
  assign array_update_85140[0] = add_84176 == 32'h0000_0000 ? array_update_85138 : array_update_85127[0];
  assign array_update_85140[1] = add_84176 == 32'h0000_0001 ? array_update_85138 : array_update_85127[1];
  assign array_update_85140[2] = add_84176 == 32'h0000_0002 ? array_update_85138 : array_update_85127[2];
  assign array_update_85140[3] = add_84176 == 32'h0000_0003 ? array_update_85138 : array_update_85127[3];
  assign array_update_85140[4] = add_84176 == 32'h0000_0004 ? array_update_85138 : array_update_85127[4];
  assign array_update_85140[5] = add_84176 == 32'h0000_0005 ? array_update_85138 : array_update_85127[5];
  assign array_update_85140[6] = add_84176 == 32'h0000_0006 ? array_update_85138 : array_update_85127[6];
  assign array_update_85140[7] = add_84176 == 32'h0000_0007 ? array_update_85138 : array_update_85127[7];
  assign array_update_85140[8] = add_84176 == 32'h0000_0008 ? array_update_85138 : array_update_85127[8];
  assign array_update_85140[9] = add_84176 == 32'h0000_0009 ? array_update_85138 : array_update_85127[9];
  assign array_index_85142 = array_update_72021[add_85139 > 32'h0000_0009 ? 4'h9 : add_85139[3:0]];
  assign array_index_85143 = array_update_85140[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_85147 = smul32b_32b_x_32b(array_index_84183[add_85139 > 32'h0000_0009 ? 4'h9 : add_85139[3:0]], array_index_85142[add_85124 > 32'h0000_0009 ? 4'h9 : add_85124[3:0]]);
  assign add_85149 = array_index_85143[add_85124 > 32'h0000_0009 ? 4'h9 : add_85124[3:0]] + smul_85147;
  assign array_update_85151[0] = add_85124 == 32'h0000_0000 ? add_85149 : array_index_85143[0];
  assign array_update_85151[1] = add_85124 == 32'h0000_0001 ? add_85149 : array_index_85143[1];
  assign array_update_85151[2] = add_85124 == 32'h0000_0002 ? add_85149 : array_index_85143[2];
  assign array_update_85151[3] = add_85124 == 32'h0000_0003 ? add_85149 : array_index_85143[3];
  assign array_update_85151[4] = add_85124 == 32'h0000_0004 ? add_85149 : array_index_85143[4];
  assign array_update_85151[5] = add_85124 == 32'h0000_0005 ? add_85149 : array_index_85143[5];
  assign array_update_85151[6] = add_85124 == 32'h0000_0006 ? add_85149 : array_index_85143[6];
  assign array_update_85151[7] = add_85124 == 32'h0000_0007 ? add_85149 : array_index_85143[7];
  assign array_update_85151[8] = add_85124 == 32'h0000_0008 ? add_85149 : array_index_85143[8];
  assign array_update_85151[9] = add_85124 == 32'h0000_0009 ? add_85149 : array_index_85143[9];
  assign add_85152 = add_85139 + 32'h0000_0001;
  assign array_update_85153[0] = add_84176 == 32'h0000_0000 ? array_update_85151 : array_update_85140[0];
  assign array_update_85153[1] = add_84176 == 32'h0000_0001 ? array_update_85151 : array_update_85140[1];
  assign array_update_85153[2] = add_84176 == 32'h0000_0002 ? array_update_85151 : array_update_85140[2];
  assign array_update_85153[3] = add_84176 == 32'h0000_0003 ? array_update_85151 : array_update_85140[3];
  assign array_update_85153[4] = add_84176 == 32'h0000_0004 ? array_update_85151 : array_update_85140[4];
  assign array_update_85153[5] = add_84176 == 32'h0000_0005 ? array_update_85151 : array_update_85140[5];
  assign array_update_85153[6] = add_84176 == 32'h0000_0006 ? array_update_85151 : array_update_85140[6];
  assign array_update_85153[7] = add_84176 == 32'h0000_0007 ? array_update_85151 : array_update_85140[7];
  assign array_update_85153[8] = add_84176 == 32'h0000_0008 ? array_update_85151 : array_update_85140[8];
  assign array_update_85153[9] = add_84176 == 32'h0000_0009 ? array_update_85151 : array_update_85140[9];
  assign array_index_85155 = array_update_72021[add_85152 > 32'h0000_0009 ? 4'h9 : add_85152[3:0]];
  assign array_index_85156 = array_update_85153[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_85160 = smul32b_32b_x_32b(array_index_84183[add_85152 > 32'h0000_0009 ? 4'h9 : add_85152[3:0]], array_index_85155[add_85124 > 32'h0000_0009 ? 4'h9 : add_85124[3:0]]);
  assign add_85162 = array_index_85156[add_85124 > 32'h0000_0009 ? 4'h9 : add_85124[3:0]] + smul_85160;
  assign array_update_85164[0] = add_85124 == 32'h0000_0000 ? add_85162 : array_index_85156[0];
  assign array_update_85164[1] = add_85124 == 32'h0000_0001 ? add_85162 : array_index_85156[1];
  assign array_update_85164[2] = add_85124 == 32'h0000_0002 ? add_85162 : array_index_85156[2];
  assign array_update_85164[3] = add_85124 == 32'h0000_0003 ? add_85162 : array_index_85156[3];
  assign array_update_85164[4] = add_85124 == 32'h0000_0004 ? add_85162 : array_index_85156[4];
  assign array_update_85164[5] = add_85124 == 32'h0000_0005 ? add_85162 : array_index_85156[5];
  assign array_update_85164[6] = add_85124 == 32'h0000_0006 ? add_85162 : array_index_85156[6];
  assign array_update_85164[7] = add_85124 == 32'h0000_0007 ? add_85162 : array_index_85156[7];
  assign array_update_85164[8] = add_85124 == 32'h0000_0008 ? add_85162 : array_index_85156[8];
  assign array_update_85164[9] = add_85124 == 32'h0000_0009 ? add_85162 : array_index_85156[9];
  assign add_85165 = add_85152 + 32'h0000_0001;
  assign array_update_85166[0] = add_84176 == 32'h0000_0000 ? array_update_85164 : array_update_85153[0];
  assign array_update_85166[1] = add_84176 == 32'h0000_0001 ? array_update_85164 : array_update_85153[1];
  assign array_update_85166[2] = add_84176 == 32'h0000_0002 ? array_update_85164 : array_update_85153[2];
  assign array_update_85166[3] = add_84176 == 32'h0000_0003 ? array_update_85164 : array_update_85153[3];
  assign array_update_85166[4] = add_84176 == 32'h0000_0004 ? array_update_85164 : array_update_85153[4];
  assign array_update_85166[5] = add_84176 == 32'h0000_0005 ? array_update_85164 : array_update_85153[5];
  assign array_update_85166[6] = add_84176 == 32'h0000_0006 ? array_update_85164 : array_update_85153[6];
  assign array_update_85166[7] = add_84176 == 32'h0000_0007 ? array_update_85164 : array_update_85153[7];
  assign array_update_85166[8] = add_84176 == 32'h0000_0008 ? array_update_85164 : array_update_85153[8];
  assign array_update_85166[9] = add_84176 == 32'h0000_0009 ? array_update_85164 : array_update_85153[9];
  assign array_index_85168 = array_update_72021[add_85165 > 32'h0000_0009 ? 4'h9 : add_85165[3:0]];
  assign array_index_85169 = array_update_85166[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_85173 = smul32b_32b_x_32b(array_index_84183[add_85165 > 32'h0000_0009 ? 4'h9 : add_85165[3:0]], array_index_85168[add_85124 > 32'h0000_0009 ? 4'h9 : add_85124[3:0]]);
  assign add_85175 = array_index_85169[add_85124 > 32'h0000_0009 ? 4'h9 : add_85124[3:0]] + smul_85173;
  assign array_update_85177[0] = add_85124 == 32'h0000_0000 ? add_85175 : array_index_85169[0];
  assign array_update_85177[1] = add_85124 == 32'h0000_0001 ? add_85175 : array_index_85169[1];
  assign array_update_85177[2] = add_85124 == 32'h0000_0002 ? add_85175 : array_index_85169[2];
  assign array_update_85177[3] = add_85124 == 32'h0000_0003 ? add_85175 : array_index_85169[3];
  assign array_update_85177[4] = add_85124 == 32'h0000_0004 ? add_85175 : array_index_85169[4];
  assign array_update_85177[5] = add_85124 == 32'h0000_0005 ? add_85175 : array_index_85169[5];
  assign array_update_85177[6] = add_85124 == 32'h0000_0006 ? add_85175 : array_index_85169[6];
  assign array_update_85177[7] = add_85124 == 32'h0000_0007 ? add_85175 : array_index_85169[7];
  assign array_update_85177[8] = add_85124 == 32'h0000_0008 ? add_85175 : array_index_85169[8];
  assign array_update_85177[9] = add_85124 == 32'h0000_0009 ? add_85175 : array_index_85169[9];
  assign add_85178 = add_85165 + 32'h0000_0001;
  assign array_update_85179[0] = add_84176 == 32'h0000_0000 ? array_update_85177 : array_update_85166[0];
  assign array_update_85179[1] = add_84176 == 32'h0000_0001 ? array_update_85177 : array_update_85166[1];
  assign array_update_85179[2] = add_84176 == 32'h0000_0002 ? array_update_85177 : array_update_85166[2];
  assign array_update_85179[3] = add_84176 == 32'h0000_0003 ? array_update_85177 : array_update_85166[3];
  assign array_update_85179[4] = add_84176 == 32'h0000_0004 ? array_update_85177 : array_update_85166[4];
  assign array_update_85179[5] = add_84176 == 32'h0000_0005 ? array_update_85177 : array_update_85166[5];
  assign array_update_85179[6] = add_84176 == 32'h0000_0006 ? array_update_85177 : array_update_85166[6];
  assign array_update_85179[7] = add_84176 == 32'h0000_0007 ? array_update_85177 : array_update_85166[7];
  assign array_update_85179[8] = add_84176 == 32'h0000_0008 ? array_update_85177 : array_update_85166[8];
  assign array_update_85179[9] = add_84176 == 32'h0000_0009 ? array_update_85177 : array_update_85166[9];
  assign array_index_85181 = array_update_72021[add_85178 > 32'h0000_0009 ? 4'h9 : add_85178[3:0]];
  assign array_index_85182 = array_update_85179[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_85186 = smul32b_32b_x_32b(array_index_84183[add_85178 > 32'h0000_0009 ? 4'h9 : add_85178[3:0]], array_index_85181[add_85124 > 32'h0000_0009 ? 4'h9 : add_85124[3:0]]);
  assign add_85188 = array_index_85182[add_85124 > 32'h0000_0009 ? 4'h9 : add_85124[3:0]] + smul_85186;
  assign array_update_85190[0] = add_85124 == 32'h0000_0000 ? add_85188 : array_index_85182[0];
  assign array_update_85190[1] = add_85124 == 32'h0000_0001 ? add_85188 : array_index_85182[1];
  assign array_update_85190[2] = add_85124 == 32'h0000_0002 ? add_85188 : array_index_85182[2];
  assign array_update_85190[3] = add_85124 == 32'h0000_0003 ? add_85188 : array_index_85182[3];
  assign array_update_85190[4] = add_85124 == 32'h0000_0004 ? add_85188 : array_index_85182[4];
  assign array_update_85190[5] = add_85124 == 32'h0000_0005 ? add_85188 : array_index_85182[5];
  assign array_update_85190[6] = add_85124 == 32'h0000_0006 ? add_85188 : array_index_85182[6];
  assign array_update_85190[7] = add_85124 == 32'h0000_0007 ? add_85188 : array_index_85182[7];
  assign array_update_85190[8] = add_85124 == 32'h0000_0008 ? add_85188 : array_index_85182[8];
  assign array_update_85190[9] = add_85124 == 32'h0000_0009 ? add_85188 : array_index_85182[9];
  assign add_85191 = add_85178 + 32'h0000_0001;
  assign array_update_85192[0] = add_84176 == 32'h0000_0000 ? array_update_85190 : array_update_85179[0];
  assign array_update_85192[1] = add_84176 == 32'h0000_0001 ? array_update_85190 : array_update_85179[1];
  assign array_update_85192[2] = add_84176 == 32'h0000_0002 ? array_update_85190 : array_update_85179[2];
  assign array_update_85192[3] = add_84176 == 32'h0000_0003 ? array_update_85190 : array_update_85179[3];
  assign array_update_85192[4] = add_84176 == 32'h0000_0004 ? array_update_85190 : array_update_85179[4];
  assign array_update_85192[5] = add_84176 == 32'h0000_0005 ? array_update_85190 : array_update_85179[5];
  assign array_update_85192[6] = add_84176 == 32'h0000_0006 ? array_update_85190 : array_update_85179[6];
  assign array_update_85192[7] = add_84176 == 32'h0000_0007 ? array_update_85190 : array_update_85179[7];
  assign array_update_85192[8] = add_84176 == 32'h0000_0008 ? array_update_85190 : array_update_85179[8];
  assign array_update_85192[9] = add_84176 == 32'h0000_0009 ? array_update_85190 : array_update_85179[9];
  assign array_index_85194 = array_update_72021[add_85191 > 32'h0000_0009 ? 4'h9 : add_85191[3:0]];
  assign array_index_85195 = array_update_85192[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_85199 = smul32b_32b_x_32b(array_index_84183[add_85191 > 32'h0000_0009 ? 4'h9 : add_85191[3:0]], array_index_85194[add_85124 > 32'h0000_0009 ? 4'h9 : add_85124[3:0]]);
  assign add_85201 = array_index_85195[add_85124 > 32'h0000_0009 ? 4'h9 : add_85124[3:0]] + smul_85199;
  assign array_update_85203[0] = add_85124 == 32'h0000_0000 ? add_85201 : array_index_85195[0];
  assign array_update_85203[1] = add_85124 == 32'h0000_0001 ? add_85201 : array_index_85195[1];
  assign array_update_85203[2] = add_85124 == 32'h0000_0002 ? add_85201 : array_index_85195[2];
  assign array_update_85203[3] = add_85124 == 32'h0000_0003 ? add_85201 : array_index_85195[3];
  assign array_update_85203[4] = add_85124 == 32'h0000_0004 ? add_85201 : array_index_85195[4];
  assign array_update_85203[5] = add_85124 == 32'h0000_0005 ? add_85201 : array_index_85195[5];
  assign array_update_85203[6] = add_85124 == 32'h0000_0006 ? add_85201 : array_index_85195[6];
  assign array_update_85203[7] = add_85124 == 32'h0000_0007 ? add_85201 : array_index_85195[7];
  assign array_update_85203[8] = add_85124 == 32'h0000_0008 ? add_85201 : array_index_85195[8];
  assign array_update_85203[9] = add_85124 == 32'h0000_0009 ? add_85201 : array_index_85195[9];
  assign add_85204 = add_85191 + 32'h0000_0001;
  assign array_update_85205[0] = add_84176 == 32'h0000_0000 ? array_update_85203 : array_update_85192[0];
  assign array_update_85205[1] = add_84176 == 32'h0000_0001 ? array_update_85203 : array_update_85192[1];
  assign array_update_85205[2] = add_84176 == 32'h0000_0002 ? array_update_85203 : array_update_85192[2];
  assign array_update_85205[3] = add_84176 == 32'h0000_0003 ? array_update_85203 : array_update_85192[3];
  assign array_update_85205[4] = add_84176 == 32'h0000_0004 ? array_update_85203 : array_update_85192[4];
  assign array_update_85205[5] = add_84176 == 32'h0000_0005 ? array_update_85203 : array_update_85192[5];
  assign array_update_85205[6] = add_84176 == 32'h0000_0006 ? array_update_85203 : array_update_85192[6];
  assign array_update_85205[7] = add_84176 == 32'h0000_0007 ? array_update_85203 : array_update_85192[7];
  assign array_update_85205[8] = add_84176 == 32'h0000_0008 ? array_update_85203 : array_update_85192[8];
  assign array_update_85205[9] = add_84176 == 32'h0000_0009 ? array_update_85203 : array_update_85192[9];
  assign array_index_85207 = array_update_72021[add_85204 > 32'h0000_0009 ? 4'h9 : add_85204[3:0]];
  assign array_index_85208 = array_update_85205[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_85212 = smul32b_32b_x_32b(array_index_84183[add_85204 > 32'h0000_0009 ? 4'h9 : add_85204[3:0]], array_index_85207[add_85124 > 32'h0000_0009 ? 4'h9 : add_85124[3:0]]);
  assign add_85214 = array_index_85208[add_85124 > 32'h0000_0009 ? 4'h9 : add_85124[3:0]] + smul_85212;
  assign array_update_85216[0] = add_85124 == 32'h0000_0000 ? add_85214 : array_index_85208[0];
  assign array_update_85216[1] = add_85124 == 32'h0000_0001 ? add_85214 : array_index_85208[1];
  assign array_update_85216[2] = add_85124 == 32'h0000_0002 ? add_85214 : array_index_85208[2];
  assign array_update_85216[3] = add_85124 == 32'h0000_0003 ? add_85214 : array_index_85208[3];
  assign array_update_85216[4] = add_85124 == 32'h0000_0004 ? add_85214 : array_index_85208[4];
  assign array_update_85216[5] = add_85124 == 32'h0000_0005 ? add_85214 : array_index_85208[5];
  assign array_update_85216[6] = add_85124 == 32'h0000_0006 ? add_85214 : array_index_85208[6];
  assign array_update_85216[7] = add_85124 == 32'h0000_0007 ? add_85214 : array_index_85208[7];
  assign array_update_85216[8] = add_85124 == 32'h0000_0008 ? add_85214 : array_index_85208[8];
  assign array_update_85216[9] = add_85124 == 32'h0000_0009 ? add_85214 : array_index_85208[9];
  assign add_85217 = add_85204 + 32'h0000_0001;
  assign array_update_85218[0] = add_84176 == 32'h0000_0000 ? array_update_85216 : array_update_85205[0];
  assign array_update_85218[1] = add_84176 == 32'h0000_0001 ? array_update_85216 : array_update_85205[1];
  assign array_update_85218[2] = add_84176 == 32'h0000_0002 ? array_update_85216 : array_update_85205[2];
  assign array_update_85218[3] = add_84176 == 32'h0000_0003 ? array_update_85216 : array_update_85205[3];
  assign array_update_85218[4] = add_84176 == 32'h0000_0004 ? array_update_85216 : array_update_85205[4];
  assign array_update_85218[5] = add_84176 == 32'h0000_0005 ? array_update_85216 : array_update_85205[5];
  assign array_update_85218[6] = add_84176 == 32'h0000_0006 ? array_update_85216 : array_update_85205[6];
  assign array_update_85218[7] = add_84176 == 32'h0000_0007 ? array_update_85216 : array_update_85205[7];
  assign array_update_85218[8] = add_84176 == 32'h0000_0008 ? array_update_85216 : array_update_85205[8];
  assign array_update_85218[9] = add_84176 == 32'h0000_0009 ? array_update_85216 : array_update_85205[9];
  assign array_index_85220 = array_update_72021[add_85217 > 32'h0000_0009 ? 4'h9 : add_85217[3:0]];
  assign array_index_85221 = array_update_85218[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_85225 = smul32b_32b_x_32b(array_index_84183[add_85217 > 32'h0000_0009 ? 4'h9 : add_85217[3:0]], array_index_85220[add_85124 > 32'h0000_0009 ? 4'h9 : add_85124[3:0]]);
  assign add_85227 = array_index_85221[add_85124 > 32'h0000_0009 ? 4'h9 : add_85124[3:0]] + smul_85225;
  assign array_update_85229[0] = add_85124 == 32'h0000_0000 ? add_85227 : array_index_85221[0];
  assign array_update_85229[1] = add_85124 == 32'h0000_0001 ? add_85227 : array_index_85221[1];
  assign array_update_85229[2] = add_85124 == 32'h0000_0002 ? add_85227 : array_index_85221[2];
  assign array_update_85229[3] = add_85124 == 32'h0000_0003 ? add_85227 : array_index_85221[3];
  assign array_update_85229[4] = add_85124 == 32'h0000_0004 ? add_85227 : array_index_85221[4];
  assign array_update_85229[5] = add_85124 == 32'h0000_0005 ? add_85227 : array_index_85221[5];
  assign array_update_85229[6] = add_85124 == 32'h0000_0006 ? add_85227 : array_index_85221[6];
  assign array_update_85229[7] = add_85124 == 32'h0000_0007 ? add_85227 : array_index_85221[7];
  assign array_update_85229[8] = add_85124 == 32'h0000_0008 ? add_85227 : array_index_85221[8];
  assign array_update_85229[9] = add_85124 == 32'h0000_0009 ? add_85227 : array_index_85221[9];
  assign add_85230 = add_85217 + 32'h0000_0001;
  assign array_update_85231[0] = add_84176 == 32'h0000_0000 ? array_update_85229 : array_update_85218[0];
  assign array_update_85231[1] = add_84176 == 32'h0000_0001 ? array_update_85229 : array_update_85218[1];
  assign array_update_85231[2] = add_84176 == 32'h0000_0002 ? array_update_85229 : array_update_85218[2];
  assign array_update_85231[3] = add_84176 == 32'h0000_0003 ? array_update_85229 : array_update_85218[3];
  assign array_update_85231[4] = add_84176 == 32'h0000_0004 ? array_update_85229 : array_update_85218[4];
  assign array_update_85231[5] = add_84176 == 32'h0000_0005 ? array_update_85229 : array_update_85218[5];
  assign array_update_85231[6] = add_84176 == 32'h0000_0006 ? array_update_85229 : array_update_85218[6];
  assign array_update_85231[7] = add_84176 == 32'h0000_0007 ? array_update_85229 : array_update_85218[7];
  assign array_update_85231[8] = add_84176 == 32'h0000_0008 ? array_update_85229 : array_update_85218[8];
  assign array_update_85231[9] = add_84176 == 32'h0000_0009 ? array_update_85229 : array_update_85218[9];
  assign array_index_85233 = array_update_72021[add_85230 > 32'h0000_0009 ? 4'h9 : add_85230[3:0]];
  assign array_index_85234 = array_update_85231[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_85238 = smul32b_32b_x_32b(array_index_84183[add_85230 > 32'h0000_0009 ? 4'h9 : add_85230[3:0]], array_index_85233[add_85124 > 32'h0000_0009 ? 4'h9 : add_85124[3:0]]);
  assign add_85240 = array_index_85234[add_85124 > 32'h0000_0009 ? 4'h9 : add_85124[3:0]] + smul_85238;
  assign array_update_85242[0] = add_85124 == 32'h0000_0000 ? add_85240 : array_index_85234[0];
  assign array_update_85242[1] = add_85124 == 32'h0000_0001 ? add_85240 : array_index_85234[1];
  assign array_update_85242[2] = add_85124 == 32'h0000_0002 ? add_85240 : array_index_85234[2];
  assign array_update_85242[3] = add_85124 == 32'h0000_0003 ? add_85240 : array_index_85234[3];
  assign array_update_85242[4] = add_85124 == 32'h0000_0004 ? add_85240 : array_index_85234[4];
  assign array_update_85242[5] = add_85124 == 32'h0000_0005 ? add_85240 : array_index_85234[5];
  assign array_update_85242[6] = add_85124 == 32'h0000_0006 ? add_85240 : array_index_85234[6];
  assign array_update_85242[7] = add_85124 == 32'h0000_0007 ? add_85240 : array_index_85234[7];
  assign array_update_85242[8] = add_85124 == 32'h0000_0008 ? add_85240 : array_index_85234[8];
  assign array_update_85242[9] = add_85124 == 32'h0000_0009 ? add_85240 : array_index_85234[9];
  assign add_85243 = add_85230 + 32'h0000_0001;
  assign array_update_85244[0] = add_84176 == 32'h0000_0000 ? array_update_85242 : array_update_85231[0];
  assign array_update_85244[1] = add_84176 == 32'h0000_0001 ? array_update_85242 : array_update_85231[1];
  assign array_update_85244[2] = add_84176 == 32'h0000_0002 ? array_update_85242 : array_update_85231[2];
  assign array_update_85244[3] = add_84176 == 32'h0000_0003 ? array_update_85242 : array_update_85231[3];
  assign array_update_85244[4] = add_84176 == 32'h0000_0004 ? array_update_85242 : array_update_85231[4];
  assign array_update_85244[5] = add_84176 == 32'h0000_0005 ? array_update_85242 : array_update_85231[5];
  assign array_update_85244[6] = add_84176 == 32'h0000_0006 ? array_update_85242 : array_update_85231[6];
  assign array_update_85244[7] = add_84176 == 32'h0000_0007 ? array_update_85242 : array_update_85231[7];
  assign array_update_85244[8] = add_84176 == 32'h0000_0008 ? array_update_85242 : array_update_85231[8];
  assign array_update_85244[9] = add_84176 == 32'h0000_0009 ? array_update_85242 : array_update_85231[9];
  assign array_index_85246 = array_update_72021[add_85243 > 32'h0000_0009 ? 4'h9 : add_85243[3:0]];
  assign array_index_85247 = array_update_85244[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_85251 = smul32b_32b_x_32b(array_index_84183[add_85243 > 32'h0000_0009 ? 4'h9 : add_85243[3:0]], array_index_85246[add_85124 > 32'h0000_0009 ? 4'h9 : add_85124[3:0]]);
  assign add_85253 = array_index_85247[add_85124 > 32'h0000_0009 ? 4'h9 : add_85124[3:0]] + smul_85251;
  assign array_update_85254[0] = add_85124 == 32'h0000_0000 ? add_85253 : array_index_85247[0];
  assign array_update_85254[1] = add_85124 == 32'h0000_0001 ? add_85253 : array_index_85247[1];
  assign array_update_85254[2] = add_85124 == 32'h0000_0002 ? add_85253 : array_index_85247[2];
  assign array_update_85254[3] = add_85124 == 32'h0000_0003 ? add_85253 : array_index_85247[3];
  assign array_update_85254[4] = add_85124 == 32'h0000_0004 ? add_85253 : array_index_85247[4];
  assign array_update_85254[5] = add_85124 == 32'h0000_0005 ? add_85253 : array_index_85247[5];
  assign array_update_85254[6] = add_85124 == 32'h0000_0006 ? add_85253 : array_index_85247[6];
  assign array_update_85254[7] = add_85124 == 32'h0000_0007 ? add_85253 : array_index_85247[7];
  assign array_update_85254[8] = add_85124 == 32'h0000_0008 ? add_85253 : array_index_85247[8];
  assign array_update_85254[9] = add_85124 == 32'h0000_0009 ? add_85253 : array_index_85247[9];
  assign array_update_85255[0] = add_84176 == 32'h0000_0000 ? array_update_85254 : array_update_85244[0];
  assign array_update_85255[1] = add_84176 == 32'h0000_0001 ? array_update_85254 : array_update_85244[1];
  assign array_update_85255[2] = add_84176 == 32'h0000_0002 ? array_update_85254 : array_update_85244[2];
  assign array_update_85255[3] = add_84176 == 32'h0000_0003 ? array_update_85254 : array_update_85244[3];
  assign array_update_85255[4] = add_84176 == 32'h0000_0004 ? array_update_85254 : array_update_85244[4];
  assign array_update_85255[5] = add_84176 == 32'h0000_0005 ? array_update_85254 : array_update_85244[5];
  assign array_update_85255[6] = add_84176 == 32'h0000_0006 ? array_update_85254 : array_update_85244[6];
  assign array_update_85255[7] = add_84176 == 32'h0000_0007 ? array_update_85254 : array_update_85244[7];
  assign array_update_85255[8] = add_84176 == 32'h0000_0008 ? array_update_85254 : array_update_85244[8];
  assign array_update_85255[9] = add_84176 == 32'h0000_0009 ? array_update_85254 : array_update_85244[9];
  assign array_index_85257 = array_update_85255[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign add_85259 = add_85124 + 32'h0000_0001;
  assign array_update_85260[0] = add_85259 == 32'h0000_0000 ? 32'h0000_0000 : array_index_85257[0];
  assign array_update_85260[1] = add_85259 == 32'h0000_0001 ? 32'h0000_0000 : array_index_85257[1];
  assign array_update_85260[2] = add_85259 == 32'h0000_0002 ? 32'h0000_0000 : array_index_85257[2];
  assign array_update_85260[3] = add_85259 == 32'h0000_0003 ? 32'h0000_0000 : array_index_85257[3];
  assign array_update_85260[4] = add_85259 == 32'h0000_0004 ? 32'h0000_0000 : array_index_85257[4];
  assign array_update_85260[5] = add_85259 == 32'h0000_0005 ? 32'h0000_0000 : array_index_85257[5];
  assign array_update_85260[6] = add_85259 == 32'h0000_0006 ? 32'h0000_0000 : array_index_85257[6];
  assign array_update_85260[7] = add_85259 == 32'h0000_0007 ? 32'h0000_0000 : array_index_85257[7];
  assign array_update_85260[8] = add_85259 == 32'h0000_0008 ? 32'h0000_0000 : array_index_85257[8];
  assign array_update_85260[9] = add_85259 == 32'h0000_0009 ? 32'h0000_0000 : array_index_85257[9];
  assign literal_85261 = 32'h0000_0000;
  assign array_update_85262[0] = add_84176 == 32'h0000_0000 ? array_update_85260 : array_update_85255[0];
  assign array_update_85262[1] = add_84176 == 32'h0000_0001 ? array_update_85260 : array_update_85255[1];
  assign array_update_85262[2] = add_84176 == 32'h0000_0002 ? array_update_85260 : array_update_85255[2];
  assign array_update_85262[3] = add_84176 == 32'h0000_0003 ? array_update_85260 : array_update_85255[3];
  assign array_update_85262[4] = add_84176 == 32'h0000_0004 ? array_update_85260 : array_update_85255[4];
  assign array_update_85262[5] = add_84176 == 32'h0000_0005 ? array_update_85260 : array_update_85255[5];
  assign array_update_85262[6] = add_84176 == 32'h0000_0006 ? array_update_85260 : array_update_85255[6];
  assign array_update_85262[7] = add_84176 == 32'h0000_0007 ? array_update_85260 : array_update_85255[7];
  assign array_update_85262[8] = add_84176 == 32'h0000_0008 ? array_update_85260 : array_update_85255[8];
  assign array_update_85262[9] = add_84176 == 32'h0000_0009 ? array_update_85260 : array_update_85255[9];
  assign array_index_85264 = array_update_72021[literal_85261 > 32'h0000_0009 ? 4'h9 : literal_85261[3:0]];
  assign array_index_85265 = array_update_85262[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_85269 = smul32b_32b_x_32b(array_index_84183[literal_85261 > 32'h0000_0009 ? 4'h9 : literal_85261[3:0]], array_index_85264[add_85259 > 32'h0000_0009 ? 4'h9 : add_85259[3:0]]);
  assign add_85271 = array_index_85265[add_85259 > 32'h0000_0009 ? 4'h9 : add_85259[3:0]] + smul_85269;
  assign array_update_85273[0] = add_85259 == 32'h0000_0000 ? add_85271 : array_index_85265[0];
  assign array_update_85273[1] = add_85259 == 32'h0000_0001 ? add_85271 : array_index_85265[1];
  assign array_update_85273[2] = add_85259 == 32'h0000_0002 ? add_85271 : array_index_85265[2];
  assign array_update_85273[3] = add_85259 == 32'h0000_0003 ? add_85271 : array_index_85265[3];
  assign array_update_85273[4] = add_85259 == 32'h0000_0004 ? add_85271 : array_index_85265[4];
  assign array_update_85273[5] = add_85259 == 32'h0000_0005 ? add_85271 : array_index_85265[5];
  assign array_update_85273[6] = add_85259 == 32'h0000_0006 ? add_85271 : array_index_85265[6];
  assign array_update_85273[7] = add_85259 == 32'h0000_0007 ? add_85271 : array_index_85265[7];
  assign array_update_85273[8] = add_85259 == 32'h0000_0008 ? add_85271 : array_index_85265[8];
  assign array_update_85273[9] = add_85259 == 32'h0000_0009 ? add_85271 : array_index_85265[9];
  assign add_85274 = literal_85261 + 32'h0000_0001;
  assign array_update_85275[0] = add_84176 == 32'h0000_0000 ? array_update_85273 : array_update_85262[0];
  assign array_update_85275[1] = add_84176 == 32'h0000_0001 ? array_update_85273 : array_update_85262[1];
  assign array_update_85275[2] = add_84176 == 32'h0000_0002 ? array_update_85273 : array_update_85262[2];
  assign array_update_85275[3] = add_84176 == 32'h0000_0003 ? array_update_85273 : array_update_85262[3];
  assign array_update_85275[4] = add_84176 == 32'h0000_0004 ? array_update_85273 : array_update_85262[4];
  assign array_update_85275[5] = add_84176 == 32'h0000_0005 ? array_update_85273 : array_update_85262[5];
  assign array_update_85275[6] = add_84176 == 32'h0000_0006 ? array_update_85273 : array_update_85262[6];
  assign array_update_85275[7] = add_84176 == 32'h0000_0007 ? array_update_85273 : array_update_85262[7];
  assign array_update_85275[8] = add_84176 == 32'h0000_0008 ? array_update_85273 : array_update_85262[8];
  assign array_update_85275[9] = add_84176 == 32'h0000_0009 ? array_update_85273 : array_update_85262[9];
  assign array_index_85277 = array_update_72021[add_85274 > 32'h0000_0009 ? 4'h9 : add_85274[3:0]];
  assign array_index_85278 = array_update_85275[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_85282 = smul32b_32b_x_32b(array_index_84183[add_85274 > 32'h0000_0009 ? 4'h9 : add_85274[3:0]], array_index_85277[add_85259 > 32'h0000_0009 ? 4'h9 : add_85259[3:0]]);
  assign add_85284 = array_index_85278[add_85259 > 32'h0000_0009 ? 4'h9 : add_85259[3:0]] + smul_85282;
  assign array_update_85286[0] = add_85259 == 32'h0000_0000 ? add_85284 : array_index_85278[0];
  assign array_update_85286[1] = add_85259 == 32'h0000_0001 ? add_85284 : array_index_85278[1];
  assign array_update_85286[2] = add_85259 == 32'h0000_0002 ? add_85284 : array_index_85278[2];
  assign array_update_85286[3] = add_85259 == 32'h0000_0003 ? add_85284 : array_index_85278[3];
  assign array_update_85286[4] = add_85259 == 32'h0000_0004 ? add_85284 : array_index_85278[4];
  assign array_update_85286[5] = add_85259 == 32'h0000_0005 ? add_85284 : array_index_85278[5];
  assign array_update_85286[6] = add_85259 == 32'h0000_0006 ? add_85284 : array_index_85278[6];
  assign array_update_85286[7] = add_85259 == 32'h0000_0007 ? add_85284 : array_index_85278[7];
  assign array_update_85286[8] = add_85259 == 32'h0000_0008 ? add_85284 : array_index_85278[8];
  assign array_update_85286[9] = add_85259 == 32'h0000_0009 ? add_85284 : array_index_85278[9];
  assign add_85287 = add_85274 + 32'h0000_0001;
  assign array_update_85288[0] = add_84176 == 32'h0000_0000 ? array_update_85286 : array_update_85275[0];
  assign array_update_85288[1] = add_84176 == 32'h0000_0001 ? array_update_85286 : array_update_85275[1];
  assign array_update_85288[2] = add_84176 == 32'h0000_0002 ? array_update_85286 : array_update_85275[2];
  assign array_update_85288[3] = add_84176 == 32'h0000_0003 ? array_update_85286 : array_update_85275[3];
  assign array_update_85288[4] = add_84176 == 32'h0000_0004 ? array_update_85286 : array_update_85275[4];
  assign array_update_85288[5] = add_84176 == 32'h0000_0005 ? array_update_85286 : array_update_85275[5];
  assign array_update_85288[6] = add_84176 == 32'h0000_0006 ? array_update_85286 : array_update_85275[6];
  assign array_update_85288[7] = add_84176 == 32'h0000_0007 ? array_update_85286 : array_update_85275[7];
  assign array_update_85288[8] = add_84176 == 32'h0000_0008 ? array_update_85286 : array_update_85275[8];
  assign array_update_85288[9] = add_84176 == 32'h0000_0009 ? array_update_85286 : array_update_85275[9];
  assign array_index_85290 = array_update_72021[add_85287 > 32'h0000_0009 ? 4'h9 : add_85287[3:0]];
  assign array_index_85291 = array_update_85288[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_85295 = smul32b_32b_x_32b(array_index_84183[add_85287 > 32'h0000_0009 ? 4'h9 : add_85287[3:0]], array_index_85290[add_85259 > 32'h0000_0009 ? 4'h9 : add_85259[3:0]]);
  assign add_85297 = array_index_85291[add_85259 > 32'h0000_0009 ? 4'h9 : add_85259[3:0]] + smul_85295;
  assign array_update_85299[0] = add_85259 == 32'h0000_0000 ? add_85297 : array_index_85291[0];
  assign array_update_85299[1] = add_85259 == 32'h0000_0001 ? add_85297 : array_index_85291[1];
  assign array_update_85299[2] = add_85259 == 32'h0000_0002 ? add_85297 : array_index_85291[2];
  assign array_update_85299[3] = add_85259 == 32'h0000_0003 ? add_85297 : array_index_85291[3];
  assign array_update_85299[4] = add_85259 == 32'h0000_0004 ? add_85297 : array_index_85291[4];
  assign array_update_85299[5] = add_85259 == 32'h0000_0005 ? add_85297 : array_index_85291[5];
  assign array_update_85299[6] = add_85259 == 32'h0000_0006 ? add_85297 : array_index_85291[6];
  assign array_update_85299[7] = add_85259 == 32'h0000_0007 ? add_85297 : array_index_85291[7];
  assign array_update_85299[8] = add_85259 == 32'h0000_0008 ? add_85297 : array_index_85291[8];
  assign array_update_85299[9] = add_85259 == 32'h0000_0009 ? add_85297 : array_index_85291[9];
  assign add_85300 = add_85287 + 32'h0000_0001;
  assign array_update_85301[0] = add_84176 == 32'h0000_0000 ? array_update_85299 : array_update_85288[0];
  assign array_update_85301[1] = add_84176 == 32'h0000_0001 ? array_update_85299 : array_update_85288[1];
  assign array_update_85301[2] = add_84176 == 32'h0000_0002 ? array_update_85299 : array_update_85288[2];
  assign array_update_85301[3] = add_84176 == 32'h0000_0003 ? array_update_85299 : array_update_85288[3];
  assign array_update_85301[4] = add_84176 == 32'h0000_0004 ? array_update_85299 : array_update_85288[4];
  assign array_update_85301[5] = add_84176 == 32'h0000_0005 ? array_update_85299 : array_update_85288[5];
  assign array_update_85301[6] = add_84176 == 32'h0000_0006 ? array_update_85299 : array_update_85288[6];
  assign array_update_85301[7] = add_84176 == 32'h0000_0007 ? array_update_85299 : array_update_85288[7];
  assign array_update_85301[8] = add_84176 == 32'h0000_0008 ? array_update_85299 : array_update_85288[8];
  assign array_update_85301[9] = add_84176 == 32'h0000_0009 ? array_update_85299 : array_update_85288[9];
  assign array_index_85303 = array_update_72021[add_85300 > 32'h0000_0009 ? 4'h9 : add_85300[3:0]];
  assign array_index_85304 = array_update_85301[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_85308 = smul32b_32b_x_32b(array_index_84183[add_85300 > 32'h0000_0009 ? 4'h9 : add_85300[3:0]], array_index_85303[add_85259 > 32'h0000_0009 ? 4'h9 : add_85259[3:0]]);
  assign add_85310 = array_index_85304[add_85259 > 32'h0000_0009 ? 4'h9 : add_85259[3:0]] + smul_85308;
  assign array_update_85312[0] = add_85259 == 32'h0000_0000 ? add_85310 : array_index_85304[0];
  assign array_update_85312[1] = add_85259 == 32'h0000_0001 ? add_85310 : array_index_85304[1];
  assign array_update_85312[2] = add_85259 == 32'h0000_0002 ? add_85310 : array_index_85304[2];
  assign array_update_85312[3] = add_85259 == 32'h0000_0003 ? add_85310 : array_index_85304[3];
  assign array_update_85312[4] = add_85259 == 32'h0000_0004 ? add_85310 : array_index_85304[4];
  assign array_update_85312[5] = add_85259 == 32'h0000_0005 ? add_85310 : array_index_85304[5];
  assign array_update_85312[6] = add_85259 == 32'h0000_0006 ? add_85310 : array_index_85304[6];
  assign array_update_85312[7] = add_85259 == 32'h0000_0007 ? add_85310 : array_index_85304[7];
  assign array_update_85312[8] = add_85259 == 32'h0000_0008 ? add_85310 : array_index_85304[8];
  assign array_update_85312[9] = add_85259 == 32'h0000_0009 ? add_85310 : array_index_85304[9];
  assign add_85313 = add_85300 + 32'h0000_0001;
  assign array_update_85314[0] = add_84176 == 32'h0000_0000 ? array_update_85312 : array_update_85301[0];
  assign array_update_85314[1] = add_84176 == 32'h0000_0001 ? array_update_85312 : array_update_85301[1];
  assign array_update_85314[2] = add_84176 == 32'h0000_0002 ? array_update_85312 : array_update_85301[2];
  assign array_update_85314[3] = add_84176 == 32'h0000_0003 ? array_update_85312 : array_update_85301[3];
  assign array_update_85314[4] = add_84176 == 32'h0000_0004 ? array_update_85312 : array_update_85301[4];
  assign array_update_85314[5] = add_84176 == 32'h0000_0005 ? array_update_85312 : array_update_85301[5];
  assign array_update_85314[6] = add_84176 == 32'h0000_0006 ? array_update_85312 : array_update_85301[6];
  assign array_update_85314[7] = add_84176 == 32'h0000_0007 ? array_update_85312 : array_update_85301[7];
  assign array_update_85314[8] = add_84176 == 32'h0000_0008 ? array_update_85312 : array_update_85301[8];
  assign array_update_85314[9] = add_84176 == 32'h0000_0009 ? array_update_85312 : array_update_85301[9];
  assign array_index_85316 = array_update_72021[add_85313 > 32'h0000_0009 ? 4'h9 : add_85313[3:0]];
  assign array_index_85317 = array_update_85314[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_85321 = smul32b_32b_x_32b(array_index_84183[add_85313 > 32'h0000_0009 ? 4'h9 : add_85313[3:0]], array_index_85316[add_85259 > 32'h0000_0009 ? 4'h9 : add_85259[3:0]]);
  assign add_85323 = array_index_85317[add_85259 > 32'h0000_0009 ? 4'h9 : add_85259[3:0]] + smul_85321;
  assign array_update_85325[0] = add_85259 == 32'h0000_0000 ? add_85323 : array_index_85317[0];
  assign array_update_85325[1] = add_85259 == 32'h0000_0001 ? add_85323 : array_index_85317[1];
  assign array_update_85325[2] = add_85259 == 32'h0000_0002 ? add_85323 : array_index_85317[2];
  assign array_update_85325[3] = add_85259 == 32'h0000_0003 ? add_85323 : array_index_85317[3];
  assign array_update_85325[4] = add_85259 == 32'h0000_0004 ? add_85323 : array_index_85317[4];
  assign array_update_85325[5] = add_85259 == 32'h0000_0005 ? add_85323 : array_index_85317[5];
  assign array_update_85325[6] = add_85259 == 32'h0000_0006 ? add_85323 : array_index_85317[6];
  assign array_update_85325[7] = add_85259 == 32'h0000_0007 ? add_85323 : array_index_85317[7];
  assign array_update_85325[8] = add_85259 == 32'h0000_0008 ? add_85323 : array_index_85317[8];
  assign array_update_85325[9] = add_85259 == 32'h0000_0009 ? add_85323 : array_index_85317[9];
  assign add_85326 = add_85313 + 32'h0000_0001;
  assign array_update_85327[0] = add_84176 == 32'h0000_0000 ? array_update_85325 : array_update_85314[0];
  assign array_update_85327[1] = add_84176 == 32'h0000_0001 ? array_update_85325 : array_update_85314[1];
  assign array_update_85327[2] = add_84176 == 32'h0000_0002 ? array_update_85325 : array_update_85314[2];
  assign array_update_85327[3] = add_84176 == 32'h0000_0003 ? array_update_85325 : array_update_85314[3];
  assign array_update_85327[4] = add_84176 == 32'h0000_0004 ? array_update_85325 : array_update_85314[4];
  assign array_update_85327[5] = add_84176 == 32'h0000_0005 ? array_update_85325 : array_update_85314[5];
  assign array_update_85327[6] = add_84176 == 32'h0000_0006 ? array_update_85325 : array_update_85314[6];
  assign array_update_85327[7] = add_84176 == 32'h0000_0007 ? array_update_85325 : array_update_85314[7];
  assign array_update_85327[8] = add_84176 == 32'h0000_0008 ? array_update_85325 : array_update_85314[8];
  assign array_update_85327[9] = add_84176 == 32'h0000_0009 ? array_update_85325 : array_update_85314[9];
  assign array_index_85329 = array_update_72021[add_85326 > 32'h0000_0009 ? 4'h9 : add_85326[3:0]];
  assign array_index_85330 = array_update_85327[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_85334 = smul32b_32b_x_32b(array_index_84183[add_85326 > 32'h0000_0009 ? 4'h9 : add_85326[3:0]], array_index_85329[add_85259 > 32'h0000_0009 ? 4'h9 : add_85259[3:0]]);
  assign add_85336 = array_index_85330[add_85259 > 32'h0000_0009 ? 4'h9 : add_85259[3:0]] + smul_85334;
  assign array_update_85338[0] = add_85259 == 32'h0000_0000 ? add_85336 : array_index_85330[0];
  assign array_update_85338[1] = add_85259 == 32'h0000_0001 ? add_85336 : array_index_85330[1];
  assign array_update_85338[2] = add_85259 == 32'h0000_0002 ? add_85336 : array_index_85330[2];
  assign array_update_85338[3] = add_85259 == 32'h0000_0003 ? add_85336 : array_index_85330[3];
  assign array_update_85338[4] = add_85259 == 32'h0000_0004 ? add_85336 : array_index_85330[4];
  assign array_update_85338[5] = add_85259 == 32'h0000_0005 ? add_85336 : array_index_85330[5];
  assign array_update_85338[6] = add_85259 == 32'h0000_0006 ? add_85336 : array_index_85330[6];
  assign array_update_85338[7] = add_85259 == 32'h0000_0007 ? add_85336 : array_index_85330[7];
  assign array_update_85338[8] = add_85259 == 32'h0000_0008 ? add_85336 : array_index_85330[8];
  assign array_update_85338[9] = add_85259 == 32'h0000_0009 ? add_85336 : array_index_85330[9];
  assign add_85339 = add_85326 + 32'h0000_0001;
  assign array_update_85340[0] = add_84176 == 32'h0000_0000 ? array_update_85338 : array_update_85327[0];
  assign array_update_85340[1] = add_84176 == 32'h0000_0001 ? array_update_85338 : array_update_85327[1];
  assign array_update_85340[2] = add_84176 == 32'h0000_0002 ? array_update_85338 : array_update_85327[2];
  assign array_update_85340[3] = add_84176 == 32'h0000_0003 ? array_update_85338 : array_update_85327[3];
  assign array_update_85340[4] = add_84176 == 32'h0000_0004 ? array_update_85338 : array_update_85327[4];
  assign array_update_85340[5] = add_84176 == 32'h0000_0005 ? array_update_85338 : array_update_85327[5];
  assign array_update_85340[6] = add_84176 == 32'h0000_0006 ? array_update_85338 : array_update_85327[6];
  assign array_update_85340[7] = add_84176 == 32'h0000_0007 ? array_update_85338 : array_update_85327[7];
  assign array_update_85340[8] = add_84176 == 32'h0000_0008 ? array_update_85338 : array_update_85327[8];
  assign array_update_85340[9] = add_84176 == 32'h0000_0009 ? array_update_85338 : array_update_85327[9];
  assign array_index_85342 = array_update_72021[add_85339 > 32'h0000_0009 ? 4'h9 : add_85339[3:0]];
  assign array_index_85343 = array_update_85340[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_85347 = smul32b_32b_x_32b(array_index_84183[add_85339 > 32'h0000_0009 ? 4'h9 : add_85339[3:0]], array_index_85342[add_85259 > 32'h0000_0009 ? 4'h9 : add_85259[3:0]]);
  assign add_85349 = array_index_85343[add_85259 > 32'h0000_0009 ? 4'h9 : add_85259[3:0]] + smul_85347;
  assign array_update_85351[0] = add_85259 == 32'h0000_0000 ? add_85349 : array_index_85343[0];
  assign array_update_85351[1] = add_85259 == 32'h0000_0001 ? add_85349 : array_index_85343[1];
  assign array_update_85351[2] = add_85259 == 32'h0000_0002 ? add_85349 : array_index_85343[2];
  assign array_update_85351[3] = add_85259 == 32'h0000_0003 ? add_85349 : array_index_85343[3];
  assign array_update_85351[4] = add_85259 == 32'h0000_0004 ? add_85349 : array_index_85343[4];
  assign array_update_85351[5] = add_85259 == 32'h0000_0005 ? add_85349 : array_index_85343[5];
  assign array_update_85351[6] = add_85259 == 32'h0000_0006 ? add_85349 : array_index_85343[6];
  assign array_update_85351[7] = add_85259 == 32'h0000_0007 ? add_85349 : array_index_85343[7];
  assign array_update_85351[8] = add_85259 == 32'h0000_0008 ? add_85349 : array_index_85343[8];
  assign array_update_85351[9] = add_85259 == 32'h0000_0009 ? add_85349 : array_index_85343[9];
  assign add_85352 = add_85339 + 32'h0000_0001;
  assign array_update_85353[0] = add_84176 == 32'h0000_0000 ? array_update_85351 : array_update_85340[0];
  assign array_update_85353[1] = add_84176 == 32'h0000_0001 ? array_update_85351 : array_update_85340[1];
  assign array_update_85353[2] = add_84176 == 32'h0000_0002 ? array_update_85351 : array_update_85340[2];
  assign array_update_85353[3] = add_84176 == 32'h0000_0003 ? array_update_85351 : array_update_85340[3];
  assign array_update_85353[4] = add_84176 == 32'h0000_0004 ? array_update_85351 : array_update_85340[4];
  assign array_update_85353[5] = add_84176 == 32'h0000_0005 ? array_update_85351 : array_update_85340[5];
  assign array_update_85353[6] = add_84176 == 32'h0000_0006 ? array_update_85351 : array_update_85340[6];
  assign array_update_85353[7] = add_84176 == 32'h0000_0007 ? array_update_85351 : array_update_85340[7];
  assign array_update_85353[8] = add_84176 == 32'h0000_0008 ? array_update_85351 : array_update_85340[8];
  assign array_update_85353[9] = add_84176 == 32'h0000_0009 ? array_update_85351 : array_update_85340[9];
  assign array_index_85355 = array_update_72021[add_85352 > 32'h0000_0009 ? 4'h9 : add_85352[3:0]];
  assign array_index_85356 = array_update_85353[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_85360 = smul32b_32b_x_32b(array_index_84183[add_85352 > 32'h0000_0009 ? 4'h9 : add_85352[3:0]], array_index_85355[add_85259 > 32'h0000_0009 ? 4'h9 : add_85259[3:0]]);
  assign add_85362 = array_index_85356[add_85259 > 32'h0000_0009 ? 4'h9 : add_85259[3:0]] + smul_85360;
  assign array_update_85364[0] = add_85259 == 32'h0000_0000 ? add_85362 : array_index_85356[0];
  assign array_update_85364[1] = add_85259 == 32'h0000_0001 ? add_85362 : array_index_85356[1];
  assign array_update_85364[2] = add_85259 == 32'h0000_0002 ? add_85362 : array_index_85356[2];
  assign array_update_85364[3] = add_85259 == 32'h0000_0003 ? add_85362 : array_index_85356[3];
  assign array_update_85364[4] = add_85259 == 32'h0000_0004 ? add_85362 : array_index_85356[4];
  assign array_update_85364[5] = add_85259 == 32'h0000_0005 ? add_85362 : array_index_85356[5];
  assign array_update_85364[6] = add_85259 == 32'h0000_0006 ? add_85362 : array_index_85356[6];
  assign array_update_85364[7] = add_85259 == 32'h0000_0007 ? add_85362 : array_index_85356[7];
  assign array_update_85364[8] = add_85259 == 32'h0000_0008 ? add_85362 : array_index_85356[8];
  assign array_update_85364[9] = add_85259 == 32'h0000_0009 ? add_85362 : array_index_85356[9];
  assign add_85365 = add_85352 + 32'h0000_0001;
  assign array_update_85366[0] = add_84176 == 32'h0000_0000 ? array_update_85364 : array_update_85353[0];
  assign array_update_85366[1] = add_84176 == 32'h0000_0001 ? array_update_85364 : array_update_85353[1];
  assign array_update_85366[2] = add_84176 == 32'h0000_0002 ? array_update_85364 : array_update_85353[2];
  assign array_update_85366[3] = add_84176 == 32'h0000_0003 ? array_update_85364 : array_update_85353[3];
  assign array_update_85366[4] = add_84176 == 32'h0000_0004 ? array_update_85364 : array_update_85353[4];
  assign array_update_85366[5] = add_84176 == 32'h0000_0005 ? array_update_85364 : array_update_85353[5];
  assign array_update_85366[6] = add_84176 == 32'h0000_0006 ? array_update_85364 : array_update_85353[6];
  assign array_update_85366[7] = add_84176 == 32'h0000_0007 ? array_update_85364 : array_update_85353[7];
  assign array_update_85366[8] = add_84176 == 32'h0000_0008 ? array_update_85364 : array_update_85353[8];
  assign array_update_85366[9] = add_84176 == 32'h0000_0009 ? array_update_85364 : array_update_85353[9];
  assign array_index_85368 = array_update_72021[add_85365 > 32'h0000_0009 ? 4'h9 : add_85365[3:0]];
  assign array_index_85369 = array_update_85366[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_85373 = smul32b_32b_x_32b(array_index_84183[add_85365 > 32'h0000_0009 ? 4'h9 : add_85365[3:0]], array_index_85368[add_85259 > 32'h0000_0009 ? 4'h9 : add_85259[3:0]]);
  assign add_85375 = array_index_85369[add_85259 > 32'h0000_0009 ? 4'h9 : add_85259[3:0]] + smul_85373;
  assign array_update_85377[0] = add_85259 == 32'h0000_0000 ? add_85375 : array_index_85369[0];
  assign array_update_85377[1] = add_85259 == 32'h0000_0001 ? add_85375 : array_index_85369[1];
  assign array_update_85377[2] = add_85259 == 32'h0000_0002 ? add_85375 : array_index_85369[2];
  assign array_update_85377[3] = add_85259 == 32'h0000_0003 ? add_85375 : array_index_85369[3];
  assign array_update_85377[4] = add_85259 == 32'h0000_0004 ? add_85375 : array_index_85369[4];
  assign array_update_85377[5] = add_85259 == 32'h0000_0005 ? add_85375 : array_index_85369[5];
  assign array_update_85377[6] = add_85259 == 32'h0000_0006 ? add_85375 : array_index_85369[6];
  assign array_update_85377[7] = add_85259 == 32'h0000_0007 ? add_85375 : array_index_85369[7];
  assign array_update_85377[8] = add_85259 == 32'h0000_0008 ? add_85375 : array_index_85369[8];
  assign array_update_85377[9] = add_85259 == 32'h0000_0009 ? add_85375 : array_index_85369[9];
  assign add_85378 = add_85365 + 32'h0000_0001;
  assign array_update_85379[0] = add_84176 == 32'h0000_0000 ? array_update_85377 : array_update_85366[0];
  assign array_update_85379[1] = add_84176 == 32'h0000_0001 ? array_update_85377 : array_update_85366[1];
  assign array_update_85379[2] = add_84176 == 32'h0000_0002 ? array_update_85377 : array_update_85366[2];
  assign array_update_85379[3] = add_84176 == 32'h0000_0003 ? array_update_85377 : array_update_85366[3];
  assign array_update_85379[4] = add_84176 == 32'h0000_0004 ? array_update_85377 : array_update_85366[4];
  assign array_update_85379[5] = add_84176 == 32'h0000_0005 ? array_update_85377 : array_update_85366[5];
  assign array_update_85379[6] = add_84176 == 32'h0000_0006 ? array_update_85377 : array_update_85366[6];
  assign array_update_85379[7] = add_84176 == 32'h0000_0007 ? array_update_85377 : array_update_85366[7];
  assign array_update_85379[8] = add_84176 == 32'h0000_0008 ? array_update_85377 : array_update_85366[8];
  assign array_update_85379[9] = add_84176 == 32'h0000_0009 ? array_update_85377 : array_update_85366[9];
  assign array_index_85381 = array_update_72021[add_85378 > 32'h0000_0009 ? 4'h9 : add_85378[3:0]];
  assign array_index_85383 = array_update_85379[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_85388 = smul32b_32b_x_32b(array_index_84183[add_85378 > 32'h0000_0009 ? 4'h9 : add_85378[3:0]], array_index_85381[add_85259 > 32'h0000_0009 ? 4'h9 : add_85259[3:0]]);
  assign add_85391 = array_index_85383[add_85259 > 32'h0000_0009 ? 4'h9 : add_85259[3:0]] + smul_85388;
  assign array_update_85393[0] = add_85259 == 32'h0000_0000 ? add_85391 : array_index_85383[0];
  assign array_update_85393[1] = add_85259 == 32'h0000_0001 ? add_85391 : array_index_85383[1];
  assign array_update_85393[2] = add_85259 == 32'h0000_0002 ? add_85391 : array_index_85383[2];
  assign array_update_85393[3] = add_85259 == 32'h0000_0003 ? add_85391 : array_index_85383[3];
  assign array_update_85393[4] = add_85259 == 32'h0000_0004 ? add_85391 : array_index_85383[4];
  assign array_update_85393[5] = add_85259 == 32'h0000_0005 ? add_85391 : array_index_85383[5];
  assign array_update_85393[6] = add_85259 == 32'h0000_0006 ? add_85391 : array_index_85383[6];
  assign array_update_85393[7] = add_85259 == 32'h0000_0007 ? add_85391 : array_index_85383[7];
  assign array_update_85393[8] = add_85259 == 32'h0000_0008 ? add_85391 : array_index_85383[8];
  assign array_update_85393[9] = add_85259 == 32'h0000_0009 ? add_85391 : array_index_85383[9];
  assign array_update_85397[0] = add_84176 == 32'h0000_0000 ? array_update_85393 : array_update_85379[0];
  assign array_update_85397[1] = add_84176 == 32'h0000_0001 ? array_update_85393 : array_update_85379[1];
  assign array_update_85397[2] = add_84176 == 32'h0000_0002 ? array_update_85393 : array_update_85379[2];
  assign array_update_85397[3] = add_84176 == 32'h0000_0003 ? array_update_85393 : array_update_85379[3];
  assign array_update_85397[4] = add_84176 == 32'h0000_0004 ? array_update_85393 : array_update_85379[4];
  assign array_update_85397[5] = add_84176 == 32'h0000_0005 ? array_update_85393 : array_update_85379[5];
  assign array_update_85397[6] = add_84176 == 32'h0000_0006 ? array_update_85393 : array_update_85379[6];
  assign array_update_85397[7] = add_84176 == 32'h0000_0007 ? array_update_85393 : array_update_85379[7];
  assign array_update_85397[8] = add_84176 == 32'h0000_0008 ? array_update_85393 : array_update_85379[8];
  assign array_update_85397[9] = add_84176 == 32'h0000_0009 ? array_update_85393 : array_update_85379[9];
  assign array_index_85401 = array_update_85397[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign add_85403 = add_85259 + 32'h0000_0001;
  assign array_update_85407[0] = add_85403 == 32'h0000_0000 ? 32'h0000_0000 : array_index_85401[0];
  assign array_update_85407[1] = add_85403 == 32'h0000_0001 ? 32'h0000_0000 : array_index_85401[1];
  assign array_update_85407[2] = add_85403 == 32'h0000_0002 ? 32'h0000_0000 : array_index_85401[2];
  assign array_update_85407[3] = add_85403 == 32'h0000_0003 ? 32'h0000_0000 : array_index_85401[3];
  assign array_update_85407[4] = add_85403 == 32'h0000_0004 ? 32'h0000_0000 : array_index_85401[4];
  assign array_update_85407[5] = add_85403 == 32'h0000_0005 ? 32'h0000_0000 : array_index_85401[5];
  assign array_update_85407[6] = add_85403 == 32'h0000_0006 ? 32'h0000_0000 : array_index_85401[6];
  assign array_update_85407[7] = add_85403 == 32'h0000_0007 ? 32'h0000_0000 : array_index_85401[7];
  assign array_update_85407[8] = add_85403 == 32'h0000_0008 ? 32'h0000_0000 : array_index_85401[8];
  assign array_update_85407[9] = add_85403 == 32'h0000_0009 ? 32'h0000_0000 : array_index_85401[9];
  assign literal_85408 = 32'h0000_0000;
  assign array_update_85411[0] = add_84176 == 32'h0000_0000 ? array_update_85407 : array_update_85397[0];
  assign array_update_85411[1] = add_84176 == 32'h0000_0001 ? array_update_85407 : array_update_85397[1];
  assign array_update_85411[2] = add_84176 == 32'h0000_0002 ? array_update_85407 : array_update_85397[2];
  assign array_update_85411[3] = add_84176 == 32'h0000_0003 ? array_update_85407 : array_update_85397[3];
  assign array_update_85411[4] = add_84176 == 32'h0000_0004 ? array_update_85407 : array_update_85397[4];
  assign array_update_85411[5] = add_84176 == 32'h0000_0005 ? array_update_85407 : array_update_85397[5];
  assign array_update_85411[6] = add_84176 == 32'h0000_0006 ? array_update_85407 : array_update_85397[6];
  assign array_update_85411[7] = add_84176 == 32'h0000_0007 ? array_update_85407 : array_update_85397[7];
  assign array_update_85411[8] = add_84176 == 32'h0000_0008 ? array_update_85407 : array_update_85397[8];
  assign array_update_85411[9] = add_84176 == 32'h0000_0009 ? array_update_85407 : array_update_85397[9];
  assign array_index_85413 = array_update_72021[literal_85408 > 32'h0000_0009 ? 4'h9 : literal_85408[3:0]];
  assign array_index_85417 = array_update_85411[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_85423 = smul32b_32b_x_32b(array_index_84183[literal_85408 > 32'h0000_0009 ? 4'h9 : literal_85408[3:0]], array_index_85413[add_85403 > 32'h0000_0009 ? 4'h9 : add_85403[3:0]]);
  assign add_85428 = array_index_85417[add_85403 > 32'h0000_0009 ? 4'h9 : add_85403[3:0]] + smul_85423;
  assign array_update_85432[0] = add_85403 == 32'h0000_0000 ? add_85428 : array_index_85417[0];
  assign array_update_85432[1] = add_85403 == 32'h0000_0001 ? add_85428 : array_index_85417[1];
  assign array_update_85432[2] = add_85403 == 32'h0000_0002 ? add_85428 : array_index_85417[2];
  assign array_update_85432[3] = add_85403 == 32'h0000_0003 ? add_85428 : array_index_85417[3];
  assign array_update_85432[4] = add_85403 == 32'h0000_0004 ? add_85428 : array_index_85417[4];
  assign array_update_85432[5] = add_85403 == 32'h0000_0005 ? add_85428 : array_index_85417[5];
  assign array_update_85432[6] = add_85403 == 32'h0000_0006 ? add_85428 : array_index_85417[6];
  assign array_update_85432[7] = add_85403 == 32'h0000_0007 ? add_85428 : array_index_85417[7];
  assign array_update_85432[8] = add_85403 == 32'h0000_0008 ? add_85428 : array_index_85417[8];
  assign array_update_85432[9] = add_85403 == 32'h0000_0009 ? add_85428 : array_index_85417[9];
  assign add_85433 = literal_85408 + 32'h0000_0001;
  assign array_update_85437[0] = add_84176 == 32'h0000_0000 ? array_update_85432 : array_update_85411[0];
  assign array_update_85437[1] = add_84176 == 32'h0000_0001 ? array_update_85432 : array_update_85411[1];
  assign array_update_85437[2] = add_84176 == 32'h0000_0002 ? array_update_85432 : array_update_85411[2];
  assign array_update_85437[3] = add_84176 == 32'h0000_0003 ? array_update_85432 : array_update_85411[3];
  assign array_update_85437[4] = add_84176 == 32'h0000_0004 ? array_update_85432 : array_update_85411[4];
  assign array_update_85437[5] = add_84176 == 32'h0000_0005 ? array_update_85432 : array_update_85411[5];
  assign array_update_85437[6] = add_84176 == 32'h0000_0006 ? array_update_85432 : array_update_85411[6];
  assign array_update_85437[7] = add_84176 == 32'h0000_0007 ? array_update_85432 : array_update_85411[7];
  assign array_update_85437[8] = add_84176 == 32'h0000_0008 ? array_update_85432 : array_update_85411[8];
  assign array_update_85437[9] = add_84176 == 32'h0000_0009 ? array_update_85432 : array_update_85411[9];
  assign array_index_85439 = array_update_72021[add_85433 > 32'h0000_0009 ? 4'h9 : add_85433[3:0]];
  assign array_index_85442 = array_update_85437[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_85449 = smul32b_32b_x_32b(array_index_84183[add_85433 > 32'h0000_0009 ? 4'h9 : add_85433[3:0]], array_index_85439[add_85403 > 32'h0000_0009 ? 4'h9 : add_85403[3:0]]);
  assign add_85453 = array_index_85442[add_85403 > 32'h0000_0009 ? 4'h9 : add_85403[3:0]] + smul_85449;
  assign array_update_85458[0] = add_85403 == 32'h0000_0000 ? add_85453 : array_index_85442[0];
  assign array_update_85458[1] = add_85403 == 32'h0000_0001 ? add_85453 : array_index_85442[1];
  assign array_update_85458[2] = add_85403 == 32'h0000_0002 ? add_85453 : array_index_85442[2];
  assign array_update_85458[3] = add_85403 == 32'h0000_0003 ? add_85453 : array_index_85442[3];
  assign array_update_85458[4] = add_85403 == 32'h0000_0004 ? add_85453 : array_index_85442[4];
  assign array_update_85458[5] = add_85403 == 32'h0000_0005 ? add_85453 : array_index_85442[5];
  assign array_update_85458[6] = add_85403 == 32'h0000_0006 ? add_85453 : array_index_85442[6];
  assign array_update_85458[7] = add_85403 == 32'h0000_0007 ? add_85453 : array_index_85442[7];
  assign array_update_85458[8] = add_85403 == 32'h0000_0008 ? add_85453 : array_index_85442[8];
  assign array_update_85458[9] = add_85403 == 32'h0000_0009 ? add_85453 : array_index_85442[9];
  assign add_85459 = add_85433 + 32'h0000_0001;
  assign array_update_85462[0] = add_84176 == 32'h0000_0000 ? array_update_85458 : array_update_85437[0];
  assign array_update_85462[1] = add_84176 == 32'h0000_0001 ? array_update_85458 : array_update_85437[1];
  assign array_update_85462[2] = add_84176 == 32'h0000_0002 ? array_update_85458 : array_update_85437[2];
  assign array_update_85462[3] = add_84176 == 32'h0000_0003 ? array_update_85458 : array_update_85437[3];
  assign array_update_85462[4] = add_84176 == 32'h0000_0004 ? array_update_85458 : array_update_85437[4];
  assign array_update_85462[5] = add_84176 == 32'h0000_0005 ? array_update_85458 : array_update_85437[5];
  assign array_update_85462[6] = add_84176 == 32'h0000_0006 ? array_update_85458 : array_update_85437[6];
  assign array_update_85462[7] = add_84176 == 32'h0000_0007 ? array_update_85458 : array_update_85437[7];
  assign array_update_85462[8] = add_84176 == 32'h0000_0008 ? array_update_85458 : array_update_85437[8];
  assign array_update_85462[9] = add_84176 == 32'h0000_0009 ? array_update_85458 : array_update_85437[9];
  assign array_index_85464 = array_update_72021[add_85459 > 32'h0000_0009 ? 4'h9 : add_85459[3:0]];
  assign array_index_85468 = array_update_85462[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_85474 = smul32b_32b_x_32b(array_index_84183[add_85459 > 32'h0000_0009 ? 4'h9 : add_85459[3:0]], array_index_85464[add_85403 > 32'h0000_0009 ? 4'h9 : add_85403[3:0]]);
  assign add_85479 = array_index_85468[add_85403 > 32'h0000_0009 ? 4'h9 : add_85403[3:0]] + smul_85474;
  assign array_update_85502[0] = add_85403 == 32'h0000_0000 ? add_85479 : array_index_85468[0];
  assign array_update_85502[1] = add_85403 == 32'h0000_0001 ? add_85479 : array_index_85468[1];
  assign array_update_85502[2] = add_85403 == 32'h0000_0002 ? add_85479 : array_index_85468[2];
  assign array_update_85502[3] = add_85403 == 32'h0000_0003 ? add_85479 : array_index_85468[3];
  assign array_update_85502[4] = add_85403 == 32'h0000_0004 ? add_85479 : array_index_85468[4];
  assign array_update_85502[5] = add_85403 == 32'h0000_0005 ? add_85479 : array_index_85468[5];
  assign array_update_85502[6] = add_85403 == 32'h0000_0006 ? add_85479 : array_index_85468[6];
  assign array_update_85502[7] = add_85403 == 32'h0000_0007 ? add_85479 : array_index_85468[7];
  assign array_update_85502[8] = add_85403 == 32'h0000_0008 ? add_85479 : array_index_85468[8];
  assign array_update_85502[9] = add_85403 == 32'h0000_0009 ? add_85479 : array_index_85468[9];
  assign add_85503 = add_85459 + 32'h0000_0001;
  assign array_update_85524[0] = add_84176 == 32'h0000_0000 ? array_update_85502 : array_update_85462[0];
  assign array_update_85524[1] = add_84176 == 32'h0000_0001 ? array_update_85502 : array_update_85462[1];
  assign array_update_85524[2] = add_84176 == 32'h0000_0002 ? array_update_85502 : array_update_85462[2];
  assign array_update_85524[3] = add_84176 == 32'h0000_0003 ? array_update_85502 : array_update_85462[3];
  assign array_update_85524[4] = add_84176 == 32'h0000_0004 ? array_update_85502 : array_update_85462[4];
  assign array_update_85524[5] = add_84176 == 32'h0000_0005 ? array_update_85502 : array_update_85462[5];
  assign array_update_85524[6] = add_84176 == 32'h0000_0006 ? array_update_85502 : array_update_85462[6];
  assign array_update_85524[7] = add_84176 == 32'h0000_0007 ? array_update_85502 : array_update_85462[7];
  assign array_update_85524[8] = add_84176 == 32'h0000_0008 ? array_update_85502 : array_update_85462[8];
  assign array_update_85524[9] = add_84176 == 32'h0000_0009 ? array_update_85502 : array_update_85462[9];
  assign array_index_85526 = array_update_72021[add_85503 > 32'h0000_0009 ? 4'h9 : add_85503[3:0]];
  assign array_index_85557 = array_update_85524[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_85581 = smul32b_32b_x_32b(array_index_84183[add_85503 > 32'h0000_0009 ? 4'h9 : add_85503[3:0]], array_index_85526[add_85403 > 32'h0000_0009 ? 4'h9 : add_85403[3:0]]);
  assign add_85613 = array_index_85557[add_85403 > 32'h0000_0009 ? 4'h9 : add_85403[3:0]] + smul_85581;
  assign array_update_85635[0] = add_85403 == 32'h0000_0000 ? add_85613 : array_index_85557[0];
  assign array_update_85635[1] = add_85403 == 32'h0000_0001 ? add_85613 : array_index_85557[1];
  assign array_update_85635[2] = add_85403 == 32'h0000_0002 ? add_85613 : array_index_85557[2];
  assign array_update_85635[3] = add_85403 == 32'h0000_0003 ? add_85613 : array_index_85557[3];
  assign array_update_85635[4] = add_85403 == 32'h0000_0004 ? add_85613 : array_index_85557[4];
  assign array_update_85635[5] = add_85403 == 32'h0000_0005 ? add_85613 : array_index_85557[5];
  assign array_update_85635[6] = add_85403 == 32'h0000_0006 ? add_85613 : array_index_85557[6];
  assign array_update_85635[7] = add_85403 == 32'h0000_0007 ? add_85613 : array_index_85557[7];
  assign array_update_85635[8] = add_85403 == 32'h0000_0008 ? add_85613 : array_index_85557[8];
  assign array_update_85635[9] = add_85403 == 32'h0000_0009 ? add_85613 : array_index_85557[9];
  assign add_85636 = add_85503 + 32'h0000_0001;
  assign array_update_85667[0] = add_84176 == 32'h0000_0000 ? array_update_85635 : array_update_85524[0];
  assign array_update_85667[1] = add_84176 == 32'h0000_0001 ? array_update_85635 : array_update_85524[1];
  assign array_update_85667[2] = add_84176 == 32'h0000_0002 ? array_update_85635 : array_update_85524[2];
  assign array_update_85667[3] = add_84176 == 32'h0000_0003 ? array_update_85635 : array_update_85524[3];
  assign array_update_85667[4] = add_84176 == 32'h0000_0004 ? array_update_85635 : array_update_85524[4];
  assign array_update_85667[5] = add_84176 == 32'h0000_0005 ? array_update_85635 : array_update_85524[5];
  assign array_update_85667[6] = add_84176 == 32'h0000_0006 ? array_update_85635 : array_update_85524[6];
  assign array_update_85667[7] = add_84176 == 32'h0000_0007 ? array_update_85635 : array_update_85524[7];
  assign array_update_85667[8] = add_84176 == 32'h0000_0008 ? array_update_85635 : array_update_85524[8];
  assign array_update_85667[9] = add_84176 == 32'h0000_0009 ? array_update_85635 : array_update_85524[9];
  assign array_index_85669 = array_update_72021[add_85636 > 32'h0000_0009 ? 4'h9 : add_85636[3:0]];
  assign array_index_85690 = array_update_85667[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_85724 = smul32b_32b_x_32b(array_index_84183[add_85636 > 32'h0000_0009 ? 4'h9 : add_85636[3:0]], array_index_85669[add_85403 > 32'h0000_0009 ? 4'h9 : add_85403[3:0]]);
  assign add_85746 = array_index_85690[add_85403 > 32'h0000_0009 ? 4'h9 : add_85403[3:0]] + smul_85724;
  assign array_update_85778[0] = add_85403 == 32'h0000_0000 ? add_85746 : array_index_85690[0];
  assign array_update_85778[1] = add_85403 == 32'h0000_0001 ? add_85746 : array_index_85690[1];
  assign array_update_85778[2] = add_85403 == 32'h0000_0002 ? add_85746 : array_index_85690[2];
  assign array_update_85778[3] = add_85403 == 32'h0000_0003 ? add_85746 : array_index_85690[3];
  assign array_update_85778[4] = add_85403 == 32'h0000_0004 ? add_85746 : array_index_85690[4];
  assign array_update_85778[5] = add_85403 == 32'h0000_0005 ? add_85746 : array_index_85690[5];
  assign array_update_85778[6] = add_85403 == 32'h0000_0006 ? add_85746 : array_index_85690[6];
  assign array_update_85778[7] = add_85403 == 32'h0000_0007 ? add_85746 : array_index_85690[7];
  assign array_update_85778[8] = add_85403 == 32'h0000_0008 ? add_85746 : array_index_85690[8];
  assign array_update_85778[9] = add_85403 == 32'h0000_0009 ? add_85746 : array_index_85690[9];
  assign add_85779 = add_85636 + 32'h0000_0001;
  assign array_update_85800[0] = add_84176 == 32'h0000_0000 ? array_update_85778 : array_update_85667[0];
  assign array_update_85800[1] = add_84176 == 32'h0000_0001 ? array_update_85778 : array_update_85667[1];
  assign array_update_85800[2] = add_84176 == 32'h0000_0002 ? array_update_85778 : array_update_85667[2];
  assign array_update_85800[3] = add_84176 == 32'h0000_0003 ? array_update_85778 : array_update_85667[3];
  assign array_update_85800[4] = add_84176 == 32'h0000_0004 ? array_update_85778 : array_update_85667[4];
  assign array_update_85800[5] = add_84176 == 32'h0000_0005 ? array_update_85778 : array_update_85667[5];
  assign array_update_85800[6] = add_84176 == 32'h0000_0006 ? array_update_85778 : array_update_85667[6];
  assign array_update_85800[7] = add_84176 == 32'h0000_0007 ? array_update_85778 : array_update_85667[7];
  assign array_update_85800[8] = add_84176 == 32'h0000_0008 ? array_update_85778 : array_update_85667[8];
  assign array_update_85800[9] = add_84176 == 32'h0000_0009 ? array_update_85778 : array_update_85667[9];
  assign array_index_85802 = array_update_72021[add_85779 > 32'h0000_0009 ? 4'h9 : add_85779[3:0]];
  assign array_index_85833 = array_update_85800[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_85857 = smul32b_32b_x_32b(array_index_84183[add_85779 > 32'h0000_0009 ? 4'h9 : add_85779[3:0]], array_index_85802[add_85403 > 32'h0000_0009 ? 4'h9 : add_85403[3:0]]);
  assign add_85889 = array_index_85833[add_85403 > 32'h0000_0009 ? 4'h9 : add_85403[3:0]] + smul_85857;
  assign array_update_85911[0] = add_85403 == 32'h0000_0000 ? add_85889 : array_index_85833[0];
  assign array_update_85911[1] = add_85403 == 32'h0000_0001 ? add_85889 : array_index_85833[1];
  assign array_update_85911[2] = add_85403 == 32'h0000_0002 ? add_85889 : array_index_85833[2];
  assign array_update_85911[3] = add_85403 == 32'h0000_0003 ? add_85889 : array_index_85833[3];
  assign array_update_85911[4] = add_85403 == 32'h0000_0004 ? add_85889 : array_index_85833[4];
  assign array_update_85911[5] = add_85403 == 32'h0000_0005 ? add_85889 : array_index_85833[5];
  assign array_update_85911[6] = add_85403 == 32'h0000_0006 ? add_85889 : array_index_85833[6];
  assign array_update_85911[7] = add_85403 == 32'h0000_0007 ? add_85889 : array_index_85833[7];
  assign array_update_85911[8] = add_85403 == 32'h0000_0008 ? add_85889 : array_index_85833[8];
  assign array_update_85911[9] = add_85403 == 32'h0000_0009 ? add_85889 : array_index_85833[9];
  assign add_85912 = add_85779 + 32'h0000_0001;
  assign array_update_85943[0] = add_84176 == 32'h0000_0000 ? array_update_85911 : array_update_85800[0];
  assign array_update_85943[1] = add_84176 == 32'h0000_0001 ? array_update_85911 : array_update_85800[1];
  assign array_update_85943[2] = add_84176 == 32'h0000_0002 ? array_update_85911 : array_update_85800[2];
  assign array_update_85943[3] = add_84176 == 32'h0000_0003 ? array_update_85911 : array_update_85800[3];
  assign array_update_85943[4] = add_84176 == 32'h0000_0004 ? array_update_85911 : array_update_85800[4];
  assign array_update_85943[5] = add_84176 == 32'h0000_0005 ? array_update_85911 : array_update_85800[5];
  assign array_update_85943[6] = add_84176 == 32'h0000_0006 ? array_update_85911 : array_update_85800[6];
  assign array_update_85943[7] = add_84176 == 32'h0000_0007 ? array_update_85911 : array_update_85800[7];
  assign array_update_85943[8] = add_84176 == 32'h0000_0008 ? array_update_85911 : array_update_85800[8];
  assign array_update_85943[9] = add_84176 == 32'h0000_0009 ? array_update_85911 : array_update_85800[9];
  assign array_index_85945 = array_update_72021[add_85912 > 32'h0000_0009 ? 4'h9 : add_85912[3:0]];
  assign array_index_85966 = array_update_85943[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_85991 = smul32b_32b_x_32b(array_index_84183[add_85912 > 32'h0000_0009 ? 4'h9 : add_85912[3:0]], array_index_85945[add_85403 > 32'h0000_0009 ? 4'h9 : add_85403[3:0]]);
  assign add_86203 = array_index_85966[add_85403 > 32'h0000_0009 ? 4'h9 : add_85403[3:0]] + smul_85991;
  assign array_update_86405[0] = add_85403 == 32'h0000_0000 ? add_86203 : array_index_85966[0];
  assign array_update_86405[1] = add_85403 == 32'h0000_0001 ? add_86203 : array_index_85966[1];
  assign array_update_86405[2] = add_85403 == 32'h0000_0002 ? add_86203 : array_index_85966[2];
  assign array_update_86405[3] = add_85403 == 32'h0000_0003 ? add_86203 : array_index_85966[3];
  assign array_update_86405[4] = add_85403 == 32'h0000_0004 ? add_86203 : array_index_85966[4];
  assign array_update_86405[5] = add_85403 == 32'h0000_0005 ? add_86203 : array_index_85966[5];
  assign array_update_86405[6] = add_85403 == 32'h0000_0006 ? add_86203 : array_index_85966[6];
  assign array_update_86405[7] = add_85403 == 32'h0000_0007 ? add_86203 : array_index_85966[7];
  assign array_update_86405[8] = add_85403 == 32'h0000_0008 ? add_86203 : array_index_85966[8];
  assign array_update_86405[9] = add_85403 == 32'h0000_0009 ? add_86203 : array_index_85966[9];
  assign add_86406 = add_85912 + 32'h0000_0001;
  assign array_update_86707[0] = add_84176 == 32'h0000_0000 ? array_update_86405 : array_update_85943[0];
  assign array_update_86707[1] = add_84176 == 32'h0000_0001 ? array_update_86405 : array_update_85943[1];
  assign array_update_86707[2] = add_84176 == 32'h0000_0002 ? array_update_86405 : array_update_85943[2];
  assign array_update_86707[3] = add_84176 == 32'h0000_0003 ? array_update_86405 : array_update_85943[3];
  assign array_update_86707[4] = add_84176 == 32'h0000_0004 ? array_update_86405 : array_update_85943[4];
  assign array_update_86707[5] = add_84176 == 32'h0000_0005 ? array_update_86405 : array_update_85943[5];
  assign array_update_86707[6] = add_84176 == 32'h0000_0006 ? array_update_86405 : array_update_85943[6];
  assign array_update_86707[7] = add_84176 == 32'h0000_0007 ? array_update_86405 : array_update_85943[7];
  assign array_update_86707[8] = add_84176 == 32'h0000_0008 ? array_update_86405 : array_update_85943[8];
  assign array_update_86707[9] = add_84176 == 32'h0000_0009 ? array_update_86405 : array_update_85943[9];
  assign array_index_86709 = array_update_72021[add_86406 > 32'h0000_0009 ? 4'h9 : add_86406[3:0]];
  assign array_index_86910 = array_update_86707[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign smul_87214 = smul32b_32b_x_32b(array_index_84183[add_86406 > 32'h0000_0009 ? 4'h9 : add_86406[3:0]], array_index_86709[add_85403 > 32'h0000_0009 ? 4'h9 : add_85403[3:0]]);
  assign add_87416 = array_index_86910[add_85403 > 32'h0000_0009 ? 4'h9 : add_85403[3:0]] + smul_87214;
  assign array_update_87718[0] = add_85403 == 32'h0000_0000 ? add_87416 : array_index_86910[0];
  assign array_update_87718[1] = add_85403 == 32'h0000_0001 ? add_87416 : array_index_86910[1];
  assign array_update_87718[2] = add_85403 == 32'h0000_0002 ? add_87416 : array_index_86910[2];
  assign array_update_87718[3] = add_85403 == 32'h0000_0003 ? add_87416 : array_index_86910[3];
  assign array_update_87718[4] = add_85403 == 32'h0000_0004 ? add_87416 : array_index_86910[4];
  assign array_update_87718[5] = add_85403 == 32'h0000_0005 ? add_87416 : array_index_86910[5];
  assign array_update_87718[6] = add_85403 == 32'h0000_0006 ? add_87416 : array_index_86910[6];
  assign array_update_87718[7] = add_85403 == 32'h0000_0007 ? add_87416 : array_index_86910[7];
  assign array_update_87718[8] = add_85403 == 32'h0000_0008 ? add_87416 : array_index_86910[8];
  assign array_update_87718[9] = add_85403 == 32'h0000_0009 ? add_87416 : array_index_86910[9];
  assign add_87719 = add_86406 + 32'h0000_0001;
  assign array_update_87920[0] = add_84176 == 32'h0000_0000 ? array_update_87718 : array_update_86707[0];
  assign array_update_87920[1] = add_84176 == 32'h0000_0001 ? array_update_87718 : array_update_86707[1];
  assign array_update_87920[2] = add_84176 == 32'h0000_0002 ? array_update_87718 : array_update_86707[2];
  assign array_update_87920[3] = add_84176 == 32'h0000_0003 ? array_update_87718 : array_update_86707[3];
  assign array_update_87920[4] = add_84176 == 32'h0000_0004 ? array_update_87718 : array_update_86707[4];
  assign array_update_87920[5] = add_84176 == 32'h0000_0005 ? array_update_87718 : array_update_86707[5];
  assign array_update_87920[6] = add_84176 == 32'h0000_0006 ? array_update_87718 : array_update_86707[6];
  assign array_update_87920[7] = add_84176 == 32'h0000_0007 ? array_update_87718 : array_update_86707[7];
  assign array_update_87920[8] = add_84176 == 32'h0000_0008 ? array_update_87718 : array_update_86707[8];
  assign array_update_87920[9] = add_84176 == 32'h0000_0009 ? array_update_87718 : array_update_86707[9];
  assign array_index_87922 = array_update_72021[add_87719 > 32'h0000_0009 ? 4'h9 : add_87719[3:0]];
  assign array_index_88245 = array_update_87920[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign literal_88243 = 32'h0000_0000;
  assign smul_88471 = smul32b_32b_x_32b(array_index_84183[add_87719 > 32'h0000_0009 ? 4'h9 : add_87719[3:0]], array_index_87922[add_85403 > 32'h0000_0009 ? 4'h9 : add_85403[3:0]]);
  assign literal_88223 = 32'h0000_0000;
  assign literal_88225 = 32'h0000_0000;
  assign literal_88227 = 32'h0000_0000;
  assign literal_88229 = 32'h0000_0000;
  assign literal_88231 = 32'h0000_0000;
  assign literal_88233 = 32'h0000_0000;
  assign literal_88235 = 32'h0000_0000;
  assign literal_88237 = 32'h0000_0000;
  assign literal_88239 = 32'h0000_0000;
  assign add_88468 = literal_88243 + 32'h0000_0001;
  assign literal_88241 = 32'h0000_0000;
  assign add_88795 = array_index_88245[add_85403 > 32'h0000_0009 ? 4'h9 : add_85403[3:0]] + smul_88471;
  assign add_88448 = literal_88223 + 32'h0000_0001;
  assign add_88450 = literal_88225 + 32'h0000_0001;
  assign add_88452 = literal_88227 + 32'h0000_0001;
  assign add_88454 = literal_88229 + 32'h0000_0001;
  assign add_88456 = literal_88231 + 32'h0000_0001;
  assign add_88458 = literal_88233 + 32'h0000_0001;
  assign add_88460 = literal_88235 + 32'h0000_0001;
  assign add_88462 = literal_88237 + 32'h0000_0001;
  assign add_88464 = literal_88239 + 32'h0000_0001;
  assign add_88792 = add_88468 + 32'h0000_0001;
  assign add_88466 = literal_88241 + 32'h0000_0001;
  assign array_update_89019[0] = add_85403 == 32'h0000_0000 ? add_88795 : array_index_88245[0];
  assign array_update_89019[1] = add_85403 == 32'h0000_0001 ? add_88795 : array_index_88245[1];
  assign array_update_89019[2] = add_85403 == 32'h0000_0002 ? add_88795 : array_index_88245[2];
  assign array_update_89019[3] = add_85403 == 32'h0000_0003 ? add_88795 : array_index_88245[3];
  assign array_update_89019[4] = add_85403 == 32'h0000_0004 ? add_88795 : array_index_88245[4];
  assign array_update_89019[5] = add_85403 == 32'h0000_0005 ? add_88795 : array_index_88245[5];
  assign array_update_89019[6] = add_85403 == 32'h0000_0006 ? add_88795 : array_index_88245[6];
  assign array_update_89019[7] = add_85403 == 32'h0000_0007 ? add_88795 : array_index_88245[7];
  assign array_update_89019[8] = add_85403 == 32'h0000_0008 ? add_88795 : array_index_88245[8];
  assign array_update_89019[9] = add_85403 == 32'h0000_0009 ? add_88795 : array_index_88245[9];
  assign add_89020 = add_87719 + 32'h0000_0001;
  assign add_88772 = add_88448 + 32'h0000_0001;
  assign add_88774 = add_88450 + 32'h0000_0001;
  assign add_88776 = add_88452 + 32'h0000_0001;
  assign add_88778 = add_88454 + 32'h0000_0001;
  assign add_88780 = add_88456 + 32'h0000_0001;
  assign add_88782 = add_88458 + 32'h0000_0001;
  assign add_88784 = add_88460 + 32'h0000_0001;
  assign add_88786 = add_88462 + 32'h0000_0001;
  assign add_88788 = add_88464 + 32'h0000_0001;
  assign add_89017 = add_88792 + 32'h0000_0001;
  assign add_88790 = add_88466 + 32'h0000_0001;
  assign array_update_89343[0] = add_84176 == 32'h0000_0000 ? array_update_89019 : array_update_87920[0];
  assign array_update_89343[1] = add_84176 == 32'h0000_0001 ? array_update_89019 : array_update_87920[1];
  assign array_update_89343[2] = add_84176 == 32'h0000_0002 ? array_update_89019 : array_update_87920[2];
  assign array_update_89343[3] = add_84176 == 32'h0000_0003 ? array_update_89019 : array_update_87920[3];
  assign array_update_89343[4] = add_84176 == 32'h0000_0004 ? array_update_89019 : array_update_87920[4];
  assign array_update_89343[5] = add_84176 == 32'h0000_0005 ? array_update_89019 : array_update_87920[5];
  assign array_update_89343[6] = add_84176 == 32'h0000_0006 ? array_update_89019 : array_update_87920[6];
  assign array_update_89343[7] = add_84176 == 32'h0000_0007 ? array_update_89019 : array_update_87920[7];
  assign array_update_89343[8] = add_84176 == 32'h0000_0008 ? array_update_89019 : array_update_87920[8];
  assign array_update_89343[9] = add_84176 == 32'h0000_0009 ? array_update_89019 : array_update_87920[9];
  assign array_index_89345 = array_update_72021[add_89020 > 32'h0000_0009 ? 4'h9 : add_89020[3:0]];
  assign add_88997 = add_88772 + 32'h0000_0001;
  assign add_88999 = add_88774 + 32'h0000_0001;
  assign add_89001 = add_88776 + 32'h0000_0001;
  assign add_89003 = add_88778 + 32'h0000_0001;
  assign add_89005 = add_88780 + 32'h0000_0001;
  assign add_89007 = add_88782 + 32'h0000_0001;
  assign add_89009 = add_88784 + 32'h0000_0001;
  assign add_89011 = add_88786 + 32'h0000_0001;
  assign add_89013 = add_88788 + 32'h0000_0001;
  assign add_89341 = add_89017 + 32'h0000_0001;
  assign add_89015 = add_88790 + 32'h0000_0001;
  assign array_index_89572 = array_update_89343[add_84176 > 32'h0000_0009 ? 4'h9 : add_84176[3:0]];
  assign add_89321 = add_88997 + 32'h0000_0001;
  assign add_89323 = add_88999 + 32'h0000_0001;
  assign add_89325 = add_89001 + 32'h0000_0001;
  assign add_89327 = add_89003 + 32'h0000_0001;
  assign add_89329 = add_89005 + 32'h0000_0001;
  assign add_89331 = add_89007 + 32'h0000_0001;
  assign add_89333 = add_89009 + 32'h0000_0001;
  assign add_89335 = add_89011 + 32'h0000_0001;
  assign add_89337 = add_89013 + 32'h0000_0001;
  assign add_89566 = add_89341 + 32'h0000_0001;
  assign add_89339 = add_89015 + 32'h0000_0001;
  assign smul_89899 = smul32b_32b_x_32b(array_index_84183[add_89020 > 32'h0000_0009 ? 4'h9 : add_89020[3:0]], array_index_89345[add_85403 > 32'h0000_0009 ? 4'h9 : add_85403[3:0]]);
  assign add_89546 = add_89321 + 32'h0000_0001;
  assign add_89548 = add_89323 + 32'h0000_0001;
  assign add_89550 = add_89325 + 32'h0000_0001;
  assign add_89552 = add_89327 + 32'h0000_0001;
  assign add_89554 = add_89329 + 32'h0000_0001;
  assign add_89556 = add_89331 + 32'h0000_0001;
  assign add_89558 = add_89333 + 32'h0000_0001;
  assign add_89560 = add_89335 + 32'h0000_0001;
  assign add_89562 = add_89337 + 32'h0000_0001;
  assign add_89895 = add_89566 + 32'h0000_0001;
  assign add_89564 = add_89339 + 32'h0000_0001;
  assign add_90127 = array_index_89572[add_85403 > 32'h0000_0009 ? 4'h9 : add_85403[3:0]] + smul_89899;
  assign add_89875 = add_89546 + 32'h0000_0001;
  assign add_89877 = add_89548 + 32'h0000_0001;
  assign add_89879 = add_89550 + 32'h0000_0001;
  assign add_89881 = add_89552 + 32'h0000_0001;
  assign add_89883 = add_89554 + 32'h0000_0001;
  assign add_89885 = add_89556 + 32'h0000_0001;
  assign add_89887 = add_89558 + 32'h0000_0001;
  assign add_89889 = add_89560 + 32'h0000_0001;
  assign add_89891 = add_89562 + 32'h0000_0001;
  assign add_90120 = add_89895 + 32'h0000_0001;
  assign add_89893 = add_89564 + 32'h0000_0001;
  assign array_update_90451[0] = add_85403 == 32'h0000_0000 ? add_90127 : array_index_89572[0];
  assign array_update_90451[1] = add_85403 == 32'h0000_0001 ? add_90127 : array_index_89572[1];
  assign array_update_90451[2] = add_85403 == 32'h0000_0002 ? add_90127 : array_index_89572[2];
  assign array_update_90451[3] = add_85403 == 32'h0000_0003 ? add_90127 : array_index_89572[3];
  assign array_update_90451[4] = add_85403 == 32'h0000_0004 ? add_90127 : array_index_89572[4];
  assign array_update_90451[5] = add_85403 == 32'h0000_0005 ? add_90127 : array_index_89572[5];
  assign array_update_90451[6] = add_85403 == 32'h0000_0006 ? add_90127 : array_index_89572[6];
  assign array_update_90451[7] = add_85403 == 32'h0000_0007 ? add_90127 : array_index_89572[7];
  assign array_update_90451[8] = add_85403 == 32'h0000_0008 ? add_90127 : array_index_89572[8];
  assign array_update_90451[9] = add_85403 == 32'h0000_0009 ? add_90127 : array_index_89572[9];
  assign add_90100 = add_89875 + 32'h0000_0001;
  assign add_90102 = add_89877 + 32'h0000_0001;
  assign add_90104 = add_89879 + 32'h0000_0001;
  assign add_90106 = add_89881 + 32'h0000_0001;
  assign add_90108 = add_89883 + 32'h0000_0001;
  assign add_90110 = add_89885 + 32'h0000_0001;
  assign add_90112 = add_89887 + 32'h0000_0001;
  assign add_90114 = add_89889 + 32'h0000_0001;
  assign add_90116 = add_89891 + 32'h0000_0001;
  assign add_90448 = add_90120 + 32'h0000_0001;
  assign add_90118 = add_89893 + 32'h0000_0001;
  assign array_update_90811[0] = add_84176 == 32'h0000_0000 ? array_update_90451 : array_update_89343[0];
  assign array_update_90811[1] = add_84176 == 32'h0000_0001 ? array_update_90451 : array_update_89343[1];
  assign array_update_90811[2] = add_84176 == 32'h0000_0002 ? array_update_90451 : array_update_89343[2];
  assign array_update_90811[3] = add_84176 == 32'h0000_0003 ? array_update_90451 : array_update_89343[3];
  assign array_update_90811[4] = add_84176 == 32'h0000_0004 ? array_update_90451 : array_update_89343[4];
  assign array_update_90811[5] = add_84176 == 32'h0000_0005 ? array_update_90451 : array_update_89343[5];
  assign array_update_90811[6] = add_84176 == 32'h0000_0006 ? array_update_90451 : array_update_89343[6];
  assign array_update_90811[7] = add_84176 == 32'h0000_0007 ? array_update_90451 : array_update_89343[7];
  assign array_update_90811[8] = add_84176 == 32'h0000_0008 ? array_update_90451 : array_update_89343[8];
  assign array_update_90811[9] = add_84176 == 32'h0000_0009 ? array_update_90451 : array_update_89343[9];
  assign add_90428 = add_90100 + 32'h0000_0001;
  assign add_90430 = add_90102 + 32'h0000_0001;
  assign add_90432 = add_90104 + 32'h0000_0001;
  assign add_90434 = add_90106 + 32'h0000_0001;
  assign add_90436 = add_90108 + 32'h0000_0001;
  assign add_90438 = add_90110 + 32'h0000_0001;
  assign add_90440 = add_90112 + 32'h0000_0001;
  assign add_90442 = add_90114 + 32'h0000_0001;
  assign add_90444 = add_90116 + 32'h0000_0001;
  assign add_90805 = add_90448 + 32'h0000_0001;
  assign add_90446 = add_90118 + 32'h0000_0001;
  assign array_index_91514 = array_update_90811[literal_88243 > 32'h0000_0009 ? 4'h9 : literal_88243[3:0]];
  assign add_90785 = add_90428 + 32'h0000_0001;
  assign array_index_91524 = array_update_90811[add_88468 > 32'h0000_0009 ? 4'h9 : add_88468[3:0]];
  assign add_90787 = add_90430 + 32'h0000_0001;
  assign array_index_91534 = array_update_90811[add_88792 > 32'h0000_0009 ? 4'h9 : add_88792[3:0]];
  assign add_90789 = add_90432 + 32'h0000_0001;
  assign array_index_91544 = array_update_90811[add_89017 > 32'h0000_0009 ? 4'h9 : add_89017[3:0]];
  assign add_90791 = add_90434 + 32'h0000_0001;
  assign array_index_91554 = array_update_90811[add_89341 > 32'h0000_0009 ? 4'h9 : add_89341[3:0]];
  assign add_90793 = add_90436 + 32'h0000_0001;
  assign array_index_91564 = array_update_90811[add_89566 > 32'h0000_0009 ? 4'h9 : add_89566[3:0]];
  assign add_90795 = add_90438 + 32'h0000_0001;
  assign array_index_91574 = array_update_90811[add_89895 > 32'h0000_0009 ? 4'h9 : add_89895[3:0]];
  assign add_90797 = add_90440 + 32'h0000_0001;
  assign array_index_91584 = array_update_90811[add_90120 > 32'h0000_0009 ? 4'h9 : add_90120[3:0]];
  assign add_90799 = add_90442 + 32'h0000_0001;
  assign array_index_91594 = array_update_90811[add_90448 > 32'h0000_0009 ? 4'h9 : add_90448[3:0]];
  assign add_90801 = add_90444 + 32'h0000_0001;
  assign array_index_91604 = array_update_90811[add_90805 > 32'h0000_0009 ? 4'h9 : add_90805[3:0]];
  assign add_90803 = add_90446 + 32'h0000_0001;
  assign out = {1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, {array_index_91514[literal_88223 > 32'h0000_0009 ? 4'h9 : literal_88223[3:0]], 1'h1}, {array_index_91514[add_88448 > 32'h0000_0009 ? 4'h9 : add_88448[3:0]], 1'h1}, {array_index_91514[add_88772 > 32'h0000_0009 ? 4'h9 : add_88772[3:0]], 1'h1}, {array_index_91514[add_88997 > 32'h0000_0009 ? 4'h9 : add_88997[3:0]], 1'h1}, {array_index_91514[add_89321 > 32'h0000_0009 ? 4'h9 : add_89321[3:0]], 1'h1}, {array_index_91514[add_89546 > 32'h0000_0009 ? 4'h9 : add_89546[3:0]], 1'h1}, {array_index_91514[add_89875 > 32'h0000_0009 ? 4'h9 : add_89875[3:0]], 1'h1}, {array_index_91514[add_90100 > 32'h0000_0009 ? 4'h9 : add_90100[3:0]], 1'h1}, {array_index_91514[add_90428 > 32'h0000_0009 ? 4'h9 : add_90428[3:0]], 1'h1}, {array_index_91514[add_90785 > 32'h0000_0009 ? 4'h9 : add_90785[3:0]], 1'h1}, {array_index_91524[literal_88225 > 32'h0000_0009 ? 4'h9 : literal_88225[3:0]], 1'h1}, {array_index_91524[add_88450 > 32'h0000_0009 ? 4'h9 : add_88450[3:0]], 1'h1}, {array_index_91524[add_88774 > 32'h0000_0009 ? 4'h9 : add_88774[3:0]], 1'h1}, {array_index_91524[add_88999 > 32'h0000_0009 ? 4'h9 : add_88999[3:0]], 1'h1}, {array_index_91524[add_89323 > 32'h0000_0009 ? 4'h9 : add_89323[3:0]], 1'h1}, {array_index_91524[add_89548 > 32'h0000_0009 ? 4'h9 : add_89548[3:0]], 1'h1}, {array_index_91524[add_89877 > 32'h0000_0009 ? 4'h9 : add_89877[3:0]], 1'h1}, {array_index_91524[add_90102 > 32'h0000_0009 ? 4'h9 : add_90102[3:0]], 1'h1}, {array_index_91524[add_90430 > 32'h0000_0009 ? 4'h9 : add_90430[3:0]], 1'h1}, {array_index_91524[add_90787 > 32'h0000_0009 ? 4'h9 : add_90787[3:0]], 1'h1}, {array_index_91534[literal_88227 > 32'h0000_0009 ? 4'h9 : literal_88227[3:0]], 1'h1}, {array_index_91534[add_88452 > 32'h0000_0009 ? 4'h9 : add_88452[3:0]], 1'h1}, {array_index_91534[add_88776 > 32'h0000_0009 ? 4'h9 : add_88776[3:0]], 1'h1}, {array_index_91534[add_89001 > 32'h0000_0009 ? 4'h9 : add_89001[3:0]], 1'h1}, {array_index_91534[add_89325 > 32'h0000_0009 ? 4'h9 : add_89325[3:0]], 1'h1}, {array_index_91534[add_89550 > 32'h0000_0009 ? 4'h9 : add_89550[3:0]], 1'h1}, {array_index_91534[add_89879 > 32'h0000_0009 ? 4'h9 : add_89879[3:0]], 1'h1}, {array_index_91534[add_90104 > 32'h0000_0009 ? 4'h9 : add_90104[3:0]], 1'h1}, {array_index_91534[add_90432 > 32'h0000_0009 ? 4'h9 : add_90432[3:0]], 1'h1}, {array_index_91534[add_90789 > 32'h0000_0009 ? 4'h9 : add_90789[3:0]], 1'h1}, {array_index_91544[literal_88229 > 32'h0000_0009 ? 4'h9 : literal_88229[3:0]], 1'h1}, {array_index_91544[add_88454 > 32'h0000_0009 ? 4'h9 : add_88454[3:0]], 1'h1}, {array_index_91544[add_88778 > 32'h0000_0009 ? 4'h9 : add_88778[3:0]], 1'h1}, {array_index_91544[add_89003 > 32'h0000_0009 ? 4'h9 : add_89003[3:0]], 1'h1}, {array_index_91544[add_89327 > 32'h0000_0009 ? 4'h9 : add_89327[3:0]], 1'h1}, {array_index_91544[add_89552 > 32'h0000_0009 ? 4'h9 : add_89552[3:0]], 1'h1}, {array_index_91544[add_89881 > 32'h0000_0009 ? 4'h9 : add_89881[3:0]], 1'h1}, {array_index_91544[add_90106 > 32'h0000_0009 ? 4'h9 : add_90106[3:0]], 1'h1}, {array_index_91544[add_90434 > 32'h0000_0009 ? 4'h9 : add_90434[3:0]], 1'h1}, {array_index_91544[add_90791 > 32'h0000_0009 ? 4'h9 : add_90791[3:0]], 1'h1}, {array_index_91554[literal_88231 > 32'h0000_0009 ? 4'h9 : literal_88231[3:0]], 1'h1}, {array_index_91554[add_88456 > 32'h0000_0009 ? 4'h9 : add_88456[3:0]], 1'h1}, {array_index_91554[add_88780 > 32'h0000_0009 ? 4'h9 : add_88780[3:0]], 1'h1}, {array_index_91554[add_89005 > 32'h0000_0009 ? 4'h9 : add_89005[3:0]], 1'h1}, {array_index_91554[add_89329 > 32'h0000_0009 ? 4'h9 : add_89329[3:0]], 1'h1}, {array_index_91554[add_89554 > 32'h0000_0009 ? 4'h9 : add_89554[3:0]], 1'h1}, {array_index_91554[add_89883 > 32'h0000_0009 ? 4'h9 : add_89883[3:0]], 1'h1}, {array_index_91554[add_90108 > 32'h0000_0009 ? 4'h9 : add_90108[3:0]], 1'h1}, {array_index_91554[add_90436 > 32'h0000_0009 ? 4'h9 : add_90436[3:0]], 1'h1}, {array_index_91554[add_90793 > 32'h0000_0009 ? 4'h9 : add_90793[3:0]], 1'h1}, {array_index_91564[literal_88233 > 32'h0000_0009 ? 4'h9 : literal_88233[3:0]], 1'h1}, {array_index_91564[add_88458 > 32'h0000_0009 ? 4'h9 : add_88458[3:0]], 1'h1}, {array_index_91564[add_88782 > 32'h0000_0009 ? 4'h9 : add_88782[3:0]], 1'h1}, {array_index_91564[add_89007 > 32'h0000_0009 ? 4'h9 : add_89007[3:0]], 1'h1}, {array_index_91564[add_89331 > 32'h0000_0009 ? 4'h9 : add_89331[3:0]], 1'h1}, {array_index_91564[add_89556 > 32'h0000_0009 ? 4'h9 : add_89556[3:0]], 1'h1}, {array_index_91564[add_89885 > 32'h0000_0009 ? 4'h9 : add_89885[3:0]], 1'h1}, {array_index_91564[add_90110 > 32'h0000_0009 ? 4'h9 : add_90110[3:0]], 1'h1}, {array_index_91564[add_90438 > 32'h0000_0009 ? 4'h9 : add_90438[3:0]], 1'h1}, {array_index_91564[add_90795 > 32'h0000_0009 ? 4'h9 : add_90795[3:0]], 1'h1}, {array_index_91574[literal_88235 > 32'h0000_0009 ? 4'h9 : literal_88235[3:0]], 1'h1}, {array_index_91574[add_88460 > 32'h0000_0009 ? 4'h9 : add_88460[3:0]], 1'h1}, {array_index_91574[add_88784 > 32'h0000_0009 ? 4'h9 : add_88784[3:0]], 1'h1}, {array_index_91574[add_89009 > 32'h0000_0009 ? 4'h9 : add_89009[3:0]], 1'h1}, {array_index_91574[add_89333 > 32'h0000_0009 ? 4'h9 : add_89333[3:0]], 1'h1}, {array_index_91574[add_89558 > 32'h0000_0009 ? 4'h9 : add_89558[3:0]], 1'h1}, {array_index_91574[add_89887 > 32'h0000_0009 ? 4'h9 : add_89887[3:0]], 1'h1}, {array_index_91574[add_90112 > 32'h0000_0009 ? 4'h9 : add_90112[3:0]], 1'h1}, {array_index_91574[add_90440 > 32'h0000_0009 ? 4'h9 : add_90440[3:0]], 1'h1}, {array_index_91574[add_90797 > 32'h0000_0009 ? 4'h9 : add_90797[3:0]], 1'h1}, {array_index_91584[literal_88237 > 32'h0000_0009 ? 4'h9 : literal_88237[3:0]], 1'h1}, {array_index_91584[add_88462 > 32'h0000_0009 ? 4'h9 : add_88462[3:0]], 1'h1}, {array_index_91584[add_88786 > 32'h0000_0009 ? 4'h9 : add_88786[3:0]], 1'h1}, {array_index_91584[add_89011 > 32'h0000_0009 ? 4'h9 : add_89011[3:0]], 1'h1}, {array_index_91584[add_89335 > 32'h0000_0009 ? 4'h9 : add_89335[3:0]], 1'h1}, {array_index_91584[add_89560 > 32'h0000_0009 ? 4'h9 : add_89560[3:0]], 1'h1}, {array_index_91584[add_89889 > 32'h0000_0009 ? 4'h9 : add_89889[3:0]], 1'h1}, {array_index_91584[add_90114 > 32'h0000_0009 ? 4'h9 : add_90114[3:0]], 1'h1}, {array_index_91584[add_90442 > 32'h0000_0009 ? 4'h9 : add_90442[3:0]], 1'h1}, {array_index_91584[add_90799 > 32'h0000_0009 ? 4'h9 : add_90799[3:0]], 1'h1}, {array_index_91594[literal_88239 > 32'h0000_0009 ? 4'h9 : literal_88239[3:0]], 1'h1}, {array_index_91594[add_88464 > 32'h0000_0009 ? 4'h9 : add_88464[3:0]], 1'h1}, {array_index_91594[add_88788 > 32'h0000_0009 ? 4'h9 : add_88788[3:0]], 1'h1}, {array_index_91594[add_89013 > 32'h0000_0009 ? 4'h9 : add_89013[3:0]], 1'h1}, {array_index_91594[add_89337 > 32'h0000_0009 ? 4'h9 : add_89337[3:0]], 1'h1}, {array_index_91594[add_89562 > 32'h0000_0009 ? 4'h9 : add_89562[3:0]], 1'h1}, {array_index_91594[add_89891 > 32'h0000_0009 ? 4'h9 : add_89891[3:0]], 1'h1}, {array_index_91594[add_90116 > 32'h0000_0009 ? 4'h9 : add_90116[3:0]], 1'h1}, {array_index_91594[add_90444 > 32'h0000_0009 ? 4'h9 : add_90444[3:0]], 1'h1}, {array_index_91594[add_90801 > 32'h0000_0009 ? 4'h9 : add_90801[3:0]], 1'h1}, {array_index_91604[literal_88241 > 32'h0000_0009 ? 4'h9 : literal_88241[3:0]], 1'h1}, {array_index_91604[add_88466 > 32'h0000_0009 ? 4'h9 : add_88466[3:0]], 1'h1}, {array_index_91604[add_88790 > 32'h0000_0009 ? 4'h9 : add_88790[3:0]], 1'h1}, {array_index_91604[add_89015 > 32'h0000_0009 ? 4'h9 : add_89015[3:0]], 1'h1}, {array_index_91604[add_89339 > 32'h0000_0009 ? 4'h9 : add_89339[3:0]], 1'h1}, {array_index_91604[add_89564 > 32'h0000_0009 ? 4'h9 : add_89564[3:0]], 1'h1}, {array_index_91604[add_89893 > 32'h0000_0009 ? 4'h9 : add_89893[3:0]], 1'h1}, {array_index_91604[add_90118 > 32'h0000_0009 ? 4'h9 : add_90118[3:0]], 1'h1}, {array_index_91604[add_90446 > 32'h0000_0009 ? 4'h9 : add_90446[3:0]], 1'h1}, {array_index_91604[add_90803 > 32'h0000_0009 ? 4'h9 : add_90803[3:0]], 1'h1}};
endmodule
