module matrix_mul_10_pipeline(
  input wire clk,
  input wire [31:0] TestBlock__A_op0,
  input wire [31:0] TestBlock__A_op1,
  input wire [31:0] TestBlock__A_op2,
  input wire [31:0] TestBlock__A_op3,
  input wire [31:0] TestBlock__A_op4,
  input wire [31:0] TestBlock__A_op5,
  input wire [31:0] TestBlock__A_op6,
  input wire [31:0] TestBlock__A_op7,
  input wire [31:0] TestBlock__A_op8,
  input wire [31:0] TestBlock__A_op9,
  input wire [31:0] TestBlock__A_op10,
  input wire [31:0] TestBlock__A_op11,
  input wire [31:0] TestBlock__A_op12,
  input wire [31:0] TestBlock__A_op13,
  input wire [31:0] TestBlock__A_op14,
  input wire [31:0] TestBlock__A_op15,
  input wire [31:0] TestBlock__A_op16,
  input wire [31:0] TestBlock__A_op17,
  input wire [31:0] TestBlock__A_op18,
  input wire [31:0] TestBlock__A_op19,
  input wire [31:0] TestBlock__A_op20,
  input wire [31:0] TestBlock__A_op21,
  input wire [31:0] TestBlock__A_op22,
  input wire [31:0] TestBlock__A_op23,
  input wire [31:0] TestBlock__A_op24,
  input wire [31:0] TestBlock__A_op25,
  input wire [31:0] TestBlock__A_op26,
  input wire [31:0] TestBlock__A_op27,
  input wire [31:0] TestBlock__A_op28,
  input wire [31:0] TestBlock__A_op29,
  input wire [31:0] TestBlock__A_op30,
  input wire [31:0] TestBlock__A_op31,
  input wire [31:0] TestBlock__A_op32,
  input wire [31:0] TestBlock__A_op33,
  input wire [31:0] TestBlock__A_op34,
  input wire [31:0] TestBlock__A_op35,
  input wire [31:0] TestBlock__A_op36,
  input wire [31:0] TestBlock__A_op37,
  input wire [31:0] TestBlock__A_op38,
  input wire [31:0] TestBlock__A_op39,
  input wire [31:0] TestBlock__A_op40,
  input wire [31:0] TestBlock__A_op41,
  input wire [31:0] TestBlock__A_op42,
  input wire [31:0] TestBlock__A_op43,
  input wire [31:0] TestBlock__A_op44,
  input wire [31:0] TestBlock__A_op45,
  input wire [31:0] TestBlock__A_op46,
  input wire [31:0] TestBlock__A_op47,
  input wire [31:0] TestBlock__A_op48,
  input wire [31:0] TestBlock__A_op49,
  input wire [31:0] TestBlock__A_op50,
  input wire [31:0] TestBlock__A_op51,
  input wire [31:0] TestBlock__A_op52,
  input wire [31:0] TestBlock__A_op53,
  input wire [31:0] TestBlock__A_op54,
  input wire [31:0] TestBlock__A_op55,
  input wire [31:0] TestBlock__A_op56,
  input wire [31:0] TestBlock__A_op57,
  input wire [31:0] TestBlock__A_op58,
  input wire [31:0] TestBlock__A_op59,
  input wire [31:0] TestBlock__A_op60,
  input wire [31:0] TestBlock__A_op61,
  input wire [31:0] TestBlock__A_op62,
  input wire [31:0] TestBlock__A_op63,
  input wire [31:0] TestBlock__A_op64,
  input wire [31:0] TestBlock__A_op65,
  input wire [31:0] TestBlock__A_op66,
  input wire [31:0] TestBlock__A_op67,
  input wire [31:0] TestBlock__A_op68,
  input wire [31:0] TestBlock__A_op69,
  input wire [31:0] TestBlock__A_op70,
  input wire [31:0] TestBlock__A_op71,
  input wire [31:0] TestBlock__A_op72,
  input wire [31:0] TestBlock__A_op73,
  input wire [31:0] TestBlock__A_op74,
  input wire [31:0] TestBlock__A_op75,
  input wire [31:0] TestBlock__A_op76,
  input wire [31:0] TestBlock__A_op77,
  input wire [31:0] TestBlock__A_op78,
  input wire [31:0] TestBlock__A_op79,
  input wire [31:0] TestBlock__A_op80,
  input wire [31:0] TestBlock__A_op81,
  input wire [31:0] TestBlock__A_op82,
  input wire [31:0] TestBlock__A_op83,
  input wire [31:0] TestBlock__A_op84,
  input wire [31:0] TestBlock__A_op85,
  input wire [31:0] TestBlock__A_op86,
  input wire [31:0] TestBlock__A_op87,
  input wire [31:0] TestBlock__A_op88,
  input wire [31:0] TestBlock__A_op89,
  input wire [31:0] TestBlock__A_op90,
  input wire [31:0] TestBlock__A_op91,
  input wire [31:0] TestBlock__A_op92,
  input wire [31:0] TestBlock__A_op93,
  input wire [31:0] TestBlock__A_op94,
  input wire [31:0] TestBlock__A_op95,
  input wire [31:0] TestBlock__A_op96,
  input wire [31:0] TestBlock__A_op97,
  input wire [31:0] TestBlock__A_op98,
  input wire [31:0] TestBlock__A_op99,
  input wire [31:0] TestBlock__B_op0,
  input wire [31:0] TestBlock__B_op1,
  input wire [31:0] TestBlock__B_op2,
  input wire [31:0] TestBlock__B_op3,
  input wire [31:0] TestBlock__B_op4,
  input wire [31:0] TestBlock__B_op5,
  input wire [31:0] TestBlock__B_op6,
  input wire [31:0] TestBlock__B_op7,
  input wire [31:0] TestBlock__B_op8,
  input wire [31:0] TestBlock__B_op9,
  input wire [31:0] TestBlock__B_op10,
  input wire [31:0] TestBlock__B_op11,
  input wire [31:0] TestBlock__B_op12,
  input wire [31:0] TestBlock__B_op13,
  input wire [31:0] TestBlock__B_op14,
  input wire [31:0] TestBlock__B_op15,
  input wire [31:0] TestBlock__B_op16,
  input wire [31:0] TestBlock__B_op17,
  input wire [31:0] TestBlock__B_op18,
  input wire [31:0] TestBlock__B_op19,
  input wire [31:0] TestBlock__B_op20,
  input wire [31:0] TestBlock__B_op21,
  input wire [31:0] TestBlock__B_op22,
  input wire [31:0] TestBlock__B_op23,
  input wire [31:0] TestBlock__B_op24,
  input wire [31:0] TestBlock__B_op25,
  input wire [31:0] TestBlock__B_op26,
  input wire [31:0] TestBlock__B_op27,
  input wire [31:0] TestBlock__B_op28,
  input wire [31:0] TestBlock__B_op29,
  input wire [31:0] TestBlock__B_op30,
  input wire [31:0] TestBlock__B_op31,
  input wire [31:0] TestBlock__B_op32,
  input wire [31:0] TestBlock__B_op33,
  input wire [31:0] TestBlock__B_op34,
  input wire [31:0] TestBlock__B_op35,
  input wire [31:0] TestBlock__B_op36,
  input wire [31:0] TestBlock__B_op37,
  input wire [31:0] TestBlock__B_op38,
  input wire [31:0] TestBlock__B_op39,
  input wire [31:0] TestBlock__B_op40,
  input wire [31:0] TestBlock__B_op41,
  input wire [31:0] TestBlock__B_op42,
  input wire [31:0] TestBlock__B_op43,
  input wire [31:0] TestBlock__B_op44,
  input wire [31:0] TestBlock__B_op45,
  input wire [31:0] TestBlock__B_op46,
  input wire [31:0] TestBlock__B_op47,
  input wire [31:0] TestBlock__B_op48,
  input wire [31:0] TestBlock__B_op49,
  input wire [31:0] TestBlock__B_op50,
  input wire [31:0] TestBlock__B_op51,
  input wire [31:0] TestBlock__B_op52,
  input wire [31:0] TestBlock__B_op53,
  input wire [31:0] TestBlock__B_op54,
  input wire [31:0] TestBlock__B_op55,
  input wire [31:0] TestBlock__B_op56,
  input wire [31:0] TestBlock__B_op57,
  input wire [31:0] TestBlock__B_op58,
  input wire [31:0] TestBlock__B_op59,
  input wire [31:0] TestBlock__B_op60,
  input wire [31:0] TestBlock__B_op61,
  input wire [31:0] TestBlock__B_op62,
  input wire [31:0] TestBlock__B_op63,
  input wire [31:0] TestBlock__B_op64,
  input wire [31:0] TestBlock__B_op65,
  input wire [31:0] TestBlock__B_op66,
  input wire [31:0] TestBlock__B_op67,
  input wire [31:0] TestBlock__B_op68,
  input wire [31:0] TestBlock__B_op69,
  input wire [31:0] TestBlock__B_op70,
  input wire [31:0] TestBlock__B_op71,
  input wire [31:0] TestBlock__B_op72,
  input wire [31:0] TestBlock__B_op73,
  input wire [31:0] TestBlock__B_op74,
  input wire [31:0] TestBlock__B_op75,
  input wire [31:0] TestBlock__B_op76,
  input wire [31:0] TestBlock__B_op77,
  input wire [31:0] TestBlock__B_op78,
  input wire [31:0] TestBlock__B_op79,
  input wire [31:0] TestBlock__B_op80,
  input wire [31:0] TestBlock__B_op81,
  input wire [31:0] TestBlock__B_op82,
  input wire [31:0] TestBlock__B_op83,
  input wire [31:0] TestBlock__B_op84,
  input wire [31:0] TestBlock__B_op85,
  input wire [31:0] TestBlock__B_op86,
  input wire [31:0] TestBlock__B_op87,
  input wire [31:0] TestBlock__B_op88,
  input wire [31:0] TestBlock__B_op89,
  input wire [31:0] TestBlock__B_op90,
  input wire [31:0] TestBlock__B_op91,
  input wire [31:0] TestBlock__B_op92,
  input wire [31:0] TestBlock__B_op93,
  input wire [31:0] TestBlock__B_op94,
  input wire [31:0] TestBlock__B_op95,
  input wire [31:0] TestBlock__B_op96,
  input wire [31:0] TestBlock__B_op97,
  input wire [31:0] TestBlock__B_op98,
  input wire [31:0] TestBlock__B_op99,
  output wire [3499:0] out
);
  // lint_off SIGNED_TYPE
  // lint_off MULTIPLY
  function automatic [31:0] smul32b_32b_x_32b (input reg [31:0] lhs, input reg [31:0] rhs);
    reg signed [31:0] signed_lhs;
    reg signed [31:0] signed_rhs;
    reg signed [31:0] signed_result;
    begin
      signed_lhs = $signed(lhs);
      signed_rhs = $signed(rhs);
      signed_result = signed_lhs * signed_rhs;
      smul32b_32b_x_32b = $unsigned(signed_result);
    end
  endfunction
  // lint_on MULTIPLY
  // lint_on SIGNED_TYPE

  // ===== Pipe stage 0:

  // Registers for pipe stage 0:
  reg [31:0] p0_TestBlock__A_op0;
  reg [31:0] p0_TestBlock__A_op1;
  reg [31:0] p0_TestBlock__A_op2;
  reg [31:0] p0_TestBlock__A_op3;
  reg [31:0] p0_TestBlock__A_op4;
  reg [31:0] p0_TestBlock__A_op5;
  reg [31:0] p0_TestBlock__A_op6;
  reg [31:0] p0_TestBlock__A_op7;
  reg [31:0] p0_TestBlock__A_op8;
  reg [31:0] p0_TestBlock__A_op9;
  reg [31:0] p0_TestBlock__A_op10;
  reg [31:0] p0_TestBlock__A_op11;
  reg [31:0] p0_TestBlock__A_op12;
  reg [31:0] p0_TestBlock__A_op13;
  reg [31:0] p0_TestBlock__A_op14;
  reg [31:0] p0_TestBlock__A_op15;
  reg [31:0] p0_TestBlock__A_op16;
  reg [31:0] p0_TestBlock__A_op17;
  reg [31:0] p0_TestBlock__A_op18;
  reg [31:0] p0_TestBlock__A_op19;
  reg [31:0] p0_TestBlock__A_op20;
  reg [31:0] p0_TestBlock__A_op21;
  reg [31:0] p0_TestBlock__A_op22;
  reg [31:0] p0_TestBlock__A_op23;
  reg [31:0] p0_TestBlock__A_op24;
  reg [31:0] p0_TestBlock__A_op25;
  reg [31:0] p0_TestBlock__A_op26;
  reg [31:0] p0_TestBlock__A_op27;
  reg [31:0] p0_TestBlock__A_op28;
  reg [31:0] p0_TestBlock__A_op29;
  reg [31:0] p0_TestBlock__A_op30;
  reg [31:0] p0_TestBlock__A_op31;
  reg [31:0] p0_TestBlock__A_op32;
  reg [31:0] p0_TestBlock__A_op33;
  reg [31:0] p0_TestBlock__A_op34;
  reg [31:0] p0_TestBlock__A_op35;
  reg [31:0] p0_TestBlock__A_op36;
  reg [31:0] p0_TestBlock__A_op37;
  reg [31:0] p0_TestBlock__A_op38;
  reg [31:0] p0_TestBlock__A_op39;
  reg [31:0] p0_TestBlock__A_op40;
  reg [31:0] p0_TestBlock__A_op41;
  reg [31:0] p0_TestBlock__A_op42;
  reg [31:0] p0_TestBlock__A_op43;
  reg [31:0] p0_TestBlock__A_op44;
  reg [31:0] p0_TestBlock__A_op45;
  reg [31:0] p0_TestBlock__A_op46;
  reg [31:0] p0_TestBlock__A_op47;
  reg [31:0] p0_TestBlock__A_op48;
  reg [31:0] p0_TestBlock__A_op49;
  reg [31:0] p0_TestBlock__A_op50;
  reg [31:0] p0_TestBlock__A_op51;
  reg [31:0] p0_TestBlock__A_op52;
  reg [31:0] p0_TestBlock__A_op53;
  reg [31:0] p0_TestBlock__A_op54;
  reg [31:0] p0_TestBlock__A_op55;
  reg [31:0] p0_TestBlock__A_op56;
  reg [31:0] p0_TestBlock__A_op57;
  reg [31:0] p0_TestBlock__A_op58;
  reg [31:0] p0_TestBlock__A_op59;
  reg [31:0] p0_TestBlock__A_op60;
  reg [31:0] p0_TestBlock__A_op61;
  reg [31:0] p0_TestBlock__A_op62;
  reg [31:0] p0_TestBlock__A_op63;
  reg [31:0] p0_TestBlock__A_op64;
  reg [31:0] p0_TestBlock__A_op65;
  reg [31:0] p0_TestBlock__A_op66;
  reg [31:0] p0_TestBlock__A_op67;
  reg [31:0] p0_TestBlock__A_op68;
  reg [31:0] p0_TestBlock__A_op69;
  reg [31:0] p0_TestBlock__A_op70;
  reg [31:0] p0_TestBlock__A_op71;
  reg [31:0] p0_TestBlock__A_op72;
  reg [31:0] p0_TestBlock__A_op73;
  reg [31:0] p0_TestBlock__A_op74;
  reg [31:0] p0_TestBlock__A_op75;
  reg [31:0] p0_TestBlock__A_op76;
  reg [31:0] p0_TestBlock__A_op77;
  reg [31:0] p0_TestBlock__A_op78;
  reg [31:0] p0_TestBlock__A_op79;
  reg [31:0] p0_TestBlock__A_op80;
  reg [31:0] p0_TestBlock__A_op81;
  reg [31:0] p0_TestBlock__A_op82;
  reg [31:0] p0_TestBlock__A_op83;
  reg [31:0] p0_TestBlock__A_op84;
  reg [31:0] p0_TestBlock__A_op85;
  reg [31:0] p0_TestBlock__A_op86;
  reg [31:0] p0_TestBlock__A_op87;
  reg [31:0] p0_TestBlock__A_op88;
  reg [31:0] p0_TestBlock__A_op89;
  reg [31:0] p0_TestBlock__A_op90;
  reg [31:0] p0_TestBlock__A_op91;
  reg [31:0] p0_TestBlock__A_op92;
  reg [31:0] p0_TestBlock__A_op93;
  reg [31:0] p0_TestBlock__A_op94;
  reg [31:0] p0_TestBlock__A_op95;
  reg [31:0] p0_TestBlock__A_op96;
  reg [31:0] p0_TestBlock__A_op97;
  reg [31:0] p0_TestBlock__A_op98;
  reg [31:0] p0_TestBlock__A_op99;
  reg [31:0] p0_TestBlock__B_op0;
  reg [31:0] p0_TestBlock__B_op1;
  reg [31:0] p0_TestBlock__B_op2;
  reg [31:0] p0_TestBlock__B_op3;
  reg [31:0] p0_TestBlock__B_op4;
  reg [31:0] p0_TestBlock__B_op5;
  reg [31:0] p0_TestBlock__B_op6;
  reg [31:0] p0_TestBlock__B_op7;
  reg [31:0] p0_TestBlock__B_op8;
  reg [31:0] p0_TestBlock__B_op9;
  reg [31:0] p0_TestBlock__B_op10;
  reg [31:0] p0_TestBlock__B_op11;
  reg [31:0] p0_TestBlock__B_op12;
  reg [31:0] p0_TestBlock__B_op13;
  reg [31:0] p0_TestBlock__B_op14;
  reg [31:0] p0_TestBlock__B_op15;
  reg [31:0] p0_TestBlock__B_op16;
  reg [31:0] p0_TestBlock__B_op17;
  reg [31:0] p0_TestBlock__B_op18;
  reg [31:0] p0_TestBlock__B_op19;
  reg [31:0] p0_TestBlock__B_op20;
  reg [31:0] p0_TestBlock__B_op21;
  reg [31:0] p0_TestBlock__B_op22;
  reg [31:0] p0_TestBlock__B_op23;
  reg [31:0] p0_TestBlock__B_op24;
  reg [31:0] p0_TestBlock__B_op25;
  reg [31:0] p0_TestBlock__B_op26;
  reg [31:0] p0_TestBlock__B_op27;
  reg [31:0] p0_TestBlock__B_op28;
  reg [31:0] p0_TestBlock__B_op29;
  reg [31:0] p0_TestBlock__B_op30;
  reg [31:0] p0_TestBlock__B_op31;
  reg [31:0] p0_TestBlock__B_op32;
  reg [31:0] p0_TestBlock__B_op33;
  reg [31:0] p0_TestBlock__B_op34;
  reg [31:0] p0_TestBlock__B_op35;
  reg [31:0] p0_TestBlock__B_op36;
  reg [31:0] p0_TestBlock__B_op37;
  reg [31:0] p0_TestBlock__B_op38;
  reg [31:0] p0_TestBlock__B_op39;
  reg [31:0] p0_TestBlock__B_op40;
  reg [31:0] p0_TestBlock__B_op41;
  reg [31:0] p0_TestBlock__B_op42;
  reg [31:0] p0_TestBlock__B_op43;
  reg [31:0] p0_TestBlock__B_op44;
  reg [31:0] p0_TestBlock__B_op45;
  reg [31:0] p0_TestBlock__B_op46;
  reg [31:0] p0_TestBlock__B_op47;
  reg [31:0] p0_TestBlock__B_op48;
  reg [31:0] p0_TestBlock__B_op49;
  reg [31:0] p0_TestBlock__B_op50;
  reg [31:0] p0_TestBlock__B_op51;
  reg [31:0] p0_TestBlock__B_op52;
  reg [31:0] p0_TestBlock__B_op53;
  reg [31:0] p0_TestBlock__B_op54;
  reg [31:0] p0_TestBlock__B_op55;
  reg [31:0] p0_TestBlock__B_op56;
  reg [31:0] p0_TestBlock__B_op57;
  reg [31:0] p0_TestBlock__B_op58;
  reg [31:0] p0_TestBlock__B_op59;
  reg [31:0] p0_TestBlock__B_op60;
  reg [31:0] p0_TestBlock__B_op61;
  reg [31:0] p0_TestBlock__B_op62;
  reg [31:0] p0_TestBlock__B_op63;
  reg [31:0] p0_TestBlock__B_op64;
  reg [31:0] p0_TestBlock__B_op65;
  reg [31:0] p0_TestBlock__B_op66;
  reg [31:0] p0_TestBlock__B_op67;
  reg [31:0] p0_TestBlock__B_op68;
  reg [31:0] p0_TestBlock__B_op69;
  reg [31:0] p0_TestBlock__B_op70;
  reg [31:0] p0_TestBlock__B_op71;
  reg [31:0] p0_TestBlock__B_op72;
  reg [31:0] p0_TestBlock__B_op73;
  reg [31:0] p0_TestBlock__B_op74;
  reg [31:0] p0_TestBlock__B_op75;
  reg [31:0] p0_TestBlock__B_op76;
  reg [31:0] p0_TestBlock__B_op77;
  reg [31:0] p0_TestBlock__B_op78;
  reg [31:0] p0_TestBlock__B_op79;
  reg [31:0] p0_TestBlock__B_op80;
  reg [31:0] p0_TestBlock__B_op81;
  reg [31:0] p0_TestBlock__B_op82;
  reg [31:0] p0_TestBlock__B_op83;
  reg [31:0] p0_TestBlock__B_op84;
  reg [31:0] p0_TestBlock__B_op85;
  reg [31:0] p0_TestBlock__B_op86;
  reg [31:0] p0_TestBlock__B_op87;
  reg [31:0] p0_TestBlock__B_op88;
  reg [31:0] p0_TestBlock__B_op89;
  reg [31:0] p0_TestBlock__B_op90;
  reg [31:0] p0_TestBlock__B_op91;
  reg [31:0] p0_TestBlock__B_op92;
  reg [31:0] p0_TestBlock__B_op93;
  reg [31:0] p0_TestBlock__B_op94;
  reg [31:0] p0_TestBlock__B_op95;
  reg [31:0] p0_TestBlock__B_op96;
  reg [31:0] p0_TestBlock__B_op97;
  reg [31:0] p0_TestBlock__B_op98;
  reg [31:0] p0_TestBlock__B_op99;
  always_ff @ (posedge clk) begin
    p0_TestBlock__A_op0 <= TestBlock__A_op0;
    p0_TestBlock__A_op1 <= TestBlock__A_op1;
    p0_TestBlock__A_op2 <= TestBlock__A_op2;
    p0_TestBlock__A_op3 <= TestBlock__A_op3;
    p0_TestBlock__A_op4 <= TestBlock__A_op4;
    p0_TestBlock__A_op5 <= TestBlock__A_op5;
    p0_TestBlock__A_op6 <= TestBlock__A_op6;
    p0_TestBlock__A_op7 <= TestBlock__A_op7;
    p0_TestBlock__A_op8 <= TestBlock__A_op8;
    p0_TestBlock__A_op9 <= TestBlock__A_op9;
    p0_TestBlock__A_op10 <= TestBlock__A_op10;
    p0_TestBlock__A_op11 <= TestBlock__A_op11;
    p0_TestBlock__A_op12 <= TestBlock__A_op12;
    p0_TestBlock__A_op13 <= TestBlock__A_op13;
    p0_TestBlock__A_op14 <= TestBlock__A_op14;
    p0_TestBlock__A_op15 <= TestBlock__A_op15;
    p0_TestBlock__A_op16 <= TestBlock__A_op16;
    p0_TestBlock__A_op17 <= TestBlock__A_op17;
    p0_TestBlock__A_op18 <= TestBlock__A_op18;
    p0_TestBlock__A_op19 <= TestBlock__A_op19;
    p0_TestBlock__A_op20 <= TestBlock__A_op20;
    p0_TestBlock__A_op21 <= TestBlock__A_op21;
    p0_TestBlock__A_op22 <= TestBlock__A_op22;
    p0_TestBlock__A_op23 <= TestBlock__A_op23;
    p0_TestBlock__A_op24 <= TestBlock__A_op24;
    p0_TestBlock__A_op25 <= TestBlock__A_op25;
    p0_TestBlock__A_op26 <= TestBlock__A_op26;
    p0_TestBlock__A_op27 <= TestBlock__A_op27;
    p0_TestBlock__A_op28 <= TestBlock__A_op28;
    p0_TestBlock__A_op29 <= TestBlock__A_op29;
    p0_TestBlock__A_op30 <= TestBlock__A_op30;
    p0_TestBlock__A_op31 <= TestBlock__A_op31;
    p0_TestBlock__A_op32 <= TestBlock__A_op32;
    p0_TestBlock__A_op33 <= TestBlock__A_op33;
    p0_TestBlock__A_op34 <= TestBlock__A_op34;
    p0_TestBlock__A_op35 <= TestBlock__A_op35;
    p0_TestBlock__A_op36 <= TestBlock__A_op36;
    p0_TestBlock__A_op37 <= TestBlock__A_op37;
    p0_TestBlock__A_op38 <= TestBlock__A_op38;
    p0_TestBlock__A_op39 <= TestBlock__A_op39;
    p0_TestBlock__A_op40 <= TestBlock__A_op40;
    p0_TestBlock__A_op41 <= TestBlock__A_op41;
    p0_TestBlock__A_op42 <= TestBlock__A_op42;
    p0_TestBlock__A_op43 <= TestBlock__A_op43;
    p0_TestBlock__A_op44 <= TestBlock__A_op44;
    p0_TestBlock__A_op45 <= TestBlock__A_op45;
    p0_TestBlock__A_op46 <= TestBlock__A_op46;
    p0_TestBlock__A_op47 <= TestBlock__A_op47;
    p0_TestBlock__A_op48 <= TestBlock__A_op48;
    p0_TestBlock__A_op49 <= TestBlock__A_op49;
    p0_TestBlock__A_op50 <= TestBlock__A_op50;
    p0_TestBlock__A_op51 <= TestBlock__A_op51;
    p0_TestBlock__A_op52 <= TestBlock__A_op52;
    p0_TestBlock__A_op53 <= TestBlock__A_op53;
    p0_TestBlock__A_op54 <= TestBlock__A_op54;
    p0_TestBlock__A_op55 <= TestBlock__A_op55;
    p0_TestBlock__A_op56 <= TestBlock__A_op56;
    p0_TestBlock__A_op57 <= TestBlock__A_op57;
    p0_TestBlock__A_op58 <= TestBlock__A_op58;
    p0_TestBlock__A_op59 <= TestBlock__A_op59;
    p0_TestBlock__A_op60 <= TestBlock__A_op60;
    p0_TestBlock__A_op61 <= TestBlock__A_op61;
    p0_TestBlock__A_op62 <= TestBlock__A_op62;
    p0_TestBlock__A_op63 <= TestBlock__A_op63;
    p0_TestBlock__A_op64 <= TestBlock__A_op64;
    p0_TestBlock__A_op65 <= TestBlock__A_op65;
    p0_TestBlock__A_op66 <= TestBlock__A_op66;
    p0_TestBlock__A_op67 <= TestBlock__A_op67;
    p0_TestBlock__A_op68 <= TestBlock__A_op68;
    p0_TestBlock__A_op69 <= TestBlock__A_op69;
    p0_TestBlock__A_op70 <= TestBlock__A_op70;
    p0_TestBlock__A_op71 <= TestBlock__A_op71;
    p0_TestBlock__A_op72 <= TestBlock__A_op72;
    p0_TestBlock__A_op73 <= TestBlock__A_op73;
    p0_TestBlock__A_op74 <= TestBlock__A_op74;
    p0_TestBlock__A_op75 <= TestBlock__A_op75;
    p0_TestBlock__A_op76 <= TestBlock__A_op76;
    p0_TestBlock__A_op77 <= TestBlock__A_op77;
    p0_TestBlock__A_op78 <= TestBlock__A_op78;
    p0_TestBlock__A_op79 <= TestBlock__A_op79;
    p0_TestBlock__A_op80 <= TestBlock__A_op80;
    p0_TestBlock__A_op81 <= TestBlock__A_op81;
    p0_TestBlock__A_op82 <= TestBlock__A_op82;
    p0_TestBlock__A_op83 <= TestBlock__A_op83;
    p0_TestBlock__A_op84 <= TestBlock__A_op84;
    p0_TestBlock__A_op85 <= TestBlock__A_op85;
    p0_TestBlock__A_op86 <= TestBlock__A_op86;
    p0_TestBlock__A_op87 <= TestBlock__A_op87;
    p0_TestBlock__A_op88 <= TestBlock__A_op88;
    p0_TestBlock__A_op89 <= TestBlock__A_op89;
    p0_TestBlock__A_op90 <= TestBlock__A_op90;
    p0_TestBlock__A_op91 <= TestBlock__A_op91;
    p0_TestBlock__A_op92 <= TestBlock__A_op92;
    p0_TestBlock__A_op93 <= TestBlock__A_op93;
    p0_TestBlock__A_op94 <= TestBlock__A_op94;
    p0_TestBlock__A_op95 <= TestBlock__A_op95;
    p0_TestBlock__A_op96 <= TestBlock__A_op96;
    p0_TestBlock__A_op97 <= TestBlock__A_op97;
    p0_TestBlock__A_op98 <= TestBlock__A_op98;
    p0_TestBlock__A_op99 <= TestBlock__A_op99;
    p0_TestBlock__B_op0 <= TestBlock__B_op0;
    p0_TestBlock__B_op1 <= TestBlock__B_op1;
    p0_TestBlock__B_op2 <= TestBlock__B_op2;
    p0_TestBlock__B_op3 <= TestBlock__B_op3;
    p0_TestBlock__B_op4 <= TestBlock__B_op4;
    p0_TestBlock__B_op5 <= TestBlock__B_op5;
    p0_TestBlock__B_op6 <= TestBlock__B_op6;
    p0_TestBlock__B_op7 <= TestBlock__B_op7;
    p0_TestBlock__B_op8 <= TestBlock__B_op8;
    p0_TestBlock__B_op9 <= TestBlock__B_op9;
    p0_TestBlock__B_op10 <= TestBlock__B_op10;
    p0_TestBlock__B_op11 <= TestBlock__B_op11;
    p0_TestBlock__B_op12 <= TestBlock__B_op12;
    p0_TestBlock__B_op13 <= TestBlock__B_op13;
    p0_TestBlock__B_op14 <= TestBlock__B_op14;
    p0_TestBlock__B_op15 <= TestBlock__B_op15;
    p0_TestBlock__B_op16 <= TestBlock__B_op16;
    p0_TestBlock__B_op17 <= TestBlock__B_op17;
    p0_TestBlock__B_op18 <= TestBlock__B_op18;
    p0_TestBlock__B_op19 <= TestBlock__B_op19;
    p0_TestBlock__B_op20 <= TestBlock__B_op20;
    p0_TestBlock__B_op21 <= TestBlock__B_op21;
    p0_TestBlock__B_op22 <= TestBlock__B_op22;
    p0_TestBlock__B_op23 <= TestBlock__B_op23;
    p0_TestBlock__B_op24 <= TestBlock__B_op24;
    p0_TestBlock__B_op25 <= TestBlock__B_op25;
    p0_TestBlock__B_op26 <= TestBlock__B_op26;
    p0_TestBlock__B_op27 <= TestBlock__B_op27;
    p0_TestBlock__B_op28 <= TestBlock__B_op28;
    p0_TestBlock__B_op29 <= TestBlock__B_op29;
    p0_TestBlock__B_op30 <= TestBlock__B_op30;
    p0_TestBlock__B_op31 <= TestBlock__B_op31;
    p0_TestBlock__B_op32 <= TestBlock__B_op32;
    p0_TestBlock__B_op33 <= TestBlock__B_op33;
    p0_TestBlock__B_op34 <= TestBlock__B_op34;
    p0_TestBlock__B_op35 <= TestBlock__B_op35;
    p0_TestBlock__B_op36 <= TestBlock__B_op36;
    p0_TestBlock__B_op37 <= TestBlock__B_op37;
    p0_TestBlock__B_op38 <= TestBlock__B_op38;
    p0_TestBlock__B_op39 <= TestBlock__B_op39;
    p0_TestBlock__B_op40 <= TestBlock__B_op40;
    p0_TestBlock__B_op41 <= TestBlock__B_op41;
    p0_TestBlock__B_op42 <= TestBlock__B_op42;
    p0_TestBlock__B_op43 <= TestBlock__B_op43;
    p0_TestBlock__B_op44 <= TestBlock__B_op44;
    p0_TestBlock__B_op45 <= TestBlock__B_op45;
    p0_TestBlock__B_op46 <= TestBlock__B_op46;
    p0_TestBlock__B_op47 <= TestBlock__B_op47;
    p0_TestBlock__B_op48 <= TestBlock__B_op48;
    p0_TestBlock__B_op49 <= TestBlock__B_op49;
    p0_TestBlock__B_op50 <= TestBlock__B_op50;
    p0_TestBlock__B_op51 <= TestBlock__B_op51;
    p0_TestBlock__B_op52 <= TestBlock__B_op52;
    p0_TestBlock__B_op53 <= TestBlock__B_op53;
    p0_TestBlock__B_op54 <= TestBlock__B_op54;
    p0_TestBlock__B_op55 <= TestBlock__B_op55;
    p0_TestBlock__B_op56 <= TestBlock__B_op56;
    p0_TestBlock__B_op57 <= TestBlock__B_op57;
    p0_TestBlock__B_op58 <= TestBlock__B_op58;
    p0_TestBlock__B_op59 <= TestBlock__B_op59;
    p0_TestBlock__B_op60 <= TestBlock__B_op60;
    p0_TestBlock__B_op61 <= TestBlock__B_op61;
    p0_TestBlock__B_op62 <= TestBlock__B_op62;
    p0_TestBlock__B_op63 <= TestBlock__B_op63;
    p0_TestBlock__B_op64 <= TestBlock__B_op64;
    p0_TestBlock__B_op65 <= TestBlock__B_op65;
    p0_TestBlock__B_op66 <= TestBlock__B_op66;
    p0_TestBlock__B_op67 <= TestBlock__B_op67;
    p0_TestBlock__B_op68 <= TestBlock__B_op68;
    p0_TestBlock__B_op69 <= TestBlock__B_op69;
    p0_TestBlock__B_op70 <= TestBlock__B_op70;
    p0_TestBlock__B_op71 <= TestBlock__B_op71;
    p0_TestBlock__B_op72 <= TestBlock__B_op72;
    p0_TestBlock__B_op73 <= TestBlock__B_op73;
    p0_TestBlock__B_op74 <= TestBlock__B_op74;
    p0_TestBlock__B_op75 <= TestBlock__B_op75;
    p0_TestBlock__B_op76 <= TestBlock__B_op76;
    p0_TestBlock__B_op77 <= TestBlock__B_op77;
    p0_TestBlock__B_op78 <= TestBlock__B_op78;
    p0_TestBlock__B_op79 <= TestBlock__B_op79;
    p0_TestBlock__B_op80 <= TestBlock__B_op80;
    p0_TestBlock__B_op81 <= TestBlock__B_op81;
    p0_TestBlock__B_op82 <= TestBlock__B_op82;
    p0_TestBlock__B_op83 <= TestBlock__B_op83;
    p0_TestBlock__B_op84 <= TestBlock__B_op84;
    p0_TestBlock__B_op85 <= TestBlock__B_op85;
    p0_TestBlock__B_op86 <= TestBlock__B_op86;
    p0_TestBlock__B_op87 <= TestBlock__B_op87;
    p0_TestBlock__B_op88 <= TestBlock__B_op88;
    p0_TestBlock__B_op89 <= TestBlock__B_op89;
    p0_TestBlock__B_op90 <= TestBlock__B_op90;
    p0_TestBlock__B_op91 <= TestBlock__B_op91;
    p0_TestBlock__B_op92 <= TestBlock__B_op92;
    p0_TestBlock__B_op93 <= TestBlock__B_op93;
    p0_TestBlock__B_op94 <= TestBlock__B_op94;
    p0_TestBlock__B_op95 <= TestBlock__B_op95;
    p0_TestBlock__B_op96 <= TestBlock__B_op96;
    p0_TestBlock__B_op97 <= TestBlock__B_op97;
    p0_TestBlock__B_op98 <= TestBlock__B_op98;
    p0_TestBlock__B_op99 <= TestBlock__B_op99;
  end

  // ===== Pipe stage 1:
  wire [31:0] p1_smul_89499_comb;
  wire [31:0] p1_smul_89500_comb;
  wire [31:0] p1_smul_89501_comb;
  wire [31:0] p1_smul_89502_comb;
  wire [31:0] p1_smul_89899_comb;
  wire [31:0] p1_smul_89900_comb;
  wire [31:0] p1_smul_89901_comb;
  wire [31:0] p1_smul_89902_comb;
  wire [31:0] p1_smul_89903_comb;
  wire [31:0] p1_smul_89904_comb;
  wire [31:0] p1_smul_89503_comb;
  wire [31:0] p1_smul_89504_comb;
  wire [31:0] p1_smul_89505_comb;
  wire [31:0] p1_smul_89506_comb;
  wire [31:0] p1_smul_89905_comb;
  wire [31:0] p1_smul_89906_comb;
  wire [31:0] p1_smul_89907_comb;
  wire [31:0] p1_smul_89908_comb;
  wire [31:0] p1_smul_89909_comb;
  wire [31:0] p1_smul_89910_comb;
  wire [31:0] p1_smul_89507_comb;
  wire [31:0] p1_smul_89508_comb;
  wire [31:0] p1_smul_89509_comb;
  wire [31:0] p1_smul_89510_comb;
  wire [31:0] p1_smul_89911_comb;
  wire [31:0] p1_smul_89912_comb;
  wire [31:0] p1_smul_89913_comb;
  wire [31:0] p1_smul_89914_comb;
  wire [31:0] p1_smul_89915_comb;
  wire [31:0] p1_smul_89916_comb;
  wire [31:0] p1_smul_89511_comb;
  wire [31:0] p1_smul_89512_comb;
  wire [31:0] p1_smul_89513_comb;
  wire [31:0] p1_smul_89514_comb;
  wire [31:0] p1_smul_89917_comb;
  wire [31:0] p1_smul_89918_comb;
  wire [31:0] p1_smul_89919_comb;
  wire [31:0] p1_smul_89920_comb;
  wire [31:0] p1_smul_89921_comb;
  wire [31:0] p1_smul_89922_comb;
  wire [31:0] p1_smul_89515_comb;
  wire [31:0] p1_smul_89516_comb;
  wire [31:0] p1_smul_89517_comb;
  wire [31:0] p1_smul_89518_comb;
  wire [31:0] p1_smul_89923_comb;
  wire [31:0] p1_smul_89924_comb;
  wire [31:0] p1_smul_89925_comb;
  wire [31:0] p1_smul_89926_comb;
  wire [31:0] p1_smul_89927_comb;
  wire [31:0] p1_smul_89928_comb;
  wire [31:0] p1_smul_89519_comb;
  wire [31:0] p1_smul_89520_comb;
  wire [31:0] p1_smul_89521_comb;
  wire [31:0] p1_smul_89522_comb;
  wire [31:0] p1_smul_89929_comb;
  wire [31:0] p1_smul_89930_comb;
  wire [31:0] p1_smul_89931_comb;
  wire [31:0] p1_smul_89932_comb;
  wire [31:0] p1_smul_89933_comb;
  wire [31:0] p1_smul_89934_comb;
  wire [31:0] p1_smul_89523_comb;
  wire [31:0] p1_smul_89524_comb;
  wire [31:0] p1_smul_89525_comb;
  wire [31:0] p1_smul_89526_comb;
  wire [31:0] p1_smul_89935_comb;
  wire [31:0] p1_smul_89936_comb;
  wire [31:0] p1_smul_89937_comb;
  wire [31:0] p1_smul_89938_comb;
  wire [31:0] p1_smul_89939_comb;
  wire [31:0] p1_smul_89940_comb;
  wire [31:0] p1_smul_89527_comb;
  wire [31:0] p1_smul_89528_comb;
  wire [31:0] p1_smul_89529_comb;
  wire [31:0] p1_smul_89530_comb;
  wire [31:0] p1_smul_89941_comb;
  wire [31:0] p1_smul_89942_comb;
  wire [31:0] p1_smul_89943_comb;
  wire [31:0] p1_smul_89944_comb;
  wire [31:0] p1_smul_89945_comb;
  wire [31:0] p1_smul_89946_comb;
  wire [31:0] p1_smul_89531_comb;
  wire [31:0] p1_smul_89532_comb;
  wire [31:0] p1_smul_89533_comb;
  wire [31:0] p1_smul_89534_comb;
  wire [31:0] p1_smul_89947_comb;
  wire [31:0] p1_smul_89948_comb;
  wire [31:0] p1_smul_89949_comb;
  wire [31:0] p1_smul_89950_comb;
  wire [31:0] p1_smul_89951_comb;
  wire [31:0] p1_smul_89952_comb;
  wire [31:0] p1_smul_89535_comb;
  wire [31:0] p1_smul_89536_comb;
  wire [31:0] p1_smul_89537_comb;
  wire [31:0] p1_smul_89538_comb;
  wire [31:0] p1_smul_89953_comb;
  wire [31:0] p1_smul_89954_comb;
  wire [31:0] p1_smul_89955_comb;
  wire [31:0] p1_smul_89956_comb;
  wire [31:0] p1_smul_89957_comb;
  wire [31:0] p1_smul_89958_comb;
  wire [31:0] p1_smul_89539_comb;
  wire [31:0] p1_smul_89540_comb;
  wire [31:0] p1_smul_89541_comb;
  wire [31:0] p1_smul_89542_comb;
  wire [31:0] p1_smul_89959_comb;
  wire [31:0] p1_smul_89960_comb;
  wire [31:0] p1_smul_89961_comb;
  wire [31:0] p1_smul_89962_comb;
  wire [31:0] p1_smul_89963_comb;
  wire [31:0] p1_smul_89964_comb;
  wire [31:0] p1_smul_89543_comb;
  wire [31:0] p1_smul_89544_comb;
  wire [31:0] p1_smul_89545_comb;
  wire [31:0] p1_smul_89546_comb;
  wire [31:0] p1_smul_89965_comb;
  wire [31:0] p1_smul_89966_comb;
  wire [31:0] p1_smul_89967_comb;
  wire [31:0] p1_smul_89968_comb;
  wire [31:0] p1_smul_89969_comb;
  wire [31:0] p1_smul_89970_comb;
  wire [31:0] p1_smul_89547_comb;
  wire [31:0] p1_smul_89548_comb;
  wire [31:0] p1_smul_89549_comb;
  wire [31:0] p1_smul_89550_comb;
  wire [31:0] p1_smul_89971_comb;
  wire [31:0] p1_smul_89972_comb;
  wire [31:0] p1_smul_89973_comb;
  wire [31:0] p1_smul_89974_comb;
  wire [31:0] p1_smul_89975_comb;
  wire [31:0] p1_smul_89976_comb;
  wire [31:0] p1_smul_89551_comb;
  wire [31:0] p1_smul_89552_comb;
  wire [31:0] p1_smul_89553_comb;
  wire [31:0] p1_smul_89554_comb;
  wire [31:0] p1_smul_89977_comb;
  wire [31:0] p1_smul_89978_comb;
  wire [31:0] p1_smul_89979_comb;
  wire [31:0] p1_smul_89980_comb;
  wire [31:0] p1_smul_89981_comb;
  wire [31:0] p1_smul_89982_comb;
  wire [31:0] p1_smul_89555_comb;
  wire [31:0] p1_smul_89556_comb;
  wire [31:0] p1_smul_89557_comb;
  wire [31:0] p1_smul_89558_comb;
  wire [31:0] p1_smul_89983_comb;
  wire [31:0] p1_smul_89984_comb;
  wire [31:0] p1_smul_89985_comb;
  wire [31:0] p1_smul_89986_comb;
  wire [31:0] p1_smul_89987_comb;
  wire [31:0] p1_smul_89988_comb;
  wire [31:0] p1_smul_89559_comb;
  wire [31:0] p1_smul_89560_comb;
  wire [31:0] p1_smul_89561_comb;
  wire [31:0] p1_smul_89562_comb;
  wire [31:0] p1_smul_89989_comb;
  wire [31:0] p1_smul_89990_comb;
  wire [31:0] p1_smul_89991_comb;
  wire [31:0] p1_smul_89992_comb;
  wire [31:0] p1_smul_89993_comb;
  wire [31:0] p1_smul_89994_comb;
  wire [31:0] p1_smul_89563_comb;
  wire [31:0] p1_smul_89564_comb;
  wire [31:0] p1_smul_89565_comb;
  wire [31:0] p1_smul_89566_comb;
  wire [31:0] p1_smul_89995_comb;
  wire [31:0] p1_smul_89996_comb;
  wire [31:0] p1_smul_89997_comb;
  wire [31:0] p1_smul_89998_comb;
  wire [31:0] p1_smul_89999_comb;
  wire [31:0] p1_smul_90000_comb;
  wire [31:0] p1_smul_89567_comb;
  wire [31:0] p1_smul_89568_comb;
  wire [31:0] p1_smul_89569_comb;
  wire [31:0] p1_smul_89570_comb;
  wire [31:0] p1_smul_90001_comb;
  wire [31:0] p1_smul_90002_comb;
  wire [31:0] p1_smul_90003_comb;
  wire [31:0] p1_smul_90004_comb;
  wire [31:0] p1_smul_90005_comb;
  wire [31:0] p1_smul_90006_comb;
  wire [31:0] p1_smul_89571_comb;
  wire [31:0] p1_smul_89572_comb;
  wire [31:0] p1_smul_89573_comb;
  wire [31:0] p1_smul_89574_comb;
  wire [31:0] p1_smul_90007_comb;
  wire [31:0] p1_smul_90008_comb;
  wire [31:0] p1_smul_90009_comb;
  wire [31:0] p1_smul_90010_comb;
  wire [31:0] p1_smul_90011_comb;
  wire [31:0] p1_smul_90012_comb;
  wire [31:0] p1_smul_89575_comb;
  wire [31:0] p1_smul_89576_comb;
  wire [31:0] p1_smul_89577_comb;
  wire [31:0] p1_smul_89578_comb;
  wire [31:0] p1_smul_90013_comb;
  wire [31:0] p1_smul_90014_comb;
  wire [31:0] p1_smul_90015_comb;
  wire [31:0] p1_smul_90016_comb;
  wire [31:0] p1_smul_90017_comb;
  wire [31:0] p1_smul_90018_comb;
  wire [31:0] p1_smul_89579_comb;
  wire [31:0] p1_smul_89580_comb;
  wire [31:0] p1_smul_89581_comb;
  wire [31:0] p1_smul_89582_comb;
  wire [31:0] p1_smul_90019_comb;
  wire [31:0] p1_smul_90020_comb;
  wire [31:0] p1_smul_90021_comb;
  wire [31:0] p1_smul_90022_comb;
  wire [31:0] p1_smul_90023_comb;
  wire [31:0] p1_smul_90024_comb;
  wire [31:0] p1_smul_89583_comb;
  wire [31:0] p1_smul_89584_comb;
  wire [31:0] p1_smul_89585_comb;
  wire [31:0] p1_smul_89586_comb;
  wire [31:0] p1_smul_90025_comb;
  wire [31:0] p1_smul_90026_comb;
  wire [31:0] p1_smul_90027_comb;
  wire [31:0] p1_smul_90028_comb;
  wire [31:0] p1_smul_90029_comb;
  wire [31:0] p1_smul_90030_comb;
  wire [31:0] p1_smul_89587_comb;
  wire [31:0] p1_smul_89588_comb;
  wire [31:0] p1_smul_89589_comb;
  wire [31:0] p1_smul_89590_comb;
  wire [31:0] p1_smul_90031_comb;
  wire [31:0] p1_smul_90032_comb;
  wire [31:0] p1_smul_90033_comb;
  wire [31:0] p1_smul_90034_comb;
  wire [31:0] p1_smul_90035_comb;
  wire [31:0] p1_smul_90036_comb;
  wire [31:0] p1_smul_89591_comb;
  wire [31:0] p1_smul_89592_comb;
  wire [31:0] p1_smul_89593_comb;
  wire [31:0] p1_smul_89594_comb;
  wire [31:0] p1_smul_90037_comb;
  wire [31:0] p1_smul_90038_comb;
  wire [31:0] p1_smul_90039_comb;
  wire [31:0] p1_smul_90040_comb;
  wire [31:0] p1_smul_90041_comb;
  wire [31:0] p1_smul_90042_comb;
  wire [31:0] p1_smul_89595_comb;
  wire [31:0] p1_smul_89596_comb;
  wire [31:0] p1_smul_89597_comb;
  wire [31:0] p1_smul_89598_comb;
  wire [31:0] p1_smul_90043_comb;
  wire [31:0] p1_smul_90044_comb;
  wire [31:0] p1_smul_90045_comb;
  wire [31:0] p1_smul_90046_comb;
  wire [31:0] p1_smul_90047_comb;
  wire [31:0] p1_smul_90048_comb;
  wire [31:0] p1_smul_89599_comb;
  wire [31:0] p1_smul_89600_comb;
  wire [31:0] p1_smul_89601_comb;
  wire [31:0] p1_smul_89602_comb;
  wire [31:0] p1_smul_90049_comb;
  wire [31:0] p1_smul_90050_comb;
  wire [31:0] p1_smul_90051_comb;
  wire [31:0] p1_smul_90052_comb;
  wire [31:0] p1_smul_90053_comb;
  wire [31:0] p1_smul_90054_comb;
  wire [31:0] p1_smul_89603_comb;
  wire [31:0] p1_smul_89604_comb;
  wire [31:0] p1_smul_89605_comb;
  wire [31:0] p1_smul_89606_comb;
  wire [31:0] p1_smul_90055_comb;
  wire [31:0] p1_smul_90056_comb;
  wire [31:0] p1_smul_90057_comb;
  wire [31:0] p1_smul_90058_comb;
  wire [31:0] p1_smul_90059_comb;
  wire [31:0] p1_smul_90060_comb;
  wire [31:0] p1_smul_89607_comb;
  wire [31:0] p1_smul_89608_comb;
  wire [31:0] p1_smul_89609_comb;
  wire [31:0] p1_smul_89610_comb;
  wire [31:0] p1_smul_90061_comb;
  wire [31:0] p1_smul_90062_comb;
  wire [31:0] p1_smul_90063_comb;
  wire [31:0] p1_smul_90064_comb;
  wire [31:0] p1_smul_90065_comb;
  wire [31:0] p1_smul_90066_comb;
  wire [31:0] p1_smul_89611_comb;
  wire [31:0] p1_smul_89612_comb;
  wire [31:0] p1_smul_89613_comb;
  wire [31:0] p1_smul_89614_comb;
  wire [31:0] p1_smul_90067_comb;
  wire [31:0] p1_smul_90068_comb;
  wire [31:0] p1_smul_90069_comb;
  wire [31:0] p1_smul_90070_comb;
  wire [31:0] p1_smul_90071_comb;
  wire [31:0] p1_smul_90072_comb;
  wire [31:0] p1_smul_89615_comb;
  wire [31:0] p1_smul_89616_comb;
  wire [31:0] p1_smul_89617_comb;
  wire [31:0] p1_smul_89618_comb;
  wire [31:0] p1_smul_90073_comb;
  wire [31:0] p1_smul_90074_comb;
  wire [31:0] p1_smul_90075_comb;
  wire [31:0] p1_smul_90076_comb;
  wire [31:0] p1_smul_90077_comb;
  wire [31:0] p1_smul_90078_comb;
  wire [31:0] p1_smul_89619_comb;
  wire [31:0] p1_smul_89620_comb;
  wire [31:0] p1_smul_89621_comb;
  wire [31:0] p1_smul_89622_comb;
  wire [31:0] p1_smul_90079_comb;
  wire [31:0] p1_smul_90080_comb;
  wire [31:0] p1_smul_90081_comb;
  wire [31:0] p1_smul_90082_comb;
  wire [31:0] p1_smul_90083_comb;
  wire [31:0] p1_smul_90084_comb;
  wire [31:0] p1_smul_89623_comb;
  wire [31:0] p1_smul_89624_comb;
  wire [31:0] p1_smul_89625_comb;
  wire [31:0] p1_smul_89626_comb;
  wire [31:0] p1_smul_90085_comb;
  wire [31:0] p1_smul_90086_comb;
  wire [31:0] p1_smul_90087_comb;
  wire [31:0] p1_smul_90088_comb;
  wire [31:0] p1_smul_90089_comb;
  wire [31:0] p1_smul_90090_comb;
  wire [31:0] p1_smul_89627_comb;
  wire [31:0] p1_smul_89628_comb;
  wire [31:0] p1_smul_89629_comb;
  wire [31:0] p1_smul_89630_comb;
  wire [31:0] p1_smul_90091_comb;
  wire [31:0] p1_smul_90092_comb;
  wire [31:0] p1_smul_90093_comb;
  wire [31:0] p1_smul_90094_comb;
  wire [31:0] p1_smul_90095_comb;
  wire [31:0] p1_smul_90096_comb;
  wire [31:0] p1_smul_89631_comb;
  wire [31:0] p1_smul_89632_comb;
  wire [31:0] p1_smul_89633_comb;
  wire [31:0] p1_smul_89634_comb;
  wire [31:0] p1_smul_90097_comb;
  wire [31:0] p1_smul_90098_comb;
  wire [31:0] p1_smul_90099_comb;
  wire [31:0] p1_smul_90100_comb;
  wire [31:0] p1_smul_90101_comb;
  wire [31:0] p1_smul_90102_comb;
  wire [31:0] p1_smul_89635_comb;
  wire [31:0] p1_smul_89636_comb;
  wire [31:0] p1_smul_89637_comb;
  wire [31:0] p1_smul_89638_comb;
  wire [31:0] p1_smul_90103_comb;
  wire [31:0] p1_smul_90104_comb;
  wire [31:0] p1_smul_90105_comb;
  wire [31:0] p1_smul_90106_comb;
  wire [31:0] p1_smul_90107_comb;
  wire [31:0] p1_smul_90108_comb;
  wire [31:0] p1_smul_89639_comb;
  wire [31:0] p1_smul_89640_comb;
  wire [31:0] p1_smul_89641_comb;
  wire [31:0] p1_smul_89642_comb;
  wire [31:0] p1_smul_90109_comb;
  wire [31:0] p1_smul_90110_comb;
  wire [31:0] p1_smul_90111_comb;
  wire [31:0] p1_smul_90112_comb;
  wire [31:0] p1_smul_90113_comb;
  wire [31:0] p1_smul_90114_comb;
  wire [31:0] p1_smul_89643_comb;
  wire [31:0] p1_smul_89644_comb;
  wire [31:0] p1_smul_89645_comb;
  wire [31:0] p1_smul_89646_comb;
  wire [31:0] p1_smul_90115_comb;
  wire [31:0] p1_smul_90116_comb;
  wire [31:0] p1_smul_90117_comb;
  wire [31:0] p1_smul_90118_comb;
  wire [31:0] p1_smul_90119_comb;
  wire [31:0] p1_smul_90120_comb;
  wire [31:0] p1_smul_89647_comb;
  wire [31:0] p1_smul_89648_comb;
  wire [31:0] p1_smul_89649_comb;
  wire [31:0] p1_smul_89650_comb;
  wire [31:0] p1_smul_90121_comb;
  wire [31:0] p1_smul_90122_comb;
  wire [31:0] p1_smul_90123_comb;
  wire [31:0] p1_smul_90124_comb;
  wire [31:0] p1_smul_90125_comb;
  wire [31:0] p1_smul_90126_comb;
  wire [31:0] p1_smul_89651_comb;
  wire [31:0] p1_smul_89652_comb;
  wire [31:0] p1_smul_89653_comb;
  wire [31:0] p1_smul_89654_comb;
  wire [31:0] p1_smul_90127_comb;
  wire [31:0] p1_smul_90128_comb;
  wire [31:0] p1_smul_90129_comb;
  wire [31:0] p1_smul_90130_comb;
  wire [31:0] p1_smul_90131_comb;
  wire [31:0] p1_smul_90132_comb;
  wire [31:0] p1_smul_89655_comb;
  wire [31:0] p1_smul_89656_comb;
  wire [31:0] p1_smul_89657_comb;
  wire [31:0] p1_smul_89658_comb;
  wire [31:0] p1_smul_90133_comb;
  wire [31:0] p1_smul_90134_comb;
  wire [31:0] p1_smul_90135_comb;
  wire [31:0] p1_smul_90136_comb;
  wire [31:0] p1_smul_90137_comb;
  wire [31:0] p1_smul_90138_comb;
  wire [31:0] p1_smul_89659_comb;
  wire [31:0] p1_smul_89660_comb;
  wire [31:0] p1_smul_89661_comb;
  wire [31:0] p1_smul_89662_comb;
  wire [31:0] p1_smul_90139_comb;
  wire [31:0] p1_smul_90140_comb;
  wire [31:0] p1_smul_90141_comb;
  wire [31:0] p1_smul_90142_comb;
  wire [31:0] p1_smul_90143_comb;
  wire [31:0] p1_smul_90144_comb;
  wire [31:0] p1_smul_89663_comb;
  wire [31:0] p1_smul_89664_comb;
  wire [31:0] p1_smul_89665_comb;
  wire [31:0] p1_smul_89666_comb;
  wire [31:0] p1_smul_90145_comb;
  wire [31:0] p1_smul_90146_comb;
  wire [31:0] p1_smul_90147_comb;
  wire [31:0] p1_smul_90148_comb;
  wire [31:0] p1_smul_90149_comb;
  wire [31:0] p1_smul_90150_comb;
  wire [31:0] p1_smul_89667_comb;
  wire [31:0] p1_smul_89668_comb;
  wire [31:0] p1_smul_89669_comb;
  wire [31:0] p1_smul_89670_comb;
  wire [31:0] p1_smul_90151_comb;
  wire [31:0] p1_smul_90152_comb;
  wire [31:0] p1_smul_90153_comb;
  wire [31:0] p1_smul_90154_comb;
  wire [31:0] p1_smul_90155_comb;
  wire [31:0] p1_smul_90156_comb;
  wire [31:0] p1_smul_89671_comb;
  wire [31:0] p1_smul_89672_comb;
  wire [31:0] p1_smul_89673_comb;
  wire [31:0] p1_smul_89674_comb;
  wire [31:0] p1_smul_90157_comb;
  wire [31:0] p1_smul_90158_comb;
  wire [31:0] p1_smul_90159_comb;
  wire [31:0] p1_smul_90160_comb;
  wire [31:0] p1_smul_90161_comb;
  wire [31:0] p1_smul_90162_comb;
  wire [31:0] p1_smul_89675_comb;
  wire [31:0] p1_smul_89676_comb;
  wire [31:0] p1_smul_89677_comb;
  wire [31:0] p1_smul_89678_comb;
  wire [31:0] p1_smul_90163_comb;
  wire [31:0] p1_smul_90164_comb;
  wire [31:0] p1_smul_90165_comb;
  wire [31:0] p1_smul_90166_comb;
  wire [31:0] p1_smul_90167_comb;
  wire [31:0] p1_smul_90168_comb;
  wire [31:0] p1_smul_89679_comb;
  wire [31:0] p1_smul_89680_comb;
  wire [31:0] p1_smul_89681_comb;
  wire [31:0] p1_smul_89682_comb;
  wire [31:0] p1_smul_90169_comb;
  wire [31:0] p1_smul_90170_comb;
  wire [31:0] p1_smul_90171_comb;
  wire [31:0] p1_smul_90172_comb;
  wire [31:0] p1_smul_90173_comb;
  wire [31:0] p1_smul_90174_comb;
  wire [31:0] p1_smul_89683_comb;
  wire [31:0] p1_smul_89684_comb;
  wire [31:0] p1_smul_89685_comb;
  wire [31:0] p1_smul_89686_comb;
  wire [31:0] p1_smul_90175_comb;
  wire [31:0] p1_smul_90176_comb;
  wire [31:0] p1_smul_90177_comb;
  wire [31:0] p1_smul_90178_comb;
  wire [31:0] p1_smul_90179_comb;
  wire [31:0] p1_smul_90180_comb;
  wire [31:0] p1_smul_89687_comb;
  wire [31:0] p1_smul_89688_comb;
  wire [31:0] p1_smul_89689_comb;
  wire [31:0] p1_smul_89690_comb;
  wire [31:0] p1_smul_90181_comb;
  wire [31:0] p1_smul_90182_comb;
  wire [31:0] p1_smul_90183_comb;
  wire [31:0] p1_smul_90184_comb;
  wire [31:0] p1_smul_90185_comb;
  wire [31:0] p1_smul_90186_comb;
  wire [31:0] p1_smul_89691_comb;
  wire [31:0] p1_smul_89692_comb;
  wire [31:0] p1_smul_89693_comb;
  wire [31:0] p1_smul_89694_comb;
  wire [31:0] p1_smul_90187_comb;
  wire [31:0] p1_smul_90188_comb;
  wire [31:0] p1_smul_90189_comb;
  wire [31:0] p1_smul_90190_comb;
  wire [31:0] p1_smul_90191_comb;
  wire [31:0] p1_smul_90192_comb;
  wire [31:0] p1_smul_89695_comb;
  wire [31:0] p1_smul_89696_comb;
  wire [31:0] p1_smul_89697_comb;
  wire [31:0] p1_smul_89698_comb;
  wire [31:0] p1_smul_90193_comb;
  wire [31:0] p1_smul_90194_comb;
  wire [31:0] p1_smul_90195_comb;
  wire [31:0] p1_smul_90196_comb;
  wire [31:0] p1_smul_90197_comb;
  wire [31:0] p1_smul_90198_comb;
  wire [31:0] p1_smul_89699_comb;
  wire [31:0] p1_smul_89700_comb;
  wire [31:0] p1_smul_89701_comb;
  wire [31:0] p1_smul_89702_comb;
  wire [31:0] p1_smul_90199_comb;
  wire [31:0] p1_smul_90200_comb;
  wire [31:0] p1_smul_90201_comb;
  wire [31:0] p1_smul_90202_comb;
  wire [31:0] p1_smul_90203_comb;
  wire [31:0] p1_smul_90204_comb;
  wire [31:0] p1_smul_89703_comb;
  wire [31:0] p1_smul_89704_comb;
  wire [31:0] p1_smul_89705_comb;
  wire [31:0] p1_smul_89706_comb;
  wire [31:0] p1_smul_90205_comb;
  wire [31:0] p1_smul_90206_comb;
  wire [31:0] p1_smul_90207_comb;
  wire [31:0] p1_smul_90208_comb;
  wire [31:0] p1_smul_90209_comb;
  wire [31:0] p1_smul_90210_comb;
  wire [31:0] p1_smul_89707_comb;
  wire [31:0] p1_smul_89708_comb;
  wire [31:0] p1_smul_89709_comb;
  wire [31:0] p1_smul_89710_comb;
  wire [31:0] p1_smul_90211_comb;
  wire [31:0] p1_smul_90212_comb;
  wire [31:0] p1_smul_90213_comb;
  wire [31:0] p1_smul_90214_comb;
  wire [31:0] p1_smul_90215_comb;
  wire [31:0] p1_smul_90216_comb;
  wire [31:0] p1_smul_89711_comb;
  wire [31:0] p1_smul_89712_comb;
  wire [31:0] p1_smul_89713_comb;
  wire [31:0] p1_smul_89714_comb;
  wire [31:0] p1_smul_90217_comb;
  wire [31:0] p1_smul_90218_comb;
  wire [31:0] p1_smul_90219_comb;
  wire [31:0] p1_smul_90220_comb;
  wire [31:0] p1_smul_90221_comb;
  wire [31:0] p1_smul_90222_comb;
  wire [31:0] p1_smul_89715_comb;
  wire [31:0] p1_smul_89716_comb;
  wire [31:0] p1_smul_89717_comb;
  wire [31:0] p1_smul_89718_comb;
  wire [31:0] p1_smul_90223_comb;
  wire [31:0] p1_smul_90224_comb;
  wire [31:0] p1_smul_90225_comb;
  wire [31:0] p1_smul_90226_comb;
  wire [31:0] p1_smul_90227_comb;
  wire [31:0] p1_smul_90228_comb;
  wire [31:0] p1_smul_89719_comb;
  wire [31:0] p1_smul_89720_comb;
  wire [31:0] p1_smul_89721_comb;
  wire [31:0] p1_smul_89722_comb;
  wire [31:0] p1_smul_90229_comb;
  wire [31:0] p1_smul_90230_comb;
  wire [31:0] p1_smul_90231_comb;
  wire [31:0] p1_smul_90232_comb;
  wire [31:0] p1_smul_90233_comb;
  wire [31:0] p1_smul_90234_comb;
  wire [31:0] p1_smul_89723_comb;
  wire [31:0] p1_smul_89724_comb;
  wire [31:0] p1_smul_89725_comb;
  wire [31:0] p1_smul_89726_comb;
  wire [31:0] p1_smul_90235_comb;
  wire [31:0] p1_smul_90236_comb;
  wire [31:0] p1_smul_90237_comb;
  wire [31:0] p1_smul_90238_comb;
  wire [31:0] p1_smul_90239_comb;
  wire [31:0] p1_smul_90240_comb;
  wire [31:0] p1_smul_89727_comb;
  wire [31:0] p1_smul_89728_comb;
  wire [31:0] p1_smul_89729_comb;
  wire [31:0] p1_smul_89730_comb;
  wire [31:0] p1_smul_90241_comb;
  wire [31:0] p1_smul_90242_comb;
  wire [31:0] p1_smul_90243_comb;
  wire [31:0] p1_smul_90244_comb;
  wire [31:0] p1_smul_90245_comb;
  wire [31:0] p1_smul_90246_comb;
  wire [31:0] p1_smul_89731_comb;
  wire [31:0] p1_smul_89732_comb;
  wire [31:0] p1_smul_89733_comb;
  wire [31:0] p1_smul_89734_comb;
  wire [31:0] p1_smul_90247_comb;
  wire [31:0] p1_smul_90248_comb;
  wire [31:0] p1_smul_90249_comb;
  wire [31:0] p1_smul_90250_comb;
  wire [31:0] p1_smul_90251_comb;
  wire [31:0] p1_smul_90252_comb;
  wire [31:0] p1_smul_89735_comb;
  wire [31:0] p1_smul_89736_comb;
  wire [31:0] p1_smul_89737_comb;
  wire [31:0] p1_smul_89738_comb;
  wire [31:0] p1_smul_90253_comb;
  wire [31:0] p1_smul_90254_comb;
  wire [31:0] p1_smul_90255_comb;
  wire [31:0] p1_smul_90256_comb;
  wire [31:0] p1_smul_90257_comb;
  wire [31:0] p1_smul_90258_comb;
  wire [31:0] p1_smul_89739_comb;
  wire [31:0] p1_smul_89740_comb;
  wire [31:0] p1_smul_89741_comb;
  wire [31:0] p1_smul_89742_comb;
  wire [31:0] p1_smul_90259_comb;
  wire [31:0] p1_smul_90260_comb;
  wire [31:0] p1_smul_90261_comb;
  wire [31:0] p1_smul_90262_comb;
  wire [31:0] p1_smul_90263_comb;
  wire [31:0] p1_smul_90264_comb;
  wire [31:0] p1_smul_89743_comb;
  wire [31:0] p1_smul_89744_comb;
  wire [31:0] p1_smul_89745_comb;
  wire [31:0] p1_smul_89746_comb;
  wire [31:0] p1_smul_90265_comb;
  wire [31:0] p1_smul_90266_comb;
  wire [31:0] p1_smul_90267_comb;
  wire [31:0] p1_smul_90268_comb;
  wire [31:0] p1_smul_90269_comb;
  wire [31:0] p1_smul_90270_comb;
  wire [31:0] p1_smul_89747_comb;
  wire [31:0] p1_smul_89748_comb;
  wire [31:0] p1_smul_89749_comb;
  wire [31:0] p1_smul_89750_comb;
  wire [31:0] p1_smul_90271_comb;
  wire [31:0] p1_smul_90272_comb;
  wire [31:0] p1_smul_90273_comb;
  wire [31:0] p1_smul_90274_comb;
  wire [31:0] p1_smul_90275_comb;
  wire [31:0] p1_smul_90276_comb;
  wire [31:0] p1_smul_89751_comb;
  wire [31:0] p1_smul_89752_comb;
  wire [31:0] p1_smul_89753_comb;
  wire [31:0] p1_smul_89754_comb;
  wire [31:0] p1_smul_90277_comb;
  wire [31:0] p1_smul_90278_comb;
  wire [31:0] p1_smul_90279_comb;
  wire [31:0] p1_smul_90280_comb;
  wire [31:0] p1_smul_90281_comb;
  wire [31:0] p1_smul_90282_comb;
  wire [31:0] p1_smul_89755_comb;
  wire [31:0] p1_smul_89756_comb;
  wire [31:0] p1_smul_89757_comb;
  wire [31:0] p1_smul_89758_comb;
  wire [31:0] p1_smul_90283_comb;
  wire [31:0] p1_smul_90284_comb;
  wire [31:0] p1_smul_90285_comb;
  wire [31:0] p1_smul_90286_comb;
  wire [31:0] p1_smul_90287_comb;
  wire [31:0] p1_smul_90288_comb;
  wire [31:0] p1_smul_89759_comb;
  wire [31:0] p1_smul_89760_comb;
  wire [31:0] p1_smul_89761_comb;
  wire [31:0] p1_smul_89762_comb;
  wire [31:0] p1_smul_90289_comb;
  wire [31:0] p1_smul_90290_comb;
  wire [31:0] p1_smul_90291_comb;
  wire [31:0] p1_smul_90292_comb;
  wire [31:0] p1_smul_90293_comb;
  wire [31:0] p1_smul_90294_comb;
  wire [31:0] p1_smul_89763_comb;
  wire [31:0] p1_smul_89764_comb;
  wire [31:0] p1_smul_89765_comb;
  wire [31:0] p1_smul_89766_comb;
  wire [31:0] p1_smul_90295_comb;
  wire [31:0] p1_smul_90296_comb;
  wire [31:0] p1_smul_90297_comb;
  wire [31:0] p1_smul_90298_comb;
  wire [31:0] p1_smul_90299_comb;
  wire [31:0] p1_smul_90300_comb;
  wire [31:0] p1_smul_89767_comb;
  wire [31:0] p1_smul_89768_comb;
  wire [31:0] p1_smul_89769_comb;
  wire [31:0] p1_smul_89770_comb;
  wire [31:0] p1_smul_90301_comb;
  wire [31:0] p1_smul_90302_comb;
  wire [31:0] p1_smul_90303_comb;
  wire [31:0] p1_smul_90304_comb;
  wire [31:0] p1_smul_90305_comb;
  wire [31:0] p1_smul_90306_comb;
  wire [31:0] p1_smul_89771_comb;
  wire [31:0] p1_smul_89772_comb;
  wire [31:0] p1_smul_89773_comb;
  wire [31:0] p1_smul_89774_comb;
  wire [31:0] p1_smul_90307_comb;
  wire [31:0] p1_smul_90308_comb;
  wire [31:0] p1_smul_90309_comb;
  wire [31:0] p1_smul_90310_comb;
  wire [31:0] p1_smul_90311_comb;
  wire [31:0] p1_smul_90312_comb;
  wire [31:0] p1_smul_89775_comb;
  wire [31:0] p1_smul_89776_comb;
  wire [31:0] p1_smul_89777_comb;
  wire [31:0] p1_smul_89778_comb;
  wire [31:0] p1_smul_90313_comb;
  wire [31:0] p1_smul_90314_comb;
  wire [31:0] p1_smul_90315_comb;
  wire [31:0] p1_smul_90316_comb;
  wire [31:0] p1_smul_90317_comb;
  wire [31:0] p1_smul_90318_comb;
  wire [31:0] p1_smul_89779_comb;
  wire [31:0] p1_smul_89780_comb;
  wire [31:0] p1_smul_89781_comb;
  wire [31:0] p1_smul_89782_comb;
  wire [31:0] p1_smul_90319_comb;
  wire [31:0] p1_smul_90320_comb;
  wire [31:0] p1_smul_90321_comb;
  wire [31:0] p1_smul_90322_comb;
  wire [31:0] p1_smul_90323_comb;
  wire [31:0] p1_smul_90324_comb;
  wire [31:0] p1_smul_89783_comb;
  wire [31:0] p1_smul_89784_comb;
  wire [31:0] p1_smul_89785_comb;
  wire [31:0] p1_smul_89786_comb;
  wire [31:0] p1_smul_90325_comb;
  wire [31:0] p1_smul_90326_comb;
  wire [31:0] p1_smul_90327_comb;
  wire [31:0] p1_smul_90328_comb;
  wire [31:0] p1_smul_90329_comb;
  wire [31:0] p1_smul_90330_comb;
  wire [31:0] p1_smul_89787_comb;
  wire [31:0] p1_smul_89788_comb;
  wire [31:0] p1_smul_89789_comb;
  wire [31:0] p1_smul_89790_comb;
  wire [31:0] p1_smul_90331_comb;
  wire [31:0] p1_smul_90332_comb;
  wire [31:0] p1_smul_90333_comb;
  wire [31:0] p1_smul_90334_comb;
  wire [31:0] p1_smul_90335_comb;
  wire [31:0] p1_smul_90336_comb;
  wire [31:0] p1_smul_89791_comb;
  wire [31:0] p1_smul_89792_comb;
  wire [31:0] p1_smul_89793_comb;
  wire [31:0] p1_smul_89794_comb;
  wire [31:0] p1_smul_90337_comb;
  wire [31:0] p1_smul_90338_comb;
  wire [31:0] p1_smul_90339_comb;
  wire [31:0] p1_smul_90340_comb;
  wire [31:0] p1_smul_90341_comb;
  wire [31:0] p1_smul_90342_comb;
  wire [31:0] p1_smul_89795_comb;
  wire [31:0] p1_smul_89796_comb;
  wire [31:0] p1_smul_89797_comb;
  wire [31:0] p1_smul_89798_comb;
  wire [31:0] p1_smul_90343_comb;
  wire [31:0] p1_smul_90344_comb;
  wire [31:0] p1_smul_90345_comb;
  wire [31:0] p1_smul_90346_comb;
  wire [31:0] p1_smul_90347_comb;
  wire [31:0] p1_smul_90348_comb;
  wire [31:0] p1_smul_89799_comb;
  wire [31:0] p1_smul_89800_comb;
  wire [31:0] p1_smul_89801_comb;
  wire [31:0] p1_smul_89802_comb;
  wire [31:0] p1_smul_90349_comb;
  wire [31:0] p1_smul_90350_comb;
  wire [31:0] p1_smul_90351_comb;
  wire [31:0] p1_smul_90352_comb;
  wire [31:0] p1_smul_90353_comb;
  wire [31:0] p1_smul_90354_comb;
  wire [31:0] p1_smul_89803_comb;
  wire [31:0] p1_smul_89804_comb;
  wire [31:0] p1_smul_89805_comb;
  wire [31:0] p1_smul_89806_comb;
  wire [31:0] p1_smul_90355_comb;
  wire [31:0] p1_smul_90356_comb;
  wire [31:0] p1_smul_90357_comb;
  wire [31:0] p1_smul_90358_comb;
  wire [31:0] p1_smul_90359_comb;
  wire [31:0] p1_smul_90360_comb;
  wire [31:0] p1_smul_89807_comb;
  wire [31:0] p1_smul_89808_comb;
  wire [31:0] p1_smul_89809_comb;
  wire [31:0] p1_smul_89810_comb;
  wire [31:0] p1_smul_90361_comb;
  wire [31:0] p1_smul_90362_comb;
  wire [31:0] p1_smul_90363_comb;
  wire [31:0] p1_smul_90364_comb;
  wire [31:0] p1_smul_90365_comb;
  wire [31:0] p1_smul_90366_comb;
  wire [31:0] p1_smul_89811_comb;
  wire [31:0] p1_smul_89812_comb;
  wire [31:0] p1_smul_89813_comb;
  wire [31:0] p1_smul_89814_comb;
  wire [31:0] p1_smul_90367_comb;
  wire [31:0] p1_smul_90368_comb;
  wire [31:0] p1_smul_90369_comb;
  wire [31:0] p1_smul_90370_comb;
  wire [31:0] p1_smul_90371_comb;
  wire [31:0] p1_smul_90372_comb;
  wire [31:0] p1_smul_89815_comb;
  wire [31:0] p1_smul_89816_comb;
  wire [31:0] p1_smul_89817_comb;
  wire [31:0] p1_smul_89818_comb;
  wire [31:0] p1_smul_90373_comb;
  wire [31:0] p1_smul_90374_comb;
  wire [31:0] p1_smul_90375_comb;
  wire [31:0] p1_smul_90376_comb;
  wire [31:0] p1_smul_90377_comb;
  wire [31:0] p1_smul_90378_comb;
  wire [31:0] p1_smul_89819_comb;
  wire [31:0] p1_smul_89820_comb;
  wire [31:0] p1_smul_89821_comb;
  wire [31:0] p1_smul_89822_comb;
  wire [31:0] p1_smul_90379_comb;
  wire [31:0] p1_smul_90380_comb;
  wire [31:0] p1_smul_90381_comb;
  wire [31:0] p1_smul_90382_comb;
  wire [31:0] p1_smul_90383_comb;
  wire [31:0] p1_smul_90384_comb;
  wire [31:0] p1_smul_89823_comb;
  wire [31:0] p1_smul_89824_comb;
  wire [31:0] p1_smul_89825_comb;
  wire [31:0] p1_smul_89826_comb;
  wire [31:0] p1_smul_90385_comb;
  wire [31:0] p1_smul_90386_comb;
  wire [31:0] p1_smul_90387_comb;
  wire [31:0] p1_smul_90388_comb;
  wire [31:0] p1_smul_90389_comb;
  wire [31:0] p1_smul_90390_comb;
  wire [31:0] p1_smul_89827_comb;
  wire [31:0] p1_smul_89828_comb;
  wire [31:0] p1_smul_89829_comb;
  wire [31:0] p1_smul_89830_comb;
  wire [31:0] p1_smul_90391_comb;
  wire [31:0] p1_smul_90392_comb;
  wire [31:0] p1_smul_90393_comb;
  wire [31:0] p1_smul_90394_comb;
  wire [31:0] p1_smul_90395_comb;
  wire [31:0] p1_smul_90396_comb;
  wire [31:0] p1_smul_89831_comb;
  wire [31:0] p1_smul_89832_comb;
  wire [31:0] p1_smul_89833_comb;
  wire [31:0] p1_smul_89834_comb;
  wire [31:0] p1_smul_90397_comb;
  wire [31:0] p1_smul_90398_comb;
  wire [31:0] p1_smul_90399_comb;
  wire [31:0] p1_smul_90400_comb;
  wire [31:0] p1_smul_90401_comb;
  wire [31:0] p1_smul_90402_comb;
  wire [31:0] p1_smul_89835_comb;
  wire [31:0] p1_smul_89836_comb;
  wire [31:0] p1_smul_89837_comb;
  wire [31:0] p1_smul_89838_comb;
  wire [31:0] p1_smul_90403_comb;
  wire [31:0] p1_smul_90404_comb;
  wire [31:0] p1_smul_90405_comb;
  wire [31:0] p1_smul_90406_comb;
  wire [31:0] p1_smul_90407_comb;
  wire [31:0] p1_smul_90408_comb;
  wire [31:0] p1_smul_89839_comb;
  wire [31:0] p1_smul_89840_comb;
  wire [31:0] p1_smul_89841_comb;
  wire [31:0] p1_smul_89842_comb;
  wire [31:0] p1_smul_90409_comb;
  wire [31:0] p1_smul_90410_comb;
  wire [31:0] p1_smul_90411_comb;
  wire [31:0] p1_smul_90412_comb;
  wire [31:0] p1_smul_90413_comb;
  wire [31:0] p1_smul_90414_comb;
  wire [31:0] p1_smul_89843_comb;
  wire [31:0] p1_smul_89844_comb;
  wire [31:0] p1_smul_89845_comb;
  wire [31:0] p1_smul_89846_comb;
  wire [31:0] p1_smul_90415_comb;
  wire [31:0] p1_smul_90416_comb;
  wire [31:0] p1_smul_90417_comb;
  wire [31:0] p1_smul_90418_comb;
  wire [31:0] p1_smul_90419_comb;
  wire [31:0] p1_smul_90420_comb;
  wire [31:0] p1_smul_89847_comb;
  wire [31:0] p1_smul_89848_comb;
  wire [31:0] p1_smul_89849_comb;
  wire [31:0] p1_smul_89850_comb;
  wire [31:0] p1_smul_90421_comb;
  wire [31:0] p1_smul_90422_comb;
  wire [31:0] p1_smul_90423_comb;
  wire [31:0] p1_smul_90424_comb;
  wire [31:0] p1_smul_90425_comb;
  wire [31:0] p1_smul_90426_comb;
  wire [31:0] p1_smul_89851_comb;
  wire [31:0] p1_smul_89852_comb;
  wire [31:0] p1_smul_89853_comb;
  wire [31:0] p1_smul_89854_comb;
  wire [31:0] p1_smul_90427_comb;
  wire [31:0] p1_smul_90428_comb;
  wire [31:0] p1_smul_90429_comb;
  wire [31:0] p1_smul_90430_comb;
  wire [31:0] p1_smul_90431_comb;
  wire [31:0] p1_smul_90432_comb;
  wire [31:0] p1_smul_89855_comb;
  wire [31:0] p1_smul_89856_comb;
  wire [31:0] p1_smul_89857_comb;
  wire [31:0] p1_smul_89858_comb;
  wire [31:0] p1_smul_90433_comb;
  wire [31:0] p1_smul_90434_comb;
  wire [31:0] p1_smul_90435_comb;
  wire [31:0] p1_smul_90436_comb;
  wire [31:0] p1_smul_90437_comb;
  wire [31:0] p1_smul_90438_comb;
  wire [31:0] p1_smul_89859_comb;
  wire [31:0] p1_smul_89860_comb;
  wire [31:0] p1_smul_89861_comb;
  wire [31:0] p1_smul_89862_comb;
  wire [31:0] p1_smul_90439_comb;
  wire [31:0] p1_smul_90440_comb;
  wire [31:0] p1_smul_90441_comb;
  wire [31:0] p1_smul_90442_comb;
  wire [31:0] p1_smul_90443_comb;
  wire [31:0] p1_smul_90444_comb;
  wire [31:0] p1_smul_89863_comb;
  wire [31:0] p1_smul_89864_comb;
  wire [31:0] p1_smul_89865_comb;
  wire [31:0] p1_smul_89866_comb;
  wire [31:0] p1_smul_90445_comb;
  wire [31:0] p1_smul_90446_comb;
  wire [31:0] p1_smul_90447_comb;
  wire [31:0] p1_smul_90448_comb;
  wire [31:0] p1_smul_90449_comb;
  wire [31:0] p1_smul_90450_comb;
  wire [31:0] p1_smul_89867_comb;
  wire [31:0] p1_smul_89868_comb;
  wire [31:0] p1_smul_89869_comb;
  wire [31:0] p1_smul_89870_comb;
  wire [31:0] p1_smul_90451_comb;
  wire [31:0] p1_smul_90452_comb;
  wire [31:0] p1_smul_90453_comb;
  wire [31:0] p1_smul_90454_comb;
  wire [31:0] p1_smul_90455_comb;
  wire [31:0] p1_smul_90456_comb;
  wire [31:0] p1_smul_89871_comb;
  wire [31:0] p1_smul_89872_comb;
  wire [31:0] p1_smul_89873_comb;
  wire [31:0] p1_smul_89874_comb;
  wire [31:0] p1_smul_90457_comb;
  wire [31:0] p1_smul_90458_comb;
  wire [31:0] p1_smul_90459_comb;
  wire [31:0] p1_smul_90460_comb;
  wire [31:0] p1_smul_90461_comb;
  wire [31:0] p1_smul_90462_comb;
  wire [31:0] p1_smul_89875_comb;
  wire [31:0] p1_smul_89876_comb;
  wire [31:0] p1_smul_89877_comb;
  wire [31:0] p1_smul_89878_comb;
  wire [31:0] p1_smul_90463_comb;
  wire [31:0] p1_smul_90464_comb;
  wire [31:0] p1_smul_90465_comb;
  wire [31:0] p1_smul_90466_comb;
  wire [31:0] p1_smul_90467_comb;
  wire [31:0] p1_smul_90468_comb;
  wire [31:0] p1_smul_89879_comb;
  wire [31:0] p1_smul_89880_comb;
  wire [31:0] p1_smul_89881_comb;
  wire [31:0] p1_smul_89882_comb;
  wire [31:0] p1_smul_90469_comb;
  wire [31:0] p1_smul_90470_comb;
  wire [31:0] p1_smul_90471_comb;
  wire [31:0] p1_smul_90472_comb;
  wire [31:0] p1_smul_90473_comb;
  wire [31:0] p1_smul_90474_comb;
  wire [31:0] p1_smul_89883_comb;
  wire [31:0] p1_smul_89884_comb;
  wire [31:0] p1_smul_89885_comb;
  wire [31:0] p1_smul_89886_comb;
  wire [31:0] p1_smul_90475_comb;
  wire [31:0] p1_smul_90476_comb;
  wire [31:0] p1_smul_90477_comb;
  wire [31:0] p1_smul_90478_comb;
  wire [31:0] p1_smul_90479_comb;
  wire [31:0] p1_smul_90480_comb;
  wire [31:0] p1_smul_89887_comb;
  wire [31:0] p1_smul_89888_comb;
  wire [31:0] p1_smul_89889_comb;
  wire [31:0] p1_smul_89890_comb;
  wire [31:0] p1_smul_90481_comb;
  wire [31:0] p1_smul_90482_comb;
  wire [31:0] p1_smul_90483_comb;
  wire [31:0] p1_smul_90484_comb;
  wire [31:0] p1_smul_90485_comb;
  wire [31:0] p1_smul_90486_comb;
  wire [31:0] p1_smul_89891_comb;
  wire [31:0] p1_smul_89892_comb;
  wire [31:0] p1_smul_89893_comb;
  wire [31:0] p1_smul_89894_comb;
  wire [31:0] p1_smul_90487_comb;
  wire [31:0] p1_smul_90488_comb;
  wire [31:0] p1_smul_90489_comb;
  wire [31:0] p1_smul_90490_comb;
  wire [31:0] p1_smul_90491_comb;
  wire [31:0] p1_smul_90492_comb;
  wire [31:0] p1_smul_89895_comb;
  wire [31:0] p1_smul_89896_comb;
  wire [31:0] p1_smul_89897_comb;
  wire [31:0] p1_smul_89898_comb;
  wire [31:0] p1_smul_90493_comb;
  wire [31:0] p1_smul_90494_comb;
  wire [31:0] p1_smul_90495_comb;
  wire [31:0] p1_smul_90496_comb;
  wire [31:0] p1_smul_90497_comb;
  wire [31:0] p1_smul_90498_comb;
  assign p1_smul_89499_comb = smul32b_32b_x_32b(p0_TestBlock__A_op0, p0_TestBlock__B_op0);
  assign p1_smul_89500_comb = smul32b_32b_x_32b(p0_TestBlock__A_op1, p0_TestBlock__B_op10);
  assign p1_smul_89501_comb = smul32b_32b_x_32b(p0_TestBlock__A_op2, p0_TestBlock__B_op20);
  assign p1_smul_89502_comb = smul32b_32b_x_32b(p0_TestBlock__A_op3, p0_TestBlock__B_op30);
  assign p1_smul_89899_comb = smul32b_32b_x_32b(p0_TestBlock__A_op4, p0_TestBlock__B_op40);
  assign p1_smul_89900_comb = smul32b_32b_x_32b(p0_TestBlock__A_op5, p0_TestBlock__B_op50);
  assign p1_smul_89901_comb = smul32b_32b_x_32b(p0_TestBlock__A_op6, p0_TestBlock__B_op60);
  assign p1_smul_89902_comb = smul32b_32b_x_32b(p0_TestBlock__A_op7, p0_TestBlock__B_op70);
  assign p1_smul_89903_comb = smul32b_32b_x_32b(p0_TestBlock__A_op8, p0_TestBlock__B_op80);
  assign p1_smul_89904_comb = smul32b_32b_x_32b(p0_TestBlock__A_op9, p0_TestBlock__B_op90);
  assign p1_smul_89503_comb = smul32b_32b_x_32b(p0_TestBlock__A_op0, p0_TestBlock__B_op1);
  assign p1_smul_89504_comb = smul32b_32b_x_32b(p0_TestBlock__A_op1, p0_TestBlock__B_op11);
  assign p1_smul_89505_comb = smul32b_32b_x_32b(p0_TestBlock__A_op2, p0_TestBlock__B_op21);
  assign p1_smul_89506_comb = smul32b_32b_x_32b(p0_TestBlock__A_op3, p0_TestBlock__B_op31);
  assign p1_smul_89905_comb = smul32b_32b_x_32b(p0_TestBlock__A_op4, p0_TestBlock__B_op41);
  assign p1_smul_89906_comb = smul32b_32b_x_32b(p0_TestBlock__A_op5, p0_TestBlock__B_op51);
  assign p1_smul_89907_comb = smul32b_32b_x_32b(p0_TestBlock__A_op6, p0_TestBlock__B_op61);
  assign p1_smul_89908_comb = smul32b_32b_x_32b(p0_TestBlock__A_op7, p0_TestBlock__B_op71);
  assign p1_smul_89909_comb = smul32b_32b_x_32b(p0_TestBlock__A_op8, p0_TestBlock__B_op81);
  assign p1_smul_89910_comb = smul32b_32b_x_32b(p0_TestBlock__A_op9, p0_TestBlock__B_op91);
  assign p1_smul_89507_comb = smul32b_32b_x_32b(p0_TestBlock__A_op0, p0_TestBlock__B_op2);
  assign p1_smul_89508_comb = smul32b_32b_x_32b(p0_TestBlock__A_op1, p0_TestBlock__B_op12);
  assign p1_smul_89509_comb = smul32b_32b_x_32b(p0_TestBlock__A_op2, p0_TestBlock__B_op22);
  assign p1_smul_89510_comb = smul32b_32b_x_32b(p0_TestBlock__A_op3, p0_TestBlock__B_op32);
  assign p1_smul_89911_comb = smul32b_32b_x_32b(p0_TestBlock__A_op4, p0_TestBlock__B_op42);
  assign p1_smul_89912_comb = smul32b_32b_x_32b(p0_TestBlock__A_op5, p0_TestBlock__B_op52);
  assign p1_smul_89913_comb = smul32b_32b_x_32b(p0_TestBlock__A_op6, p0_TestBlock__B_op62);
  assign p1_smul_89914_comb = smul32b_32b_x_32b(p0_TestBlock__A_op7, p0_TestBlock__B_op72);
  assign p1_smul_89915_comb = smul32b_32b_x_32b(p0_TestBlock__A_op8, p0_TestBlock__B_op82);
  assign p1_smul_89916_comb = smul32b_32b_x_32b(p0_TestBlock__A_op9, p0_TestBlock__B_op92);
  assign p1_smul_89511_comb = smul32b_32b_x_32b(p0_TestBlock__A_op0, p0_TestBlock__B_op3);
  assign p1_smul_89512_comb = smul32b_32b_x_32b(p0_TestBlock__A_op1, p0_TestBlock__B_op13);
  assign p1_smul_89513_comb = smul32b_32b_x_32b(p0_TestBlock__A_op2, p0_TestBlock__B_op23);
  assign p1_smul_89514_comb = smul32b_32b_x_32b(p0_TestBlock__A_op3, p0_TestBlock__B_op33);
  assign p1_smul_89917_comb = smul32b_32b_x_32b(p0_TestBlock__A_op4, p0_TestBlock__B_op43);
  assign p1_smul_89918_comb = smul32b_32b_x_32b(p0_TestBlock__A_op5, p0_TestBlock__B_op53);
  assign p1_smul_89919_comb = smul32b_32b_x_32b(p0_TestBlock__A_op6, p0_TestBlock__B_op63);
  assign p1_smul_89920_comb = smul32b_32b_x_32b(p0_TestBlock__A_op7, p0_TestBlock__B_op73);
  assign p1_smul_89921_comb = smul32b_32b_x_32b(p0_TestBlock__A_op8, p0_TestBlock__B_op83);
  assign p1_smul_89922_comb = smul32b_32b_x_32b(p0_TestBlock__A_op9, p0_TestBlock__B_op93);
  assign p1_smul_89515_comb = smul32b_32b_x_32b(p0_TestBlock__A_op0, p0_TestBlock__B_op4);
  assign p1_smul_89516_comb = smul32b_32b_x_32b(p0_TestBlock__A_op1, p0_TestBlock__B_op14);
  assign p1_smul_89517_comb = smul32b_32b_x_32b(p0_TestBlock__A_op2, p0_TestBlock__B_op24);
  assign p1_smul_89518_comb = smul32b_32b_x_32b(p0_TestBlock__A_op3, p0_TestBlock__B_op34);
  assign p1_smul_89923_comb = smul32b_32b_x_32b(p0_TestBlock__A_op4, p0_TestBlock__B_op44);
  assign p1_smul_89924_comb = smul32b_32b_x_32b(p0_TestBlock__A_op5, p0_TestBlock__B_op54);
  assign p1_smul_89925_comb = smul32b_32b_x_32b(p0_TestBlock__A_op6, p0_TestBlock__B_op64);
  assign p1_smul_89926_comb = smul32b_32b_x_32b(p0_TestBlock__A_op7, p0_TestBlock__B_op74);
  assign p1_smul_89927_comb = smul32b_32b_x_32b(p0_TestBlock__A_op8, p0_TestBlock__B_op84);
  assign p1_smul_89928_comb = smul32b_32b_x_32b(p0_TestBlock__A_op9, p0_TestBlock__B_op94);
  assign p1_smul_89519_comb = smul32b_32b_x_32b(p0_TestBlock__A_op0, p0_TestBlock__B_op5);
  assign p1_smul_89520_comb = smul32b_32b_x_32b(p0_TestBlock__A_op1, p0_TestBlock__B_op15);
  assign p1_smul_89521_comb = smul32b_32b_x_32b(p0_TestBlock__A_op2, p0_TestBlock__B_op25);
  assign p1_smul_89522_comb = smul32b_32b_x_32b(p0_TestBlock__A_op3, p0_TestBlock__B_op35);
  assign p1_smul_89929_comb = smul32b_32b_x_32b(p0_TestBlock__A_op4, p0_TestBlock__B_op45);
  assign p1_smul_89930_comb = smul32b_32b_x_32b(p0_TestBlock__A_op5, p0_TestBlock__B_op55);
  assign p1_smul_89931_comb = smul32b_32b_x_32b(p0_TestBlock__A_op6, p0_TestBlock__B_op65);
  assign p1_smul_89932_comb = smul32b_32b_x_32b(p0_TestBlock__A_op7, p0_TestBlock__B_op75);
  assign p1_smul_89933_comb = smul32b_32b_x_32b(p0_TestBlock__A_op8, p0_TestBlock__B_op85);
  assign p1_smul_89934_comb = smul32b_32b_x_32b(p0_TestBlock__A_op9, p0_TestBlock__B_op95);
  assign p1_smul_89523_comb = smul32b_32b_x_32b(p0_TestBlock__A_op0, p0_TestBlock__B_op6);
  assign p1_smul_89524_comb = smul32b_32b_x_32b(p0_TestBlock__A_op1, p0_TestBlock__B_op16);
  assign p1_smul_89525_comb = smul32b_32b_x_32b(p0_TestBlock__A_op2, p0_TestBlock__B_op26);
  assign p1_smul_89526_comb = smul32b_32b_x_32b(p0_TestBlock__A_op3, p0_TestBlock__B_op36);
  assign p1_smul_89935_comb = smul32b_32b_x_32b(p0_TestBlock__A_op4, p0_TestBlock__B_op46);
  assign p1_smul_89936_comb = smul32b_32b_x_32b(p0_TestBlock__A_op5, p0_TestBlock__B_op56);
  assign p1_smul_89937_comb = smul32b_32b_x_32b(p0_TestBlock__A_op6, p0_TestBlock__B_op66);
  assign p1_smul_89938_comb = smul32b_32b_x_32b(p0_TestBlock__A_op7, p0_TestBlock__B_op76);
  assign p1_smul_89939_comb = smul32b_32b_x_32b(p0_TestBlock__A_op8, p0_TestBlock__B_op86);
  assign p1_smul_89940_comb = smul32b_32b_x_32b(p0_TestBlock__A_op9, p0_TestBlock__B_op96);
  assign p1_smul_89527_comb = smul32b_32b_x_32b(p0_TestBlock__A_op0, p0_TestBlock__B_op7);
  assign p1_smul_89528_comb = smul32b_32b_x_32b(p0_TestBlock__A_op1, p0_TestBlock__B_op17);
  assign p1_smul_89529_comb = smul32b_32b_x_32b(p0_TestBlock__A_op2, p0_TestBlock__B_op27);
  assign p1_smul_89530_comb = smul32b_32b_x_32b(p0_TestBlock__A_op3, p0_TestBlock__B_op37);
  assign p1_smul_89941_comb = smul32b_32b_x_32b(p0_TestBlock__A_op4, p0_TestBlock__B_op47);
  assign p1_smul_89942_comb = smul32b_32b_x_32b(p0_TestBlock__A_op5, p0_TestBlock__B_op57);
  assign p1_smul_89943_comb = smul32b_32b_x_32b(p0_TestBlock__A_op6, p0_TestBlock__B_op67);
  assign p1_smul_89944_comb = smul32b_32b_x_32b(p0_TestBlock__A_op7, p0_TestBlock__B_op77);
  assign p1_smul_89945_comb = smul32b_32b_x_32b(p0_TestBlock__A_op8, p0_TestBlock__B_op87);
  assign p1_smul_89946_comb = smul32b_32b_x_32b(p0_TestBlock__A_op9, p0_TestBlock__B_op97);
  assign p1_smul_89531_comb = smul32b_32b_x_32b(p0_TestBlock__A_op0, p0_TestBlock__B_op8);
  assign p1_smul_89532_comb = smul32b_32b_x_32b(p0_TestBlock__A_op1, p0_TestBlock__B_op18);
  assign p1_smul_89533_comb = smul32b_32b_x_32b(p0_TestBlock__A_op2, p0_TestBlock__B_op28);
  assign p1_smul_89534_comb = smul32b_32b_x_32b(p0_TestBlock__A_op3, p0_TestBlock__B_op38);
  assign p1_smul_89947_comb = smul32b_32b_x_32b(p0_TestBlock__A_op4, p0_TestBlock__B_op48);
  assign p1_smul_89948_comb = smul32b_32b_x_32b(p0_TestBlock__A_op5, p0_TestBlock__B_op58);
  assign p1_smul_89949_comb = smul32b_32b_x_32b(p0_TestBlock__A_op6, p0_TestBlock__B_op68);
  assign p1_smul_89950_comb = smul32b_32b_x_32b(p0_TestBlock__A_op7, p0_TestBlock__B_op78);
  assign p1_smul_89951_comb = smul32b_32b_x_32b(p0_TestBlock__A_op8, p0_TestBlock__B_op88);
  assign p1_smul_89952_comb = smul32b_32b_x_32b(p0_TestBlock__A_op9, p0_TestBlock__B_op98);
  assign p1_smul_89535_comb = smul32b_32b_x_32b(p0_TestBlock__A_op0, p0_TestBlock__B_op9);
  assign p1_smul_89536_comb = smul32b_32b_x_32b(p0_TestBlock__A_op1, p0_TestBlock__B_op19);
  assign p1_smul_89537_comb = smul32b_32b_x_32b(p0_TestBlock__A_op2, p0_TestBlock__B_op29);
  assign p1_smul_89538_comb = smul32b_32b_x_32b(p0_TestBlock__A_op3, p0_TestBlock__B_op39);
  assign p1_smul_89953_comb = smul32b_32b_x_32b(p0_TestBlock__A_op4, p0_TestBlock__B_op49);
  assign p1_smul_89954_comb = smul32b_32b_x_32b(p0_TestBlock__A_op5, p0_TestBlock__B_op59);
  assign p1_smul_89955_comb = smul32b_32b_x_32b(p0_TestBlock__A_op6, p0_TestBlock__B_op69);
  assign p1_smul_89956_comb = smul32b_32b_x_32b(p0_TestBlock__A_op7, p0_TestBlock__B_op79);
  assign p1_smul_89957_comb = smul32b_32b_x_32b(p0_TestBlock__A_op8, p0_TestBlock__B_op89);
  assign p1_smul_89958_comb = smul32b_32b_x_32b(p0_TestBlock__A_op9, p0_TestBlock__B_op99);
  assign p1_smul_89539_comb = smul32b_32b_x_32b(p0_TestBlock__A_op10, p0_TestBlock__B_op0);
  assign p1_smul_89540_comb = smul32b_32b_x_32b(p0_TestBlock__A_op11, p0_TestBlock__B_op10);
  assign p1_smul_89541_comb = smul32b_32b_x_32b(p0_TestBlock__A_op12, p0_TestBlock__B_op20);
  assign p1_smul_89542_comb = smul32b_32b_x_32b(p0_TestBlock__A_op13, p0_TestBlock__B_op30);
  assign p1_smul_89959_comb = smul32b_32b_x_32b(p0_TestBlock__A_op14, p0_TestBlock__B_op40);
  assign p1_smul_89960_comb = smul32b_32b_x_32b(p0_TestBlock__A_op15, p0_TestBlock__B_op50);
  assign p1_smul_89961_comb = smul32b_32b_x_32b(p0_TestBlock__A_op16, p0_TestBlock__B_op60);
  assign p1_smul_89962_comb = smul32b_32b_x_32b(p0_TestBlock__A_op17, p0_TestBlock__B_op70);
  assign p1_smul_89963_comb = smul32b_32b_x_32b(p0_TestBlock__A_op18, p0_TestBlock__B_op80);
  assign p1_smul_89964_comb = smul32b_32b_x_32b(p0_TestBlock__A_op19, p0_TestBlock__B_op90);
  assign p1_smul_89543_comb = smul32b_32b_x_32b(p0_TestBlock__A_op10, p0_TestBlock__B_op1);
  assign p1_smul_89544_comb = smul32b_32b_x_32b(p0_TestBlock__A_op11, p0_TestBlock__B_op11);
  assign p1_smul_89545_comb = smul32b_32b_x_32b(p0_TestBlock__A_op12, p0_TestBlock__B_op21);
  assign p1_smul_89546_comb = smul32b_32b_x_32b(p0_TestBlock__A_op13, p0_TestBlock__B_op31);
  assign p1_smul_89965_comb = smul32b_32b_x_32b(p0_TestBlock__A_op14, p0_TestBlock__B_op41);
  assign p1_smul_89966_comb = smul32b_32b_x_32b(p0_TestBlock__A_op15, p0_TestBlock__B_op51);
  assign p1_smul_89967_comb = smul32b_32b_x_32b(p0_TestBlock__A_op16, p0_TestBlock__B_op61);
  assign p1_smul_89968_comb = smul32b_32b_x_32b(p0_TestBlock__A_op17, p0_TestBlock__B_op71);
  assign p1_smul_89969_comb = smul32b_32b_x_32b(p0_TestBlock__A_op18, p0_TestBlock__B_op81);
  assign p1_smul_89970_comb = smul32b_32b_x_32b(p0_TestBlock__A_op19, p0_TestBlock__B_op91);
  assign p1_smul_89547_comb = smul32b_32b_x_32b(p0_TestBlock__A_op10, p0_TestBlock__B_op2);
  assign p1_smul_89548_comb = smul32b_32b_x_32b(p0_TestBlock__A_op11, p0_TestBlock__B_op12);
  assign p1_smul_89549_comb = smul32b_32b_x_32b(p0_TestBlock__A_op12, p0_TestBlock__B_op22);
  assign p1_smul_89550_comb = smul32b_32b_x_32b(p0_TestBlock__A_op13, p0_TestBlock__B_op32);
  assign p1_smul_89971_comb = smul32b_32b_x_32b(p0_TestBlock__A_op14, p0_TestBlock__B_op42);
  assign p1_smul_89972_comb = smul32b_32b_x_32b(p0_TestBlock__A_op15, p0_TestBlock__B_op52);
  assign p1_smul_89973_comb = smul32b_32b_x_32b(p0_TestBlock__A_op16, p0_TestBlock__B_op62);
  assign p1_smul_89974_comb = smul32b_32b_x_32b(p0_TestBlock__A_op17, p0_TestBlock__B_op72);
  assign p1_smul_89975_comb = smul32b_32b_x_32b(p0_TestBlock__A_op18, p0_TestBlock__B_op82);
  assign p1_smul_89976_comb = smul32b_32b_x_32b(p0_TestBlock__A_op19, p0_TestBlock__B_op92);
  assign p1_smul_89551_comb = smul32b_32b_x_32b(p0_TestBlock__A_op10, p0_TestBlock__B_op3);
  assign p1_smul_89552_comb = smul32b_32b_x_32b(p0_TestBlock__A_op11, p0_TestBlock__B_op13);
  assign p1_smul_89553_comb = smul32b_32b_x_32b(p0_TestBlock__A_op12, p0_TestBlock__B_op23);
  assign p1_smul_89554_comb = smul32b_32b_x_32b(p0_TestBlock__A_op13, p0_TestBlock__B_op33);
  assign p1_smul_89977_comb = smul32b_32b_x_32b(p0_TestBlock__A_op14, p0_TestBlock__B_op43);
  assign p1_smul_89978_comb = smul32b_32b_x_32b(p0_TestBlock__A_op15, p0_TestBlock__B_op53);
  assign p1_smul_89979_comb = smul32b_32b_x_32b(p0_TestBlock__A_op16, p0_TestBlock__B_op63);
  assign p1_smul_89980_comb = smul32b_32b_x_32b(p0_TestBlock__A_op17, p0_TestBlock__B_op73);
  assign p1_smul_89981_comb = smul32b_32b_x_32b(p0_TestBlock__A_op18, p0_TestBlock__B_op83);
  assign p1_smul_89982_comb = smul32b_32b_x_32b(p0_TestBlock__A_op19, p0_TestBlock__B_op93);
  assign p1_smul_89555_comb = smul32b_32b_x_32b(p0_TestBlock__A_op10, p0_TestBlock__B_op4);
  assign p1_smul_89556_comb = smul32b_32b_x_32b(p0_TestBlock__A_op11, p0_TestBlock__B_op14);
  assign p1_smul_89557_comb = smul32b_32b_x_32b(p0_TestBlock__A_op12, p0_TestBlock__B_op24);
  assign p1_smul_89558_comb = smul32b_32b_x_32b(p0_TestBlock__A_op13, p0_TestBlock__B_op34);
  assign p1_smul_89983_comb = smul32b_32b_x_32b(p0_TestBlock__A_op14, p0_TestBlock__B_op44);
  assign p1_smul_89984_comb = smul32b_32b_x_32b(p0_TestBlock__A_op15, p0_TestBlock__B_op54);
  assign p1_smul_89985_comb = smul32b_32b_x_32b(p0_TestBlock__A_op16, p0_TestBlock__B_op64);
  assign p1_smul_89986_comb = smul32b_32b_x_32b(p0_TestBlock__A_op17, p0_TestBlock__B_op74);
  assign p1_smul_89987_comb = smul32b_32b_x_32b(p0_TestBlock__A_op18, p0_TestBlock__B_op84);
  assign p1_smul_89988_comb = smul32b_32b_x_32b(p0_TestBlock__A_op19, p0_TestBlock__B_op94);
  assign p1_smul_89559_comb = smul32b_32b_x_32b(p0_TestBlock__A_op10, p0_TestBlock__B_op5);
  assign p1_smul_89560_comb = smul32b_32b_x_32b(p0_TestBlock__A_op11, p0_TestBlock__B_op15);
  assign p1_smul_89561_comb = smul32b_32b_x_32b(p0_TestBlock__A_op12, p0_TestBlock__B_op25);
  assign p1_smul_89562_comb = smul32b_32b_x_32b(p0_TestBlock__A_op13, p0_TestBlock__B_op35);
  assign p1_smul_89989_comb = smul32b_32b_x_32b(p0_TestBlock__A_op14, p0_TestBlock__B_op45);
  assign p1_smul_89990_comb = smul32b_32b_x_32b(p0_TestBlock__A_op15, p0_TestBlock__B_op55);
  assign p1_smul_89991_comb = smul32b_32b_x_32b(p0_TestBlock__A_op16, p0_TestBlock__B_op65);
  assign p1_smul_89992_comb = smul32b_32b_x_32b(p0_TestBlock__A_op17, p0_TestBlock__B_op75);
  assign p1_smul_89993_comb = smul32b_32b_x_32b(p0_TestBlock__A_op18, p0_TestBlock__B_op85);
  assign p1_smul_89994_comb = smul32b_32b_x_32b(p0_TestBlock__A_op19, p0_TestBlock__B_op95);
  assign p1_smul_89563_comb = smul32b_32b_x_32b(p0_TestBlock__A_op10, p0_TestBlock__B_op6);
  assign p1_smul_89564_comb = smul32b_32b_x_32b(p0_TestBlock__A_op11, p0_TestBlock__B_op16);
  assign p1_smul_89565_comb = smul32b_32b_x_32b(p0_TestBlock__A_op12, p0_TestBlock__B_op26);
  assign p1_smul_89566_comb = smul32b_32b_x_32b(p0_TestBlock__A_op13, p0_TestBlock__B_op36);
  assign p1_smul_89995_comb = smul32b_32b_x_32b(p0_TestBlock__A_op14, p0_TestBlock__B_op46);
  assign p1_smul_89996_comb = smul32b_32b_x_32b(p0_TestBlock__A_op15, p0_TestBlock__B_op56);
  assign p1_smul_89997_comb = smul32b_32b_x_32b(p0_TestBlock__A_op16, p0_TestBlock__B_op66);
  assign p1_smul_89998_comb = smul32b_32b_x_32b(p0_TestBlock__A_op17, p0_TestBlock__B_op76);
  assign p1_smul_89999_comb = smul32b_32b_x_32b(p0_TestBlock__A_op18, p0_TestBlock__B_op86);
  assign p1_smul_90000_comb = smul32b_32b_x_32b(p0_TestBlock__A_op19, p0_TestBlock__B_op96);
  assign p1_smul_89567_comb = smul32b_32b_x_32b(p0_TestBlock__A_op10, p0_TestBlock__B_op7);
  assign p1_smul_89568_comb = smul32b_32b_x_32b(p0_TestBlock__A_op11, p0_TestBlock__B_op17);
  assign p1_smul_89569_comb = smul32b_32b_x_32b(p0_TestBlock__A_op12, p0_TestBlock__B_op27);
  assign p1_smul_89570_comb = smul32b_32b_x_32b(p0_TestBlock__A_op13, p0_TestBlock__B_op37);
  assign p1_smul_90001_comb = smul32b_32b_x_32b(p0_TestBlock__A_op14, p0_TestBlock__B_op47);
  assign p1_smul_90002_comb = smul32b_32b_x_32b(p0_TestBlock__A_op15, p0_TestBlock__B_op57);
  assign p1_smul_90003_comb = smul32b_32b_x_32b(p0_TestBlock__A_op16, p0_TestBlock__B_op67);
  assign p1_smul_90004_comb = smul32b_32b_x_32b(p0_TestBlock__A_op17, p0_TestBlock__B_op77);
  assign p1_smul_90005_comb = smul32b_32b_x_32b(p0_TestBlock__A_op18, p0_TestBlock__B_op87);
  assign p1_smul_90006_comb = smul32b_32b_x_32b(p0_TestBlock__A_op19, p0_TestBlock__B_op97);
  assign p1_smul_89571_comb = smul32b_32b_x_32b(p0_TestBlock__A_op10, p0_TestBlock__B_op8);
  assign p1_smul_89572_comb = smul32b_32b_x_32b(p0_TestBlock__A_op11, p0_TestBlock__B_op18);
  assign p1_smul_89573_comb = smul32b_32b_x_32b(p0_TestBlock__A_op12, p0_TestBlock__B_op28);
  assign p1_smul_89574_comb = smul32b_32b_x_32b(p0_TestBlock__A_op13, p0_TestBlock__B_op38);
  assign p1_smul_90007_comb = smul32b_32b_x_32b(p0_TestBlock__A_op14, p0_TestBlock__B_op48);
  assign p1_smul_90008_comb = smul32b_32b_x_32b(p0_TestBlock__A_op15, p0_TestBlock__B_op58);
  assign p1_smul_90009_comb = smul32b_32b_x_32b(p0_TestBlock__A_op16, p0_TestBlock__B_op68);
  assign p1_smul_90010_comb = smul32b_32b_x_32b(p0_TestBlock__A_op17, p0_TestBlock__B_op78);
  assign p1_smul_90011_comb = smul32b_32b_x_32b(p0_TestBlock__A_op18, p0_TestBlock__B_op88);
  assign p1_smul_90012_comb = smul32b_32b_x_32b(p0_TestBlock__A_op19, p0_TestBlock__B_op98);
  assign p1_smul_89575_comb = smul32b_32b_x_32b(p0_TestBlock__A_op10, p0_TestBlock__B_op9);
  assign p1_smul_89576_comb = smul32b_32b_x_32b(p0_TestBlock__A_op11, p0_TestBlock__B_op19);
  assign p1_smul_89577_comb = smul32b_32b_x_32b(p0_TestBlock__A_op12, p0_TestBlock__B_op29);
  assign p1_smul_89578_comb = smul32b_32b_x_32b(p0_TestBlock__A_op13, p0_TestBlock__B_op39);
  assign p1_smul_90013_comb = smul32b_32b_x_32b(p0_TestBlock__A_op14, p0_TestBlock__B_op49);
  assign p1_smul_90014_comb = smul32b_32b_x_32b(p0_TestBlock__A_op15, p0_TestBlock__B_op59);
  assign p1_smul_90015_comb = smul32b_32b_x_32b(p0_TestBlock__A_op16, p0_TestBlock__B_op69);
  assign p1_smul_90016_comb = smul32b_32b_x_32b(p0_TestBlock__A_op17, p0_TestBlock__B_op79);
  assign p1_smul_90017_comb = smul32b_32b_x_32b(p0_TestBlock__A_op18, p0_TestBlock__B_op89);
  assign p1_smul_90018_comb = smul32b_32b_x_32b(p0_TestBlock__A_op19, p0_TestBlock__B_op99);
  assign p1_smul_89579_comb = smul32b_32b_x_32b(p0_TestBlock__A_op20, p0_TestBlock__B_op0);
  assign p1_smul_89580_comb = smul32b_32b_x_32b(p0_TestBlock__A_op21, p0_TestBlock__B_op10);
  assign p1_smul_89581_comb = smul32b_32b_x_32b(p0_TestBlock__A_op22, p0_TestBlock__B_op20);
  assign p1_smul_89582_comb = smul32b_32b_x_32b(p0_TestBlock__A_op23, p0_TestBlock__B_op30);
  assign p1_smul_90019_comb = smul32b_32b_x_32b(p0_TestBlock__A_op24, p0_TestBlock__B_op40);
  assign p1_smul_90020_comb = smul32b_32b_x_32b(p0_TestBlock__A_op25, p0_TestBlock__B_op50);
  assign p1_smul_90021_comb = smul32b_32b_x_32b(p0_TestBlock__A_op26, p0_TestBlock__B_op60);
  assign p1_smul_90022_comb = smul32b_32b_x_32b(p0_TestBlock__A_op27, p0_TestBlock__B_op70);
  assign p1_smul_90023_comb = smul32b_32b_x_32b(p0_TestBlock__A_op28, p0_TestBlock__B_op80);
  assign p1_smul_90024_comb = smul32b_32b_x_32b(p0_TestBlock__A_op29, p0_TestBlock__B_op90);
  assign p1_smul_89583_comb = smul32b_32b_x_32b(p0_TestBlock__A_op20, p0_TestBlock__B_op1);
  assign p1_smul_89584_comb = smul32b_32b_x_32b(p0_TestBlock__A_op21, p0_TestBlock__B_op11);
  assign p1_smul_89585_comb = smul32b_32b_x_32b(p0_TestBlock__A_op22, p0_TestBlock__B_op21);
  assign p1_smul_89586_comb = smul32b_32b_x_32b(p0_TestBlock__A_op23, p0_TestBlock__B_op31);
  assign p1_smul_90025_comb = smul32b_32b_x_32b(p0_TestBlock__A_op24, p0_TestBlock__B_op41);
  assign p1_smul_90026_comb = smul32b_32b_x_32b(p0_TestBlock__A_op25, p0_TestBlock__B_op51);
  assign p1_smul_90027_comb = smul32b_32b_x_32b(p0_TestBlock__A_op26, p0_TestBlock__B_op61);
  assign p1_smul_90028_comb = smul32b_32b_x_32b(p0_TestBlock__A_op27, p0_TestBlock__B_op71);
  assign p1_smul_90029_comb = smul32b_32b_x_32b(p0_TestBlock__A_op28, p0_TestBlock__B_op81);
  assign p1_smul_90030_comb = smul32b_32b_x_32b(p0_TestBlock__A_op29, p0_TestBlock__B_op91);
  assign p1_smul_89587_comb = smul32b_32b_x_32b(p0_TestBlock__A_op20, p0_TestBlock__B_op2);
  assign p1_smul_89588_comb = smul32b_32b_x_32b(p0_TestBlock__A_op21, p0_TestBlock__B_op12);
  assign p1_smul_89589_comb = smul32b_32b_x_32b(p0_TestBlock__A_op22, p0_TestBlock__B_op22);
  assign p1_smul_89590_comb = smul32b_32b_x_32b(p0_TestBlock__A_op23, p0_TestBlock__B_op32);
  assign p1_smul_90031_comb = smul32b_32b_x_32b(p0_TestBlock__A_op24, p0_TestBlock__B_op42);
  assign p1_smul_90032_comb = smul32b_32b_x_32b(p0_TestBlock__A_op25, p0_TestBlock__B_op52);
  assign p1_smul_90033_comb = smul32b_32b_x_32b(p0_TestBlock__A_op26, p0_TestBlock__B_op62);
  assign p1_smul_90034_comb = smul32b_32b_x_32b(p0_TestBlock__A_op27, p0_TestBlock__B_op72);
  assign p1_smul_90035_comb = smul32b_32b_x_32b(p0_TestBlock__A_op28, p0_TestBlock__B_op82);
  assign p1_smul_90036_comb = smul32b_32b_x_32b(p0_TestBlock__A_op29, p0_TestBlock__B_op92);
  assign p1_smul_89591_comb = smul32b_32b_x_32b(p0_TestBlock__A_op20, p0_TestBlock__B_op3);
  assign p1_smul_89592_comb = smul32b_32b_x_32b(p0_TestBlock__A_op21, p0_TestBlock__B_op13);
  assign p1_smul_89593_comb = smul32b_32b_x_32b(p0_TestBlock__A_op22, p0_TestBlock__B_op23);
  assign p1_smul_89594_comb = smul32b_32b_x_32b(p0_TestBlock__A_op23, p0_TestBlock__B_op33);
  assign p1_smul_90037_comb = smul32b_32b_x_32b(p0_TestBlock__A_op24, p0_TestBlock__B_op43);
  assign p1_smul_90038_comb = smul32b_32b_x_32b(p0_TestBlock__A_op25, p0_TestBlock__B_op53);
  assign p1_smul_90039_comb = smul32b_32b_x_32b(p0_TestBlock__A_op26, p0_TestBlock__B_op63);
  assign p1_smul_90040_comb = smul32b_32b_x_32b(p0_TestBlock__A_op27, p0_TestBlock__B_op73);
  assign p1_smul_90041_comb = smul32b_32b_x_32b(p0_TestBlock__A_op28, p0_TestBlock__B_op83);
  assign p1_smul_90042_comb = smul32b_32b_x_32b(p0_TestBlock__A_op29, p0_TestBlock__B_op93);
  assign p1_smul_89595_comb = smul32b_32b_x_32b(p0_TestBlock__A_op20, p0_TestBlock__B_op4);
  assign p1_smul_89596_comb = smul32b_32b_x_32b(p0_TestBlock__A_op21, p0_TestBlock__B_op14);
  assign p1_smul_89597_comb = smul32b_32b_x_32b(p0_TestBlock__A_op22, p0_TestBlock__B_op24);
  assign p1_smul_89598_comb = smul32b_32b_x_32b(p0_TestBlock__A_op23, p0_TestBlock__B_op34);
  assign p1_smul_90043_comb = smul32b_32b_x_32b(p0_TestBlock__A_op24, p0_TestBlock__B_op44);
  assign p1_smul_90044_comb = smul32b_32b_x_32b(p0_TestBlock__A_op25, p0_TestBlock__B_op54);
  assign p1_smul_90045_comb = smul32b_32b_x_32b(p0_TestBlock__A_op26, p0_TestBlock__B_op64);
  assign p1_smul_90046_comb = smul32b_32b_x_32b(p0_TestBlock__A_op27, p0_TestBlock__B_op74);
  assign p1_smul_90047_comb = smul32b_32b_x_32b(p0_TestBlock__A_op28, p0_TestBlock__B_op84);
  assign p1_smul_90048_comb = smul32b_32b_x_32b(p0_TestBlock__A_op29, p0_TestBlock__B_op94);
  assign p1_smul_89599_comb = smul32b_32b_x_32b(p0_TestBlock__A_op20, p0_TestBlock__B_op5);
  assign p1_smul_89600_comb = smul32b_32b_x_32b(p0_TestBlock__A_op21, p0_TestBlock__B_op15);
  assign p1_smul_89601_comb = smul32b_32b_x_32b(p0_TestBlock__A_op22, p0_TestBlock__B_op25);
  assign p1_smul_89602_comb = smul32b_32b_x_32b(p0_TestBlock__A_op23, p0_TestBlock__B_op35);
  assign p1_smul_90049_comb = smul32b_32b_x_32b(p0_TestBlock__A_op24, p0_TestBlock__B_op45);
  assign p1_smul_90050_comb = smul32b_32b_x_32b(p0_TestBlock__A_op25, p0_TestBlock__B_op55);
  assign p1_smul_90051_comb = smul32b_32b_x_32b(p0_TestBlock__A_op26, p0_TestBlock__B_op65);
  assign p1_smul_90052_comb = smul32b_32b_x_32b(p0_TestBlock__A_op27, p0_TestBlock__B_op75);
  assign p1_smul_90053_comb = smul32b_32b_x_32b(p0_TestBlock__A_op28, p0_TestBlock__B_op85);
  assign p1_smul_90054_comb = smul32b_32b_x_32b(p0_TestBlock__A_op29, p0_TestBlock__B_op95);
  assign p1_smul_89603_comb = smul32b_32b_x_32b(p0_TestBlock__A_op20, p0_TestBlock__B_op6);
  assign p1_smul_89604_comb = smul32b_32b_x_32b(p0_TestBlock__A_op21, p0_TestBlock__B_op16);
  assign p1_smul_89605_comb = smul32b_32b_x_32b(p0_TestBlock__A_op22, p0_TestBlock__B_op26);
  assign p1_smul_89606_comb = smul32b_32b_x_32b(p0_TestBlock__A_op23, p0_TestBlock__B_op36);
  assign p1_smul_90055_comb = smul32b_32b_x_32b(p0_TestBlock__A_op24, p0_TestBlock__B_op46);
  assign p1_smul_90056_comb = smul32b_32b_x_32b(p0_TestBlock__A_op25, p0_TestBlock__B_op56);
  assign p1_smul_90057_comb = smul32b_32b_x_32b(p0_TestBlock__A_op26, p0_TestBlock__B_op66);
  assign p1_smul_90058_comb = smul32b_32b_x_32b(p0_TestBlock__A_op27, p0_TestBlock__B_op76);
  assign p1_smul_90059_comb = smul32b_32b_x_32b(p0_TestBlock__A_op28, p0_TestBlock__B_op86);
  assign p1_smul_90060_comb = smul32b_32b_x_32b(p0_TestBlock__A_op29, p0_TestBlock__B_op96);
  assign p1_smul_89607_comb = smul32b_32b_x_32b(p0_TestBlock__A_op20, p0_TestBlock__B_op7);
  assign p1_smul_89608_comb = smul32b_32b_x_32b(p0_TestBlock__A_op21, p0_TestBlock__B_op17);
  assign p1_smul_89609_comb = smul32b_32b_x_32b(p0_TestBlock__A_op22, p0_TestBlock__B_op27);
  assign p1_smul_89610_comb = smul32b_32b_x_32b(p0_TestBlock__A_op23, p0_TestBlock__B_op37);
  assign p1_smul_90061_comb = smul32b_32b_x_32b(p0_TestBlock__A_op24, p0_TestBlock__B_op47);
  assign p1_smul_90062_comb = smul32b_32b_x_32b(p0_TestBlock__A_op25, p0_TestBlock__B_op57);
  assign p1_smul_90063_comb = smul32b_32b_x_32b(p0_TestBlock__A_op26, p0_TestBlock__B_op67);
  assign p1_smul_90064_comb = smul32b_32b_x_32b(p0_TestBlock__A_op27, p0_TestBlock__B_op77);
  assign p1_smul_90065_comb = smul32b_32b_x_32b(p0_TestBlock__A_op28, p0_TestBlock__B_op87);
  assign p1_smul_90066_comb = smul32b_32b_x_32b(p0_TestBlock__A_op29, p0_TestBlock__B_op97);
  assign p1_smul_89611_comb = smul32b_32b_x_32b(p0_TestBlock__A_op20, p0_TestBlock__B_op8);
  assign p1_smul_89612_comb = smul32b_32b_x_32b(p0_TestBlock__A_op21, p0_TestBlock__B_op18);
  assign p1_smul_89613_comb = smul32b_32b_x_32b(p0_TestBlock__A_op22, p0_TestBlock__B_op28);
  assign p1_smul_89614_comb = smul32b_32b_x_32b(p0_TestBlock__A_op23, p0_TestBlock__B_op38);
  assign p1_smul_90067_comb = smul32b_32b_x_32b(p0_TestBlock__A_op24, p0_TestBlock__B_op48);
  assign p1_smul_90068_comb = smul32b_32b_x_32b(p0_TestBlock__A_op25, p0_TestBlock__B_op58);
  assign p1_smul_90069_comb = smul32b_32b_x_32b(p0_TestBlock__A_op26, p0_TestBlock__B_op68);
  assign p1_smul_90070_comb = smul32b_32b_x_32b(p0_TestBlock__A_op27, p0_TestBlock__B_op78);
  assign p1_smul_90071_comb = smul32b_32b_x_32b(p0_TestBlock__A_op28, p0_TestBlock__B_op88);
  assign p1_smul_90072_comb = smul32b_32b_x_32b(p0_TestBlock__A_op29, p0_TestBlock__B_op98);
  assign p1_smul_89615_comb = smul32b_32b_x_32b(p0_TestBlock__A_op20, p0_TestBlock__B_op9);
  assign p1_smul_89616_comb = smul32b_32b_x_32b(p0_TestBlock__A_op21, p0_TestBlock__B_op19);
  assign p1_smul_89617_comb = smul32b_32b_x_32b(p0_TestBlock__A_op22, p0_TestBlock__B_op29);
  assign p1_smul_89618_comb = smul32b_32b_x_32b(p0_TestBlock__A_op23, p0_TestBlock__B_op39);
  assign p1_smul_90073_comb = smul32b_32b_x_32b(p0_TestBlock__A_op24, p0_TestBlock__B_op49);
  assign p1_smul_90074_comb = smul32b_32b_x_32b(p0_TestBlock__A_op25, p0_TestBlock__B_op59);
  assign p1_smul_90075_comb = smul32b_32b_x_32b(p0_TestBlock__A_op26, p0_TestBlock__B_op69);
  assign p1_smul_90076_comb = smul32b_32b_x_32b(p0_TestBlock__A_op27, p0_TestBlock__B_op79);
  assign p1_smul_90077_comb = smul32b_32b_x_32b(p0_TestBlock__A_op28, p0_TestBlock__B_op89);
  assign p1_smul_90078_comb = smul32b_32b_x_32b(p0_TestBlock__A_op29, p0_TestBlock__B_op99);
  assign p1_smul_89619_comb = smul32b_32b_x_32b(p0_TestBlock__A_op30, p0_TestBlock__B_op0);
  assign p1_smul_89620_comb = smul32b_32b_x_32b(p0_TestBlock__A_op31, p0_TestBlock__B_op10);
  assign p1_smul_89621_comb = smul32b_32b_x_32b(p0_TestBlock__A_op32, p0_TestBlock__B_op20);
  assign p1_smul_89622_comb = smul32b_32b_x_32b(p0_TestBlock__A_op33, p0_TestBlock__B_op30);
  assign p1_smul_90079_comb = smul32b_32b_x_32b(p0_TestBlock__A_op34, p0_TestBlock__B_op40);
  assign p1_smul_90080_comb = smul32b_32b_x_32b(p0_TestBlock__A_op35, p0_TestBlock__B_op50);
  assign p1_smul_90081_comb = smul32b_32b_x_32b(p0_TestBlock__A_op36, p0_TestBlock__B_op60);
  assign p1_smul_90082_comb = smul32b_32b_x_32b(p0_TestBlock__A_op37, p0_TestBlock__B_op70);
  assign p1_smul_90083_comb = smul32b_32b_x_32b(p0_TestBlock__A_op38, p0_TestBlock__B_op80);
  assign p1_smul_90084_comb = smul32b_32b_x_32b(p0_TestBlock__A_op39, p0_TestBlock__B_op90);
  assign p1_smul_89623_comb = smul32b_32b_x_32b(p0_TestBlock__A_op30, p0_TestBlock__B_op1);
  assign p1_smul_89624_comb = smul32b_32b_x_32b(p0_TestBlock__A_op31, p0_TestBlock__B_op11);
  assign p1_smul_89625_comb = smul32b_32b_x_32b(p0_TestBlock__A_op32, p0_TestBlock__B_op21);
  assign p1_smul_89626_comb = smul32b_32b_x_32b(p0_TestBlock__A_op33, p0_TestBlock__B_op31);
  assign p1_smul_90085_comb = smul32b_32b_x_32b(p0_TestBlock__A_op34, p0_TestBlock__B_op41);
  assign p1_smul_90086_comb = smul32b_32b_x_32b(p0_TestBlock__A_op35, p0_TestBlock__B_op51);
  assign p1_smul_90087_comb = smul32b_32b_x_32b(p0_TestBlock__A_op36, p0_TestBlock__B_op61);
  assign p1_smul_90088_comb = smul32b_32b_x_32b(p0_TestBlock__A_op37, p0_TestBlock__B_op71);
  assign p1_smul_90089_comb = smul32b_32b_x_32b(p0_TestBlock__A_op38, p0_TestBlock__B_op81);
  assign p1_smul_90090_comb = smul32b_32b_x_32b(p0_TestBlock__A_op39, p0_TestBlock__B_op91);
  assign p1_smul_89627_comb = smul32b_32b_x_32b(p0_TestBlock__A_op30, p0_TestBlock__B_op2);
  assign p1_smul_89628_comb = smul32b_32b_x_32b(p0_TestBlock__A_op31, p0_TestBlock__B_op12);
  assign p1_smul_89629_comb = smul32b_32b_x_32b(p0_TestBlock__A_op32, p0_TestBlock__B_op22);
  assign p1_smul_89630_comb = smul32b_32b_x_32b(p0_TestBlock__A_op33, p0_TestBlock__B_op32);
  assign p1_smul_90091_comb = smul32b_32b_x_32b(p0_TestBlock__A_op34, p0_TestBlock__B_op42);
  assign p1_smul_90092_comb = smul32b_32b_x_32b(p0_TestBlock__A_op35, p0_TestBlock__B_op52);
  assign p1_smul_90093_comb = smul32b_32b_x_32b(p0_TestBlock__A_op36, p0_TestBlock__B_op62);
  assign p1_smul_90094_comb = smul32b_32b_x_32b(p0_TestBlock__A_op37, p0_TestBlock__B_op72);
  assign p1_smul_90095_comb = smul32b_32b_x_32b(p0_TestBlock__A_op38, p0_TestBlock__B_op82);
  assign p1_smul_90096_comb = smul32b_32b_x_32b(p0_TestBlock__A_op39, p0_TestBlock__B_op92);
  assign p1_smul_89631_comb = smul32b_32b_x_32b(p0_TestBlock__A_op30, p0_TestBlock__B_op3);
  assign p1_smul_89632_comb = smul32b_32b_x_32b(p0_TestBlock__A_op31, p0_TestBlock__B_op13);
  assign p1_smul_89633_comb = smul32b_32b_x_32b(p0_TestBlock__A_op32, p0_TestBlock__B_op23);
  assign p1_smul_89634_comb = smul32b_32b_x_32b(p0_TestBlock__A_op33, p0_TestBlock__B_op33);
  assign p1_smul_90097_comb = smul32b_32b_x_32b(p0_TestBlock__A_op34, p0_TestBlock__B_op43);
  assign p1_smul_90098_comb = smul32b_32b_x_32b(p0_TestBlock__A_op35, p0_TestBlock__B_op53);
  assign p1_smul_90099_comb = smul32b_32b_x_32b(p0_TestBlock__A_op36, p0_TestBlock__B_op63);
  assign p1_smul_90100_comb = smul32b_32b_x_32b(p0_TestBlock__A_op37, p0_TestBlock__B_op73);
  assign p1_smul_90101_comb = smul32b_32b_x_32b(p0_TestBlock__A_op38, p0_TestBlock__B_op83);
  assign p1_smul_90102_comb = smul32b_32b_x_32b(p0_TestBlock__A_op39, p0_TestBlock__B_op93);
  assign p1_smul_89635_comb = smul32b_32b_x_32b(p0_TestBlock__A_op30, p0_TestBlock__B_op4);
  assign p1_smul_89636_comb = smul32b_32b_x_32b(p0_TestBlock__A_op31, p0_TestBlock__B_op14);
  assign p1_smul_89637_comb = smul32b_32b_x_32b(p0_TestBlock__A_op32, p0_TestBlock__B_op24);
  assign p1_smul_89638_comb = smul32b_32b_x_32b(p0_TestBlock__A_op33, p0_TestBlock__B_op34);
  assign p1_smul_90103_comb = smul32b_32b_x_32b(p0_TestBlock__A_op34, p0_TestBlock__B_op44);
  assign p1_smul_90104_comb = smul32b_32b_x_32b(p0_TestBlock__A_op35, p0_TestBlock__B_op54);
  assign p1_smul_90105_comb = smul32b_32b_x_32b(p0_TestBlock__A_op36, p0_TestBlock__B_op64);
  assign p1_smul_90106_comb = smul32b_32b_x_32b(p0_TestBlock__A_op37, p0_TestBlock__B_op74);
  assign p1_smul_90107_comb = smul32b_32b_x_32b(p0_TestBlock__A_op38, p0_TestBlock__B_op84);
  assign p1_smul_90108_comb = smul32b_32b_x_32b(p0_TestBlock__A_op39, p0_TestBlock__B_op94);
  assign p1_smul_89639_comb = smul32b_32b_x_32b(p0_TestBlock__A_op30, p0_TestBlock__B_op5);
  assign p1_smul_89640_comb = smul32b_32b_x_32b(p0_TestBlock__A_op31, p0_TestBlock__B_op15);
  assign p1_smul_89641_comb = smul32b_32b_x_32b(p0_TestBlock__A_op32, p0_TestBlock__B_op25);
  assign p1_smul_89642_comb = smul32b_32b_x_32b(p0_TestBlock__A_op33, p0_TestBlock__B_op35);
  assign p1_smul_90109_comb = smul32b_32b_x_32b(p0_TestBlock__A_op34, p0_TestBlock__B_op45);
  assign p1_smul_90110_comb = smul32b_32b_x_32b(p0_TestBlock__A_op35, p0_TestBlock__B_op55);
  assign p1_smul_90111_comb = smul32b_32b_x_32b(p0_TestBlock__A_op36, p0_TestBlock__B_op65);
  assign p1_smul_90112_comb = smul32b_32b_x_32b(p0_TestBlock__A_op37, p0_TestBlock__B_op75);
  assign p1_smul_90113_comb = smul32b_32b_x_32b(p0_TestBlock__A_op38, p0_TestBlock__B_op85);
  assign p1_smul_90114_comb = smul32b_32b_x_32b(p0_TestBlock__A_op39, p0_TestBlock__B_op95);
  assign p1_smul_89643_comb = smul32b_32b_x_32b(p0_TestBlock__A_op30, p0_TestBlock__B_op6);
  assign p1_smul_89644_comb = smul32b_32b_x_32b(p0_TestBlock__A_op31, p0_TestBlock__B_op16);
  assign p1_smul_89645_comb = smul32b_32b_x_32b(p0_TestBlock__A_op32, p0_TestBlock__B_op26);
  assign p1_smul_89646_comb = smul32b_32b_x_32b(p0_TestBlock__A_op33, p0_TestBlock__B_op36);
  assign p1_smul_90115_comb = smul32b_32b_x_32b(p0_TestBlock__A_op34, p0_TestBlock__B_op46);
  assign p1_smul_90116_comb = smul32b_32b_x_32b(p0_TestBlock__A_op35, p0_TestBlock__B_op56);
  assign p1_smul_90117_comb = smul32b_32b_x_32b(p0_TestBlock__A_op36, p0_TestBlock__B_op66);
  assign p1_smul_90118_comb = smul32b_32b_x_32b(p0_TestBlock__A_op37, p0_TestBlock__B_op76);
  assign p1_smul_90119_comb = smul32b_32b_x_32b(p0_TestBlock__A_op38, p0_TestBlock__B_op86);
  assign p1_smul_90120_comb = smul32b_32b_x_32b(p0_TestBlock__A_op39, p0_TestBlock__B_op96);
  assign p1_smul_89647_comb = smul32b_32b_x_32b(p0_TestBlock__A_op30, p0_TestBlock__B_op7);
  assign p1_smul_89648_comb = smul32b_32b_x_32b(p0_TestBlock__A_op31, p0_TestBlock__B_op17);
  assign p1_smul_89649_comb = smul32b_32b_x_32b(p0_TestBlock__A_op32, p0_TestBlock__B_op27);
  assign p1_smul_89650_comb = smul32b_32b_x_32b(p0_TestBlock__A_op33, p0_TestBlock__B_op37);
  assign p1_smul_90121_comb = smul32b_32b_x_32b(p0_TestBlock__A_op34, p0_TestBlock__B_op47);
  assign p1_smul_90122_comb = smul32b_32b_x_32b(p0_TestBlock__A_op35, p0_TestBlock__B_op57);
  assign p1_smul_90123_comb = smul32b_32b_x_32b(p0_TestBlock__A_op36, p0_TestBlock__B_op67);
  assign p1_smul_90124_comb = smul32b_32b_x_32b(p0_TestBlock__A_op37, p0_TestBlock__B_op77);
  assign p1_smul_90125_comb = smul32b_32b_x_32b(p0_TestBlock__A_op38, p0_TestBlock__B_op87);
  assign p1_smul_90126_comb = smul32b_32b_x_32b(p0_TestBlock__A_op39, p0_TestBlock__B_op97);
  assign p1_smul_89651_comb = smul32b_32b_x_32b(p0_TestBlock__A_op30, p0_TestBlock__B_op8);
  assign p1_smul_89652_comb = smul32b_32b_x_32b(p0_TestBlock__A_op31, p0_TestBlock__B_op18);
  assign p1_smul_89653_comb = smul32b_32b_x_32b(p0_TestBlock__A_op32, p0_TestBlock__B_op28);
  assign p1_smul_89654_comb = smul32b_32b_x_32b(p0_TestBlock__A_op33, p0_TestBlock__B_op38);
  assign p1_smul_90127_comb = smul32b_32b_x_32b(p0_TestBlock__A_op34, p0_TestBlock__B_op48);
  assign p1_smul_90128_comb = smul32b_32b_x_32b(p0_TestBlock__A_op35, p0_TestBlock__B_op58);
  assign p1_smul_90129_comb = smul32b_32b_x_32b(p0_TestBlock__A_op36, p0_TestBlock__B_op68);
  assign p1_smul_90130_comb = smul32b_32b_x_32b(p0_TestBlock__A_op37, p0_TestBlock__B_op78);
  assign p1_smul_90131_comb = smul32b_32b_x_32b(p0_TestBlock__A_op38, p0_TestBlock__B_op88);
  assign p1_smul_90132_comb = smul32b_32b_x_32b(p0_TestBlock__A_op39, p0_TestBlock__B_op98);
  assign p1_smul_89655_comb = smul32b_32b_x_32b(p0_TestBlock__A_op30, p0_TestBlock__B_op9);
  assign p1_smul_89656_comb = smul32b_32b_x_32b(p0_TestBlock__A_op31, p0_TestBlock__B_op19);
  assign p1_smul_89657_comb = smul32b_32b_x_32b(p0_TestBlock__A_op32, p0_TestBlock__B_op29);
  assign p1_smul_89658_comb = smul32b_32b_x_32b(p0_TestBlock__A_op33, p0_TestBlock__B_op39);
  assign p1_smul_90133_comb = smul32b_32b_x_32b(p0_TestBlock__A_op34, p0_TestBlock__B_op49);
  assign p1_smul_90134_comb = smul32b_32b_x_32b(p0_TestBlock__A_op35, p0_TestBlock__B_op59);
  assign p1_smul_90135_comb = smul32b_32b_x_32b(p0_TestBlock__A_op36, p0_TestBlock__B_op69);
  assign p1_smul_90136_comb = smul32b_32b_x_32b(p0_TestBlock__A_op37, p0_TestBlock__B_op79);
  assign p1_smul_90137_comb = smul32b_32b_x_32b(p0_TestBlock__A_op38, p0_TestBlock__B_op89);
  assign p1_smul_90138_comb = smul32b_32b_x_32b(p0_TestBlock__A_op39, p0_TestBlock__B_op99);
  assign p1_smul_89659_comb = smul32b_32b_x_32b(p0_TestBlock__A_op40, p0_TestBlock__B_op0);
  assign p1_smul_89660_comb = smul32b_32b_x_32b(p0_TestBlock__A_op41, p0_TestBlock__B_op10);
  assign p1_smul_89661_comb = smul32b_32b_x_32b(p0_TestBlock__A_op42, p0_TestBlock__B_op20);
  assign p1_smul_89662_comb = smul32b_32b_x_32b(p0_TestBlock__A_op43, p0_TestBlock__B_op30);
  assign p1_smul_90139_comb = smul32b_32b_x_32b(p0_TestBlock__A_op44, p0_TestBlock__B_op40);
  assign p1_smul_90140_comb = smul32b_32b_x_32b(p0_TestBlock__A_op45, p0_TestBlock__B_op50);
  assign p1_smul_90141_comb = smul32b_32b_x_32b(p0_TestBlock__A_op46, p0_TestBlock__B_op60);
  assign p1_smul_90142_comb = smul32b_32b_x_32b(p0_TestBlock__A_op47, p0_TestBlock__B_op70);
  assign p1_smul_90143_comb = smul32b_32b_x_32b(p0_TestBlock__A_op48, p0_TestBlock__B_op80);
  assign p1_smul_90144_comb = smul32b_32b_x_32b(p0_TestBlock__A_op49, p0_TestBlock__B_op90);
  assign p1_smul_89663_comb = smul32b_32b_x_32b(p0_TestBlock__A_op40, p0_TestBlock__B_op1);
  assign p1_smul_89664_comb = smul32b_32b_x_32b(p0_TestBlock__A_op41, p0_TestBlock__B_op11);
  assign p1_smul_89665_comb = smul32b_32b_x_32b(p0_TestBlock__A_op42, p0_TestBlock__B_op21);
  assign p1_smul_89666_comb = smul32b_32b_x_32b(p0_TestBlock__A_op43, p0_TestBlock__B_op31);
  assign p1_smul_90145_comb = smul32b_32b_x_32b(p0_TestBlock__A_op44, p0_TestBlock__B_op41);
  assign p1_smul_90146_comb = smul32b_32b_x_32b(p0_TestBlock__A_op45, p0_TestBlock__B_op51);
  assign p1_smul_90147_comb = smul32b_32b_x_32b(p0_TestBlock__A_op46, p0_TestBlock__B_op61);
  assign p1_smul_90148_comb = smul32b_32b_x_32b(p0_TestBlock__A_op47, p0_TestBlock__B_op71);
  assign p1_smul_90149_comb = smul32b_32b_x_32b(p0_TestBlock__A_op48, p0_TestBlock__B_op81);
  assign p1_smul_90150_comb = smul32b_32b_x_32b(p0_TestBlock__A_op49, p0_TestBlock__B_op91);
  assign p1_smul_89667_comb = smul32b_32b_x_32b(p0_TestBlock__A_op40, p0_TestBlock__B_op2);
  assign p1_smul_89668_comb = smul32b_32b_x_32b(p0_TestBlock__A_op41, p0_TestBlock__B_op12);
  assign p1_smul_89669_comb = smul32b_32b_x_32b(p0_TestBlock__A_op42, p0_TestBlock__B_op22);
  assign p1_smul_89670_comb = smul32b_32b_x_32b(p0_TestBlock__A_op43, p0_TestBlock__B_op32);
  assign p1_smul_90151_comb = smul32b_32b_x_32b(p0_TestBlock__A_op44, p0_TestBlock__B_op42);
  assign p1_smul_90152_comb = smul32b_32b_x_32b(p0_TestBlock__A_op45, p0_TestBlock__B_op52);
  assign p1_smul_90153_comb = smul32b_32b_x_32b(p0_TestBlock__A_op46, p0_TestBlock__B_op62);
  assign p1_smul_90154_comb = smul32b_32b_x_32b(p0_TestBlock__A_op47, p0_TestBlock__B_op72);
  assign p1_smul_90155_comb = smul32b_32b_x_32b(p0_TestBlock__A_op48, p0_TestBlock__B_op82);
  assign p1_smul_90156_comb = smul32b_32b_x_32b(p0_TestBlock__A_op49, p0_TestBlock__B_op92);
  assign p1_smul_89671_comb = smul32b_32b_x_32b(p0_TestBlock__A_op40, p0_TestBlock__B_op3);
  assign p1_smul_89672_comb = smul32b_32b_x_32b(p0_TestBlock__A_op41, p0_TestBlock__B_op13);
  assign p1_smul_89673_comb = smul32b_32b_x_32b(p0_TestBlock__A_op42, p0_TestBlock__B_op23);
  assign p1_smul_89674_comb = smul32b_32b_x_32b(p0_TestBlock__A_op43, p0_TestBlock__B_op33);
  assign p1_smul_90157_comb = smul32b_32b_x_32b(p0_TestBlock__A_op44, p0_TestBlock__B_op43);
  assign p1_smul_90158_comb = smul32b_32b_x_32b(p0_TestBlock__A_op45, p0_TestBlock__B_op53);
  assign p1_smul_90159_comb = smul32b_32b_x_32b(p0_TestBlock__A_op46, p0_TestBlock__B_op63);
  assign p1_smul_90160_comb = smul32b_32b_x_32b(p0_TestBlock__A_op47, p0_TestBlock__B_op73);
  assign p1_smul_90161_comb = smul32b_32b_x_32b(p0_TestBlock__A_op48, p0_TestBlock__B_op83);
  assign p1_smul_90162_comb = smul32b_32b_x_32b(p0_TestBlock__A_op49, p0_TestBlock__B_op93);
  assign p1_smul_89675_comb = smul32b_32b_x_32b(p0_TestBlock__A_op40, p0_TestBlock__B_op4);
  assign p1_smul_89676_comb = smul32b_32b_x_32b(p0_TestBlock__A_op41, p0_TestBlock__B_op14);
  assign p1_smul_89677_comb = smul32b_32b_x_32b(p0_TestBlock__A_op42, p0_TestBlock__B_op24);
  assign p1_smul_89678_comb = smul32b_32b_x_32b(p0_TestBlock__A_op43, p0_TestBlock__B_op34);
  assign p1_smul_90163_comb = smul32b_32b_x_32b(p0_TestBlock__A_op44, p0_TestBlock__B_op44);
  assign p1_smul_90164_comb = smul32b_32b_x_32b(p0_TestBlock__A_op45, p0_TestBlock__B_op54);
  assign p1_smul_90165_comb = smul32b_32b_x_32b(p0_TestBlock__A_op46, p0_TestBlock__B_op64);
  assign p1_smul_90166_comb = smul32b_32b_x_32b(p0_TestBlock__A_op47, p0_TestBlock__B_op74);
  assign p1_smul_90167_comb = smul32b_32b_x_32b(p0_TestBlock__A_op48, p0_TestBlock__B_op84);
  assign p1_smul_90168_comb = smul32b_32b_x_32b(p0_TestBlock__A_op49, p0_TestBlock__B_op94);
  assign p1_smul_89679_comb = smul32b_32b_x_32b(p0_TestBlock__A_op40, p0_TestBlock__B_op5);
  assign p1_smul_89680_comb = smul32b_32b_x_32b(p0_TestBlock__A_op41, p0_TestBlock__B_op15);
  assign p1_smul_89681_comb = smul32b_32b_x_32b(p0_TestBlock__A_op42, p0_TestBlock__B_op25);
  assign p1_smul_89682_comb = smul32b_32b_x_32b(p0_TestBlock__A_op43, p0_TestBlock__B_op35);
  assign p1_smul_90169_comb = smul32b_32b_x_32b(p0_TestBlock__A_op44, p0_TestBlock__B_op45);
  assign p1_smul_90170_comb = smul32b_32b_x_32b(p0_TestBlock__A_op45, p0_TestBlock__B_op55);
  assign p1_smul_90171_comb = smul32b_32b_x_32b(p0_TestBlock__A_op46, p0_TestBlock__B_op65);
  assign p1_smul_90172_comb = smul32b_32b_x_32b(p0_TestBlock__A_op47, p0_TestBlock__B_op75);
  assign p1_smul_90173_comb = smul32b_32b_x_32b(p0_TestBlock__A_op48, p0_TestBlock__B_op85);
  assign p1_smul_90174_comb = smul32b_32b_x_32b(p0_TestBlock__A_op49, p0_TestBlock__B_op95);
  assign p1_smul_89683_comb = smul32b_32b_x_32b(p0_TestBlock__A_op40, p0_TestBlock__B_op6);
  assign p1_smul_89684_comb = smul32b_32b_x_32b(p0_TestBlock__A_op41, p0_TestBlock__B_op16);
  assign p1_smul_89685_comb = smul32b_32b_x_32b(p0_TestBlock__A_op42, p0_TestBlock__B_op26);
  assign p1_smul_89686_comb = smul32b_32b_x_32b(p0_TestBlock__A_op43, p0_TestBlock__B_op36);
  assign p1_smul_90175_comb = smul32b_32b_x_32b(p0_TestBlock__A_op44, p0_TestBlock__B_op46);
  assign p1_smul_90176_comb = smul32b_32b_x_32b(p0_TestBlock__A_op45, p0_TestBlock__B_op56);
  assign p1_smul_90177_comb = smul32b_32b_x_32b(p0_TestBlock__A_op46, p0_TestBlock__B_op66);
  assign p1_smul_90178_comb = smul32b_32b_x_32b(p0_TestBlock__A_op47, p0_TestBlock__B_op76);
  assign p1_smul_90179_comb = smul32b_32b_x_32b(p0_TestBlock__A_op48, p0_TestBlock__B_op86);
  assign p1_smul_90180_comb = smul32b_32b_x_32b(p0_TestBlock__A_op49, p0_TestBlock__B_op96);
  assign p1_smul_89687_comb = smul32b_32b_x_32b(p0_TestBlock__A_op40, p0_TestBlock__B_op7);
  assign p1_smul_89688_comb = smul32b_32b_x_32b(p0_TestBlock__A_op41, p0_TestBlock__B_op17);
  assign p1_smul_89689_comb = smul32b_32b_x_32b(p0_TestBlock__A_op42, p0_TestBlock__B_op27);
  assign p1_smul_89690_comb = smul32b_32b_x_32b(p0_TestBlock__A_op43, p0_TestBlock__B_op37);
  assign p1_smul_90181_comb = smul32b_32b_x_32b(p0_TestBlock__A_op44, p0_TestBlock__B_op47);
  assign p1_smul_90182_comb = smul32b_32b_x_32b(p0_TestBlock__A_op45, p0_TestBlock__B_op57);
  assign p1_smul_90183_comb = smul32b_32b_x_32b(p0_TestBlock__A_op46, p0_TestBlock__B_op67);
  assign p1_smul_90184_comb = smul32b_32b_x_32b(p0_TestBlock__A_op47, p0_TestBlock__B_op77);
  assign p1_smul_90185_comb = smul32b_32b_x_32b(p0_TestBlock__A_op48, p0_TestBlock__B_op87);
  assign p1_smul_90186_comb = smul32b_32b_x_32b(p0_TestBlock__A_op49, p0_TestBlock__B_op97);
  assign p1_smul_89691_comb = smul32b_32b_x_32b(p0_TestBlock__A_op40, p0_TestBlock__B_op8);
  assign p1_smul_89692_comb = smul32b_32b_x_32b(p0_TestBlock__A_op41, p0_TestBlock__B_op18);
  assign p1_smul_89693_comb = smul32b_32b_x_32b(p0_TestBlock__A_op42, p0_TestBlock__B_op28);
  assign p1_smul_89694_comb = smul32b_32b_x_32b(p0_TestBlock__A_op43, p0_TestBlock__B_op38);
  assign p1_smul_90187_comb = smul32b_32b_x_32b(p0_TestBlock__A_op44, p0_TestBlock__B_op48);
  assign p1_smul_90188_comb = smul32b_32b_x_32b(p0_TestBlock__A_op45, p0_TestBlock__B_op58);
  assign p1_smul_90189_comb = smul32b_32b_x_32b(p0_TestBlock__A_op46, p0_TestBlock__B_op68);
  assign p1_smul_90190_comb = smul32b_32b_x_32b(p0_TestBlock__A_op47, p0_TestBlock__B_op78);
  assign p1_smul_90191_comb = smul32b_32b_x_32b(p0_TestBlock__A_op48, p0_TestBlock__B_op88);
  assign p1_smul_90192_comb = smul32b_32b_x_32b(p0_TestBlock__A_op49, p0_TestBlock__B_op98);
  assign p1_smul_89695_comb = smul32b_32b_x_32b(p0_TestBlock__A_op40, p0_TestBlock__B_op9);
  assign p1_smul_89696_comb = smul32b_32b_x_32b(p0_TestBlock__A_op41, p0_TestBlock__B_op19);
  assign p1_smul_89697_comb = smul32b_32b_x_32b(p0_TestBlock__A_op42, p0_TestBlock__B_op29);
  assign p1_smul_89698_comb = smul32b_32b_x_32b(p0_TestBlock__A_op43, p0_TestBlock__B_op39);
  assign p1_smul_90193_comb = smul32b_32b_x_32b(p0_TestBlock__A_op44, p0_TestBlock__B_op49);
  assign p1_smul_90194_comb = smul32b_32b_x_32b(p0_TestBlock__A_op45, p0_TestBlock__B_op59);
  assign p1_smul_90195_comb = smul32b_32b_x_32b(p0_TestBlock__A_op46, p0_TestBlock__B_op69);
  assign p1_smul_90196_comb = smul32b_32b_x_32b(p0_TestBlock__A_op47, p0_TestBlock__B_op79);
  assign p1_smul_90197_comb = smul32b_32b_x_32b(p0_TestBlock__A_op48, p0_TestBlock__B_op89);
  assign p1_smul_90198_comb = smul32b_32b_x_32b(p0_TestBlock__A_op49, p0_TestBlock__B_op99);
  assign p1_smul_89699_comb = smul32b_32b_x_32b(p0_TestBlock__A_op50, p0_TestBlock__B_op0);
  assign p1_smul_89700_comb = smul32b_32b_x_32b(p0_TestBlock__A_op51, p0_TestBlock__B_op10);
  assign p1_smul_89701_comb = smul32b_32b_x_32b(p0_TestBlock__A_op52, p0_TestBlock__B_op20);
  assign p1_smul_89702_comb = smul32b_32b_x_32b(p0_TestBlock__A_op53, p0_TestBlock__B_op30);
  assign p1_smul_90199_comb = smul32b_32b_x_32b(p0_TestBlock__A_op54, p0_TestBlock__B_op40);
  assign p1_smul_90200_comb = smul32b_32b_x_32b(p0_TestBlock__A_op55, p0_TestBlock__B_op50);
  assign p1_smul_90201_comb = smul32b_32b_x_32b(p0_TestBlock__A_op56, p0_TestBlock__B_op60);
  assign p1_smul_90202_comb = smul32b_32b_x_32b(p0_TestBlock__A_op57, p0_TestBlock__B_op70);
  assign p1_smul_90203_comb = smul32b_32b_x_32b(p0_TestBlock__A_op58, p0_TestBlock__B_op80);
  assign p1_smul_90204_comb = smul32b_32b_x_32b(p0_TestBlock__A_op59, p0_TestBlock__B_op90);
  assign p1_smul_89703_comb = smul32b_32b_x_32b(p0_TestBlock__A_op50, p0_TestBlock__B_op1);
  assign p1_smul_89704_comb = smul32b_32b_x_32b(p0_TestBlock__A_op51, p0_TestBlock__B_op11);
  assign p1_smul_89705_comb = smul32b_32b_x_32b(p0_TestBlock__A_op52, p0_TestBlock__B_op21);
  assign p1_smul_89706_comb = smul32b_32b_x_32b(p0_TestBlock__A_op53, p0_TestBlock__B_op31);
  assign p1_smul_90205_comb = smul32b_32b_x_32b(p0_TestBlock__A_op54, p0_TestBlock__B_op41);
  assign p1_smul_90206_comb = smul32b_32b_x_32b(p0_TestBlock__A_op55, p0_TestBlock__B_op51);
  assign p1_smul_90207_comb = smul32b_32b_x_32b(p0_TestBlock__A_op56, p0_TestBlock__B_op61);
  assign p1_smul_90208_comb = smul32b_32b_x_32b(p0_TestBlock__A_op57, p0_TestBlock__B_op71);
  assign p1_smul_90209_comb = smul32b_32b_x_32b(p0_TestBlock__A_op58, p0_TestBlock__B_op81);
  assign p1_smul_90210_comb = smul32b_32b_x_32b(p0_TestBlock__A_op59, p0_TestBlock__B_op91);
  assign p1_smul_89707_comb = smul32b_32b_x_32b(p0_TestBlock__A_op50, p0_TestBlock__B_op2);
  assign p1_smul_89708_comb = smul32b_32b_x_32b(p0_TestBlock__A_op51, p0_TestBlock__B_op12);
  assign p1_smul_89709_comb = smul32b_32b_x_32b(p0_TestBlock__A_op52, p0_TestBlock__B_op22);
  assign p1_smul_89710_comb = smul32b_32b_x_32b(p0_TestBlock__A_op53, p0_TestBlock__B_op32);
  assign p1_smul_90211_comb = smul32b_32b_x_32b(p0_TestBlock__A_op54, p0_TestBlock__B_op42);
  assign p1_smul_90212_comb = smul32b_32b_x_32b(p0_TestBlock__A_op55, p0_TestBlock__B_op52);
  assign p1_smul_90213_comb = smul32b_32b_x_32b(p0_TestBlock__A_op56, p0_TestBlock__B_op62);
  assign p1_smul_90214_comb = smul32b_32b_x_32b(p0_TestBlock__A_op57, p0_TestBlock__B_op72);
  assign p1_smul_90215_comb = smul32b_32b_x_32b(p0_TestBlock__A_op58, p0_TestBlock__B_op82);
  assign p1_smul_90216_comb = smul32b_32b_x_32b(p0_TestBlock__A_op59, p0_TestBlock__B_op92);
  assign p1_smul_89711_comb = smul32b_32b_x_32b(p0_TestBlock__A_op50, p0_TestBlock__B_op3);
  assign p1_smul_89712_comb = smul32b_32b_x_32b(p0_TestBlock__A_op51, p0_TestBlock__B_op13);
  assign p1_smul_89713_comb = smul32b_32b_x_32b(p0_TestBlock__A_op52, p0_TestBlock__B_op23);
  assign p1_smul_89714_comb = smul32b_32b_x_32b(p0_TestBlock__A_op53, p0_TestBlock__B_op33);
  assign p1_smul_90217_comb = smul32b_32b_x_32b(p0_TestBlock__A_op54, p0_TestBlock__B_op43);
  assign p1_smul_90218_comb = smul32b_32b_x_32b(p0_TestBlock__A_op55, p0_TestBlock__B_op53);
  assign p1_smul_90219_comb = smul32b_32b_x_32b(p0_TestBlock__A_op56, p0_TestBlock__B_op63);
  assign p1_smul_90220_comb = smul32b_32b_x_32b(p0_TestBlock__A_op57, p0_TestBlock__B_op73);
  assign p1_smul_90221_comb = smul32b_32b_x_32b(p0_TestBlock__A_op58, p0_TestBlock__B_op83);
  assign p1_smul_90222_comb = smul32b_32b_x_32b(p0_TestBlock__A_op59, p0_TestBlock__B_op93);
  assign p1_smul_89715_comb = smul32b_32b_x_32b(p0_TestBlock__A_op50, p0_TestBlock__B_op4);
  assign p1_smul_89716_comb = smul32b_32b_x_32b(p0_TestBlock__A_op51, p0_TestBlock__B_op14);
  assign p1_smul_89717_comb = smul32b_32b_x_32b(p0_TestBlock__A_op52, p0_TestBlock__B_op24);
  assign p1_smul_89718_comb = smul32b_32b_x_32b(p0_TestBlock__A_op53, p0_TestBlock__B_op34);
  assign p1_smul_90223_comb = smul32b_32b_x_32b(p0_TestBlock__A_op54, p0_TestBlock__B_op44);
  assign p1_smul_90224_comb = smul32b_32b_x_32b(p0_TestBlock__A_op55, p0_TestBlock__B_op54);
  assign p1_smul_90225_comb = smul32b_32b_x_32b(p0_TestBlock__A_op56, p0_TestBlock__B_op64);
  assign p1_smul_90226_comb = smul32b_32b_x_32b(p0_TestBlock__A_op57, p0_TestBlock__B_op74);
  assign p1_smul_90227_comb = smul32b_32b_x_32b(p0_TestBlock__A_op58, p0_TestBlock__B_op84);
  assign p1_smul_90228_comb = smul32b_32b_x_32b(p0_TestBlock__A_op59, p0_TestBlock__B_op94);
  assign p1_smul_89719_comb = smul32b_32b_x_32b(p0_TestBlock__A_op50, p0_TestBlock__B_op5);
  assign p1_smul_89720_comb = smul32b_32b_x_32b(p0_TestBlock__A_op51, p0_TestBlock__B_op15);
  assign p1_smul_89721_comb = smul32b_32b_x_32b(p0_TestBlock__A_op52, p0_TestBlock__B_op25);
  assign p1_smul_89722_comb = smul32b_32b_x_32b(p0_TestBlock__A_op53, p0_TestBlock__B_op35);
  assign p1_smul_90229_comb = smul32b_32b_x_32b(p0_TestBlock__A_op54, p0_TestBlock__B_op45);
  assign p1_smul_90230_comb = smul32b_32b_x_32b(p0_TestBlock__A_op55, p0_TestBlock__B_op55);
  assign p1_smul_90231_comb = smul32b_32b_x_32b(p0_TestBlock__A_op56, p0_TestBlock__B_op65);
  assign p1_smul_90232_comb = smul32b_32b_x_32b(p0_TestBlock__A_op57, p0_TestBlock__B_op75);
  assign p1_smul_90233_comb = smul32b_32b_x_32b(p0_TestBlock__A_op58, p0_TestBlock__B_op85);
  assign p1_smul_90234_comb = smul32b_32b_x_32b(p0_TestBlock__A_op59, p0_TestBlock__B_op95);
  assign p1_smul_89723_comb = smul32b_32b_x_32b(p0_TestBlock__A_op50, p0_TestBlock__B_op6);
  assign p1_smul_89724_comb = smul32b_32b_x_32b(p0_TestBlock__A_op51, p0_TestBlock__B_op16);
  assign p1_smul_89725_comb = smul32b_32b_x_32b(p0_TestBlock__A_op52, p0_TestBlock__B_op26);
  assign p1_smul_89726_comb = smul32b_32b_x_32b(p0_TestBlock__A_op53, p0_TestBlock__B_op36);
  assign p1_smul_90235_comb = smul32b_32b_x_32b(p0_TestBlock__A_op54, p0_TestBlock__B_op46);
  assign p1_smul_90236_comb = smul32b_32b_x_32b(p0_TestBlock__A_op55, p0_TestBlock__B_op56);
  assign p1_smul_90237_comb = smul32b_32b_x_32b(p0_TestBlock__A_op56, p0_TestBlock__B_op66);
  assign p1_smul_90238_comb = smul32b_32b_x_32b(p0_TestBlock__A_op57, p0_TestBlock__B_op76);
  assign p1_smul_90239_comb = smul32b_32b_x_32b(p0_TestBlock__A_op58, p0_TestBlock__B_op86);
  assign p1_smul_90240_comb = smul32b_32b_x_32b(p0_TestBlock__A_op59, p0_TestBlock__B_op96);
  assign p1_smul_89727_comb = smul32b_32b_x_32b(p0_TestBlock__A_op50, p0_TestBlock__B_op7);
  assign p1_smul_89728_comb = smul32b_32b_x_32b(p0_TestBlock__A_op51, p0_TestBlock__B_op17);
  assign p1_smul_89729_comb = smul32b_32b_x_32b(p0_TestBlock__A_op52, p0_TestBlock__B_op27);
  assign p1_smul_89730_comb = smul32b_32b_x_32b(p0_TestBlock__A_op53, p0_TestBlock__B_op37);
  assign p1_smul_90241_comb = smul32b_32b_x_32b(p0_TestBlock__A_op54, p0_TestBlock__B_op47);
  assign p1_smul_90242_comb = smul32b_32b_x_32b(p0_TestBlock__A_op55, p0_TestBlock__B_op57);
  assign p1_smul_90243_comb = smul32b_32b_x_32b(p0_TestBlock__A_op56, p0_TestBlock__B_op67);
  assign p1_smul_90244_comb = smul32b_32b_x_32b(p0_TestBlock__A_op57, p0_TestBlock__B_op77);
  assign p1_smul_90245_comb = smul32b_32b_x_32b(p0_TestBlock__A_op58, p0_TestBlock__B_op87);
  assign p1_smul_90246_comb = smul32b_32b_x_32b(p0_TestBlock__A_op59, p0_TestBlock__B_op97);
  assign p1_smul_89731_comb = smul32b_32b_x_32b(p0_TestBlock__A_op50, p0_TestBlock__B_op8);
  assign p1_smul_89732_comb = smul32b_32b_x_32b(p0_TestBlock__A_op51, p0_TestBlock__B_op18);
  assign p1_smul_89733_comb = smul32b_32b_x_32b(p0_TestBlock__A_op52, p0_TestBlock__B_op28);
  assign p1_smul_89734_comb = smul32b_32b_x_32b(p0_TestBlock__A_op53, p0_TestBlock__B_op38);
  assign p1_smul_90247_comb = smul32b_32b_x_32b(p0_TestBlock__A_op54, p0_TestBlock__B_op48);
  assign p1_smul_90248_comb = smul32b_32b_x_32b(p0_TestBlock__A_op55, p0_TestBlock__B_op58);
  assign p1_smul_90249_comb = smul32b_32b_x_32b(p0_TestBlock__A_op56, p0_TestBlock__B_op68);
  assign p1_smul_90250_comb = smul32b_32b_x_32b(p0_TestBlock__A_op57, p0_TestBlock__B_op78);
  assign p1_smul_90251_comb = smul32b_32b_x_32b(p0_TestBlock__A_op58, p0_TestBlock__B_op88);
  assign p1_smul_90252_comb = smul32b_32b_x_32b(p0_TestBlock__A_op59, p0_TestBlock__B_op98);
  assign p1_smul_89735_comb = smul32b_32b_x_32b(p0_TestBlock__A_op50, p0_TestBlock__B_op9);
  assign p1_smul_89736_comb = smul32b_32b_x_32b(p0_TestBlock__A_op51, p0_TestBlock__B_op19);
  assign p1_smul_89737_comb = smul32b_32b_x_32b(p0_TestBlock__A_op52, p0_TestBlock__B_op29);
  assign p1_smul_89738_comb = smul32b_32b_x_32b(p0_TestBlock__A_op53, p0_TestBlock__B_op39);
  assign p1_smul_90253_comb = smul32b_32b_x_32b(p0_TestBlock__A_op54, p0_TestBlock__B_op49);
  assign p1_smul_90254_comb = smul32b_32b_x_32b(p0_TestBlock__A_op55, p0_TestBlock__B_op59);
  assign p1_smul_90255_comb = smul32b_32b_x_32b(p0_TestBlock__A_op56, p0_TestBlock__B_op69);
  assign p1_smul_90256_comb = smul32b_32b_x_32b(p0_TestBlock__A_op57, p0_TestBlock__B_op79);
  assign p1_smul_90257_comb = smul32b_32b_x_32b(p0_TestBlock__A_op58, p0_TestBlock__B_op89);
  assign p1_smul_90258_comb = smul32b_32b_x_32b(p0_TestBlock__A_op59, p0_TestBlock__B_op99);
  assign p1_smul_89739_comb = smul32b_32b_x_32b(p0_TestBlock__A_op60, p0_TestBlock__B_op0);
  assign p1_smul_89740_comb = smul32b_32b_x_32b(p0_TestBlock__A_op61, p0_TestBlock__B_op10);
  assign p1_smul_89741_comb = smul32b_32b_x_32b(p0_TestBlock__A_op62, p0_TestBlock__B_op20);
  assign p1_smul_89742_comb = smul32b_32b_x_32b(p0_TestBlock__A_op63, p0_TestBlock__B_op30);
  assign p1_smul_90259_comb = smul32b_32b_x_32b(p0_TestBlock__A_op64, p0_TestBlock__B_op40);
  assign p1_smul_90260_comb = smul32b_32b_x_32b(p0_TestBlock__A_op65, p0_TestBlock__B_op50);
  assign p1_smul_90261_comb = smul32b_32b_x_32b(p0_TestBlock__A_op66, p0_TestBlock__B_op60);
  assign p1_smul_90262_comb = smul32b_32b_x_32b(p0_TestBlock__A_op67, p0_TestBlock__B_op70);
  assign p1_smul_90263_comb = smul32b_32b_x_32b(p0_TestBlock__A_op68, p0_TestBlock__B_op80);
  assign p1_smul_90264_comb = smul32b_32b_x_32b(p0_TestBlock__A_op69, p0_TestBlock__B_op90);
  assign p1_smul_89743_comb = smul32b_32b_x_32b(p0_TestBlock__A_op60, p0_TestBlock__B_op1);
  assign p1_smul_89744_comb = smul32b_32b_x_32b(p0_TestBlock__A_op61, p0_TestBlock__B_op11);
  assign p1_smul_89745_comb = smul32b_32b_x_32b(p0_TestBlock__A_op62, p0_TestBlock__B_op21);
  assign p1_smul_89746_comb = smul32b_32b_x_32b(p0_TestBlock__A_op63, p0_TestBlock__B_op31);
  assign p1_smul_90265_comb = smul32b_32b_x_32b(p0_TestBlock__A_op64, p0_TestBlock__B_op41);
  assign p1_smul_90266_comb = smul32b_32b_x_32b(p0_TestBlock__A_op65, p0_TestBlock__B_op51);
  assign p1_smul_90267_comb = smul32b_32b_x_32b(p0_TestBlock__A_op66, p0_TestBlock__B_op61);
  assign p1_smul_90268_comb = smul32b_32b_x_32b(p0_TestBlock__A_op67, p0_TestBlock__B_op71);
  assign p1_smul_90269_comb = smul32b_32b_x_32b(p0_TestBlock__A_op68, p0_TestBlock__B_op81);
  assign p1_smul_90270_comb = smul32b_32b_x_32b(p0_TestBlock__A_op69, p0_TestBlock__B_op91);
  assign p1_smul_89747_comb = smul32b_32b_x_32b(p0_TestBlock__A_op60, p0_TestBlock__B_op2);
  assign p1_smul_89748_comb = smul32b_32b_x_32b(p0_TestBlock__A_op61, p0_TestBlock__B_op12);
  assign p1_smul_89749_comb = smul32b_32b_x_32b(p0_TestBlock__A_op62, p0_TestBlock__B_op22);
  assign p1_smul_89750_comb = smul32b_32b_x_32b(p0_TestBlock__A_op63, p0_TestBlock__B_op32);
  assign p1_smul_90271_comb = smul32b_32b_x_32b(p0_TestBlock__A_op64, p0_TestBlock__B_op42);
  assign p1_smul_90272_comb = smul32b_32b_x_32b(p0_TestBlock__A_op65, p0_TestBlock__B_op52);
  assign p1_smul_90273_comb = smul32b_32b_x_32b(p0_TestBlock__A_op66, p0_TestBlock__B_op62);
  assign p1_smul_90274_comb = smul32b_32b_x_32b(p0_TestBlock__A_op67, p0_TestBlock__B_op72);
  assign p1_smul_90275_comb = smul32b_32b_x_32b(p0_TestBlock__A_op68, p0_TestBlock__B_op82);
  assign p1_smul_90276_comb = smul32b_32b_x_32b(p0_TestBlock__A_op69, p0_TestBlock__B_op92);
  assign p1_smul_89751_comb = smul32b_32b_x_32b(p0_TestBlock__A_op60, p0_TestBlock__B_op3);
  assign p1_smul_89752_comb = smul32b_32b_x_32b(p0_TestBlock__A_op61, p0_TestBlock__B_op13);
  assign p1_smul_89753_comb = smul32b_32b_x_32b(p0_TestBlock__A_op62, p0_TestBlock__B_op23);
  assign p1_smul_89754_comb = smul32b_32b_x_32b(p0_TestBlock__A_op63, p0_TestBlock__B_op33);
  assign p1_smul_90277_comb = smul32b_32b_x_32b(p0_TestBlock__A_op64, p0_TestBlock__B_op43);
  assign p1_smul_90278_comb = smul32b_32b_x_32b(p0_TestBlock__A_op65, p0_TestBlock__B_op53);
  assign p1_smul_90279_comb = smul32b_32b_x_32b(p0_TestBlock__A_op66, p0_TestBlock__B_op63);
  assign p1_smul_90280_comb = smul32b_32b_x_32b(p0_TestBlock__A_op67, p0_TestBlock__B_op73);
  assign p1_smul_90281_comb = smul32b_32b_x_32b(p0_TestBlock__A_op68, p0_TestBlock__B_op83);
  assign p1_smul_90282_comb = smul32b_32b_x_32b(p0_TestBlock__A_op69, p0_TestBlock__B_op93);
  assign p1_smul_89755_comb = smul32b_32b_x_32b(p0_TestBlock__A_op60, p0_TestBlock__B_op4);
  assign p1_smul_89756_comb = smul32b_32b_x_32b(p0_TestBlock__A_op61, p0_TestBlock__B_op14);
  assign p1_smul_89757_comb = smul32b_32b_x_32b(p0_TestBlock__A_op62, p0_TestBlock__B_op24);
  assign p1_smul_89758_comb = smul32b_32b_x_32b(p0_TestBlock__A_op63, p0_TestBlock__B_op34);
  assign p1_smul_90283_comb = smul32b_32b_x_32b(p0_TestBlock__A_op64, p0_TestBlock__B_op44);
  assign p1_smul_90284_comb = smul32b_32b_x_32b(p0_TestBlock__A_op65, p0_TestBlock__B_op54);
  assign p1_smul_90285_comb = smul32b_32b_x_32b(p0_TestBlock__A_op66, p0_TestBlock__B_op64);
  assign p1_smul_90286_comb = smul32b_32b_x_32b(p0_TestBlock__A_op67, p0_TestBlock__B_op74);
  assign p1_smul_90287_comb = smul32b_32b_x_32b(p0_TestBlock__A_op68, p0_TestBlock__B_op84);
  assign p1_smul_90288_comb = smul32b_32b_x_32b(p0_TestBlock__A_op69, p0_TestBlock__B_op94);
  assign p1_smul_89759_comb = smul32b_32b_x_32b(p0_TestBlock__A_op60, p0_TestBlock__B_op5);
  assign p1_smul_89760_comb = smul32b_32b_x_32b(p0_TestBlock__A_op61, p0_TestBlock__B_op15);
  assign p1_smul_89761_comb = smul32b_32b_x_32b(p0_TestBlock__A_op62, p0_TestBlock__B_op25);
  assign p1_smul_89762_comb = smul32b_32b_x_32b(p0_TestBlock__A_op63, p0_TestBlock__B_op35);
  assign p1_smul_90289_comb = smul32b_32b_x_32b(p0_TestBlock__A_op64, p0_TestBlock__B_op45);
  assign p1_smul_90290_comb = smul32b_32b_x_32b(p0_TestBlock__A_op65, p0_TestBlock__B_op55);
  assign p1_smul_90291_comb = smul32b_32b_x_32b(p0_TestBlock__A_op66, p0_TestBlock__B_op65);
  assign p1_smul_90292_comb = smul32b_32b_x_32b(p0_TestBlock__A_op67, p0_TestBlock__B_op75);
  assign p1_smul_90293_comb = smul32b_32b_x_32b(p0_TestBlock__A_op68, p0_TestBlock__B_op85);
  assign p1_smul_90294_comb = smul32b_32b_x_32b(p0_TestBlock__A_op69, p0_TestBlock__B_op95);
  assign p1_smul_89763_comb = smul32b_32b_x_32b(p0_TestBlock__A_op60, p0_TestBlock__B_op6);
  assign p1_smul_89764_comb = smul32b_32b_x_32b(p0_TestBlock__A_op61, p0_TestBlock__B_op16);
  assign p1_smul_89765_comb = smul32b_32b_x_32b(p0_TestBlock__A_op62, p0_TestBlock__B_op26);
  assign p1_smul_89766_comb = smul32b_32b_x_32b(p0_TestBlock__A_op63, p0_TestBlock__B_op36);
  assign p1_smul_90295_comb = smul32b_32b_x_32b(p0_TestBlock__A_op64, p0_TestBlock__B_op46);
  assign p1_smul_90296_comb = smul32b_32b_x_32b(p0_TestBlock__A_op65, p0_TestBlock__B_op56);
  assign p1_smul_90297_comb = smul32b_32b_x_32b(p0_TestBlock__A_op66, p0_TestBlock__B_op66);
  assign p1_smul_90298_comb = smul32b_32b_x_32b(p0_TestBlock__A_op67, p0_TestBlock__B_op76);
  assign p1_smul_90299_comb = smul32b_32b_x_32b(p0_TestBlock__A_op68, p0_TestBlock__B_op86);
  assign p1_smul_90300_comb = smul32b_32b_x_32b(p0_TestBlock__A_op69, p0_TestBlock__B_op96);
  assign p1_smul_89767_comb = smul32b_32b_x_32b(p0_TestBlock__A_op60, p0_TestBlock__B_op7);
  assign p1_smul_89768_comb = smul32b_32b_x_32b(p0_TestBlock__A_op61, p0_TestBlock__B_op17);
  assign p1_smul_89769_comb = smul32b_32b_x_32b(p0_TestBlock__A_op62, p0_TestBlock__B_op27);
  assign p1_smul_89770_comb = smul32b_32b_x_32b(p0_TestBlock__A_op63, p0_TestBlock__B_op37);
  assign p1_smul_90301_comb = smul32b_32b_x_32b(p0_TestBlock__A_op64, p0_TestBlock__B_op47);
  assign p1_smul_90302_comb = smul32b_32b_x_32b(p0_TestBlock__A_op65, p0_TestBlock__B_op57);
  assign p1_smul_90303_comb = smul32b_32b_x_32b(p0_TestBlock__A_op66, p0_TestBlock__B_op67);
  assign p1_smul_90304_comb = smul32b_32b_x_32b(p0_TestBlock__A_op67, p0_TestBlock__B_op77);
  assign p1_smul_90305_comb = smul32b_32b_x_32b(p0_TestBlock__A_op68, p0_TestBlock__B_op87);
  assign p1_smul_90306_comb = smul32b_32b_x_32b(p0_TestBlock__A_op69, p0_TestBlock__B_op97);
  assign p1_smul_89771_comb = smul32b_32b_x_32b(p0_TestBlock__A_op60, p0_TestBlock__B_op8);
  assign p1_smul_89772_comb = smul32b_32b_x_32b(p0_TestBlock__A_op61, p0_TestBlock__B_op18);
  assign p1_smul_89773_comb = smul32b_32b_x_32b(p0_TestBlock__A_op62, p0_TestBlock__B_op28);
  assign p1_smul_89774_comb = smul32b_32b_x_32b(p0_TestBlock__A_op63, p0_TestBlock__B_op38);
  assign p1_smul_90307_comb = smul32b_32b_x_32b(p0_TestBlock__A_op64, p0_TestBlock__B_op48);
  assign p1_smul_90308_comb = smul32b_32b_x_32b(p0_TestBlock__A_op65, p0_TestBlock__B_op58);
  assign p1_smul_90309_comb = smul32b_32b_x_32b(p0_TestBlock__A_op66, p0_TestBlock__B_op68);
  assign p1_smul_90310_comb = smul32b_32b_x_32b(p0_TestBlock__A_op67, p0_TestBlock__B_op78);
  assign p1_smul_90311_comb = smul32b_32b_x_32b(p0_TestBlock__A_op68, p0_TestBlock__B_op88);
  assign p1_smul_90312_comb = smul32b_32b_x_32b(p0_TestBlock__A_op69, p0_TestBlock__B_op98);
  assign p1_smul_89775_comb = smul32b_32b_x_32b(p0_TestBlock__A_op60, p0_TestBlock__B_op9);
  assign p1_smul_89776_comb = smul32b_32b_x_32b(p0_TestBlock__A_op61, p0_TestBlock__B_op19);
  assign p1_smul_89777_comb = smul32b_32b_x_32b(p0_TestBlock__A_op62, p0_TestBlock__B_op29);
  assign p1_smul_89778_comb = smul32b_32b_x_32b(p0_TestBlock__A_op63, p0_TestBlock__B_op39);
  assign p1_smul_90313_comb = smul32b_32b_x_32b(p0_TestBlock__A_op64, p0_TestBlock__B_op49);
  assign p1_smul_90314_comb = smul32b_32b_x_32b(p0_TestBlock__A_op65, p0_TestBlock__B_op59);
  assign p1_smul_90315_comb = smul32b_32b_x_32b(p0_TestBlock__A_op66, p0_TestBlock__B_op69);
  assign p1_smul_90316_comb = smul32b_32b_x_32b(p0_TestBlock__A_op67, p0_TestBlock__B_op79);
  assign p1_smul_90317_comb = smul32b_32b_x_32b(p0_TestBlock__A_op68, p0_TestBlock__B_op89);
  assign p1_smul_90318_comb = smul32b_32b_x_32b(p0_TestBlock__A_op69, p0_TestBlock__B_op99);
  assign p1_smul_89779_comb = smul32b_32b_x_32b(p0_TestBlock__A_op70, p0_TestBlock__B_op0);
  assign p1_smul_89780_comb = smul32b_32b_x_32b(p0_TestBlock__A_op71, p0_TestBlock__B_op10);
  assign p1_smul_89781_comb = smul32b_32b_x_32b(p0_TestBlock__A_op72, p0_TestBlock__B_op20);
  assign p1_smul_89782_comb = smul32b_32b_x_32b(p0_TestBlock__A_op73, p0_TestBlock__B_op30);
  assign p1_smul_90319_comb = smul32b_32b_x_32b(p0_TestBlock__A_op74, p0_TestBlock__B_op40);
  assign p1_smul_90320_comb = smul32b_32b_x_32b(p0_TestBlock__A_op75, p0_TestBlock__B_op50);
  assign p1_smul_90321_comb = smul32b_32b_x_32b(p0_TestBlock__A_op76, p0_TestBlock__B_op60);
  assign p1_smul_90322_comb = smul32b_32b_x_32b(p0_TestBlock__A_op77, p0_TestBlock__B_op70);
  assign p1_smul_90323_comb = smul32b_32b_x_32b(p0_TestBlock__A_op78, p0_TestBlock__B_op80);
  assign p1_smul_90324_comb = smul32b_32b_x_32b(p0_TestBlock__A_op79, p0_TestBlock__B_op90);
  assign p1_smul_89783_comb = smul32b_32b_x_32b(p0_TestBlock__A_op70, p0_TestBlock__B_op1);
  assign p1_smul_89784_comb = smul32b_32b_x_32b(p0_TestBlock__A_op71, p0_TestBlock__B_op11);
  assign p1_smul_89785_comb = smul32b_32b_x_32b(p0_TestBlock__A_op72, p0_TestBlock__B_op21);
  assign p1_smul_89786_comb = smul32b_32b_x_32b(p0_TestBlock__A_op73, p0_TestBlock__B_op31);
  assign p1_smul_90325_comb = smul32b_32b_x_32b(p0_TestBlock__A_op74, p0_TestBlock__B_op41);
  assign p1_smul_90326_comb = smul32b_32b_x_32b(p0_TestBlock__A_op75, p0_TestBlock__B_op51);
  assign p1_smul_90327_comb = smul32b_32b_x_32b(p0_TestBlock__A_op76, p0_TestBlock__B_op61);
  assign p1_smul_90328_comb = smul32b_32b_x_32b(p0_TestBlock__A_op77, p0_TestBlock__B_op71);
  assign p1_smul_90329_comb = smul32b_32b_x_32b(p0_TestBlock__A_op78, p0_TestBlock__B_op81);
  assign p1_smul_90330_comb = smul32b_32b_x_32b(p0_TestBlock__A_op79, p0_TestBlock__B_op91);
  assign p1_smul_89787_comb = smul32b_32b_x_32b(p0_TestBlock__A_op70, p0_TestBlock__B_op2);
  assign p1_smul_89788_comb = smul32b_32b_x_32b(p0_TestBlock__A_op71, p0_TestBlock__B_op12);
  assign p1_smul_89789_comb = smul32b_32b_x_32b(p0_TestBlock__A_op72, p0_TestBlock__B_op22);
  assign p1_smul_89790_comb = smul32b_32b_x_32b(p0_TestBlock__A_op73, p0_TestBlock__B_op32);
  assign p1_smul_90331_comb = smul32b_32b_x_32b(p0_TestBlock__A_op74, p0_TestBlock__B_op42);
  assign p1_smul_90332_comb = smul32b_32b_x_32b(p0_TestBlock__A_op75, p0_TestBlock__B_op52);
  assign p1_smul_90333_comb = smul32b_32b_x_32b(p0_TestBlock__A_op76, p0_TestBlock__B_op62);
  assign p1_smul_90334_comb = smul32b_32b_x_32b(p0_TestBlock__A_op77, p0_TestBlock__B_op72);
  assign p1_smul_90335_comb = smul32b_32b_x_32b(p0_TestBlock__A_op78, p0_TestBlock__B_op82);
  assign p1_smul_90336_comb = smul32b_32b_x_32b(p0_TestBlock__A_op79, p0_TestBlock__B_op92);
  assign p1_smul_89791_comb = smul32b_32b_x_32b(p0_TestBlock__A_op70, p0_TestBlock__B_op3);
  assign p1_smul_89792_comb = smul32b_32b_x_32b(p0_TestBlock__A_op71, p0_TestBlock__B_op13);
  assign p1_smul_89793_comb = smul32b_32b_x_32b(p0_TestBlock__A_op72, p0_TestBlock__B_op23);
  assign p1_smul_89794_comb = smul32b_32b_x_32b(p0_TestBlock__A_op73, p0_TestBlock__B_op33);
  assign p1_smul_90337_comb = smul32b_32b_x_32b(p0_TestBlock__A_op74, p0_TestBlock__B_op43);
  assign p1_smul_90338_comb = smul32b_32b_x_32b(p0_TestBlock__A_op75, p0_TestBlock__B_op53);
  assign p1_smul_90339_comb = smul32b_32b_x_32b(p0_TestBlock__A_op76, p0_TestBlock__B_op63);
  assign p1_smul_90340_comb = smul32b_32b_x_32b(p0_TestBlock__A_op77, p0_TestBlock__B_op73);
  assign p1_smul_90341_comb = smul32b_32b_x_32b(p0_TestBlock__A_op78, p0_TestBlock__B_op83);
  assign p1_smul_90342_comb = smul32b_32b_x_32b(p0_TestBlock__A_op79, p0_TestBlock__B_op93);
  assign p1_smul_89795_comb = smul32b_32b_x_32b(p0_TestBlock__A_op70, p0_TestBlock__B_op4);
  assign p1_smul_89796_comb = smul32b_32b_x_32b(p0_TestBlock__A_op71, p0_TestBlock__B_op14);
  assign p1_smul_89797_comb = smul32b_32b_x_32b(p0_TestBlock__A_op72, p0_TestBlock__B_op24);
  assign p1_smul_89798_comb = smul32b_32b_x_32b(p0_TestBlock__A_op73, p0_TestBlock__B_op34);
  assign p1_smul_90343_comb = smul32b_32b_x_32b(p0_TestBlock__A_op74, p0_TestBlock__B_op44);
  assign p1_smul_90344_comb = smul32b_32b_x_32b(p0_TestBlock__A_op75, p0_TestBlock__B_op54);
  assign p1_smul_90345_comb = smul32b_32b_x_32b(p0_TestBlock__A_op76, p0_TestBlock__B_op64);
  assign p1_smul_90346_comb = smul32b_32b_x_32b(p0_TestBlock__A_op77, p0_TestBlock__B_op74);
  assign p1_smul_90347_comb = smul32b_32b_x_32b(p0_TestBlock__A_op78, p0_TestBlock__B_op84);
  assign p1_smul_90348_comb = smul32b_32b_x_32b(p0_TestBlock__A_op79, p0_TestBlock__B_op94);
  assign p1_smul_89799_comb = smul32b_32b_x_32b(p0_TestBlock__A_op70, p0_TestBlock__B_op5);
  assign p1_smul_89800_comb = smul32b_32b_x_32b(p0_TestBlock__A_op71, p0_TestBlock__B_op15);
  assign p1_smul_89801_comb = smul32b_32b_x_32b(p0_TestBlock__A_op72, p0_TestBlock__B_op25);
  assign p1_smul_89802_comb = smul32b_32b_x_32b(p0_TestBlock__A_op73, p0_TestBlock__B_op35);
  assign p1_smul_90349_comb = smul32b_32b_x_32b(p0_TestBlock__A_op74, p0_TestBlock__B_op45);
  assign p1_smul_90350_comb = smul32b_32b_x_32b(p0_TestBlock__A_op75, p0_TestBlock__B_op55);
  assign p1_smul_90351_comb = smul32b_32b_x_32b(p0_TestBlock__A_op76, p0_TestBlock__B_op65);
  assign p1_smul_90352_comb = smul32b_32b_x_32b(p0_TestBlock__A_op77, p0_TestBlock__B_op75);
  assign p1_smul_90353_comb = smul32b_32b_x_32b(p0_TestBlock__A_op78, p0_TestBlock__B_op85);
  assign p1_smul_90354_comb = smul32b_32b_x_32b(p0_TestBlock__A_op79, p0_TestBlock__B_op95);
  assign p1_smul_89803_comb = smul32b_32b_x_32b(p0_TestBlock__A_op70, p0_TestBlock__B_op6);
  assign p1_smul_89804_comb = smul32b_32b_x_32b(p0_TestBlock__A_op71, p0_TestBlock__B_op16);
  assign p1_smul_89805_comb = smul32b_32b_x_32b(p0_TestBlock__A_op72, p0_TestBlock__B_op26);
  assign p1_smul_89806_comb = smul32b_32b_x_32b(p0_TestBlock__A_op73, p0_TestBlock__B_op36);
  assign p1_smul_90355_comb = smul32b_32b_x_32b(p0_TestBlock__A_op74, p0_TestBlock__B_op46);
  assign p1_smul_90356_comb = smul32b_32b_x_32b(p0_TestBlock__A_op75, p0_TestBlock__B_op56);
  assign p1_smul_90357_comb = smul32b_32b_x_32b(p0_TestBlock__A_op76, p0_TestBlock__B_op66);
  assign p1_smul_90358_comb = smul32b_32b_x_32b(p0_TestBlock__A_op77, p0_TestBlock__B_op76);
  assign p1_smul_90359_comb = smul32b_32b_x_32b(p0_TestBlock__A_op78, p0_TestBlock__B_op86);
  assign p1_smul_90360_comb = smul32b_32b_x_32b(p0_TestBlock__A_op79, p0_TestBlock__B_op96);
  assign p1_smul_89807_comb = smul32b_32b_x_32b(p0_TestBlock__A_op70, p0_TestBlock__B_op7);
  assign p1_smul_89808_comb = smul32b_32b_x_32b(p0_TestBlock__A_op71, p0_TestBlock__B_op17);
  assign p1_smul_89809_comb = smul32b_32b_x_32b(p0_TestBlock__A_op72, p0_TestBlock__B_op27);
  assign p1_smul_89810_comb = smul32b_32b_x_32b(p0_TestBlock__A_op73, p0_TestBlock__B_op37);
  assign p1_smul_90361_comb = smul32b_32b_x_32b(p0_TestBlock__A_op74, p0_TestBlock__B_op47);
  assign p1_smul_90362_comb = smul32b_32b_x_32b(p0_TestBlock__A_op75, p0_TestBlock__B_op57);
  assign p1_smul_90363_comb = smul32b_32b_x_32b(p0_TestBlock__A_op76, p0_TestBlock__B_op67);
  assign p1_smul_90364_comb = smul32b_32b_x_32b(p0_TestBlock__A_op77, p0_TestBlock__B_op77);
  assign p1_smul_90365_comb = smul32b_32b_x_32b(p0_TestBlock__A_op78, p0_TestBlock__B_op87);
  assign p1_smul_90366_comb = smul32b_32b_x_32b(p0_TestBlock__A_op79, p0_TestBlock__B_op97);
  assign p1_smul_89811_comb = smul32b_32b_x_32b(p0_TestBlock__A_op70, p0_TestBlock__B_op8);
  assign p1_smul_89812_comb = smul32b_32b_x_32b(p0_TestBlock__A_op71, p0_TestBlock__B_op18);
  assign p1_smul_89813_comb = smul32b_32b_x_32b(p0_TestBlock__A_op72, p0_TestBlock__B_op28);
  assign p1_smul_89814_comb = smul32b_32b_x_32b(p0_TestBlock__A_op73, p0_TestBlock__B_op38);
  assign p1_smul_90367_comb = smul32b_32b_x_32b(p0_TestBlock__A_op74, p0_TestBlock__B_op48);
  assign p1_smul_90368_comb = smul32b_32b_x_32b(p0_TestBlock__A_op75, p0_TestBlock__B_op58);
  assign p1_smul_90369_comb = smul32b_32b_x_32b(p0_TestBlock__A_op76, p0_TestBlock__B_op68);
  assign p1_smul_90370_comb = smul32b_32b_x_32b(p0_TestBlock__A_op77, p0_TestBlock__B_op78);
  assign p1_smul_90371_comb = smul32b_32b_x_32b(p0_TestBlock__A_op78, p0_TestBlock__B_op88);
  assign p1_smul_90372_comb = smul32b_32b_x_32b(p0_TestBlock__A_op79, p0_TestBlock__B_op98);
  assign p1_smul_89815_comb = smul32b_32b_x_32b(p0_TestBlock__A_op70, p0_TestBlock__B_op9);
  assign p1_smul_89816_comb = smul32b_32b_x_32b(p0_TestBlock__A_op71, p0_TestBlock__B_op19);
  assign p1_smul_89817_comb = smul32b_32b_x_32b(p0_TestBlock__A_op72, p0_TestBlock__B_op29);
  assign p1_smul_89818_comb = smul32b_32b_x_32b(p0_TestBlock__A_op73, p0_TestBlock__B_op39);
  assign p1_smul_90373_comb = smul32b_32b_x_32b(p0_TestBlock__A_op74, p0_TestBlock__B_op49);
  assign p1_smul_90374_comb = smul32b_32b_x_32b(p0_TestBlock__A_op75, p0_TestBlock__B_op59);
  assign p1_smul_90375_comb = smul32b_32b_x_32b(p0_TestBlock__A_op76, p0_TestBlock__B_op69);
  assign p1_smul_90376_comb = smul32b_32b_x_32b(p0_TestBlock__A_op77, p0_TestBlock__B_op79);
  assign p1_smul_90377_comb = smul32b_32b_x_32b(p0_TestBlock__A_op78, p0_TestBlock__B_op89);
  assign p1_smul_90378_comb = smul32b_32b_x_32b(p0_TestBlock__A_op79, p0_TestBlock__B_op99);
  assign p1_smul_89819_comb = smul32b_32b_x_32b(p0_TestBlock__A_op80, p0_TestBlock__B_op0);
  assign p1_smul_89820_comb = smul32b_32b_x_32b(p0_TestBlock__A_op81, p0_TestBlock__B_op10);
  assign p1_smul_89821_comb = smul32b_32b_x_32b(p0_TestBlock__A_op82, p0_TestBlock__B_op20);
  assign p1_smul_89822_comb = smul32b_32b_x_32b(p0_TestBlock__A_op83, p0_TestBlock__B_op30);
  assign p1_smul_90379_comb = smul32b_32b_x_32b(p0_TestBlock__A_op84, p0_TestBlock__B_op40);
  assign p1_smul_90380_comb = smul32b_32b_x_32b(p0_TestBlock__A_op85, p0_TestBlock__B_op50);
  assign p1_smul_90381_comb = smul32b_32b_x_32b(p0_TestBlock__A_op86, p0_TestBlock__B_op60);
  assign p1_smul_90382_comb = smul32b_32b_x_32b(p0_TestBlock__A_op87, p0_TestBlock__B_op70);
  assign p1_smul_90383_comb = smul32b_32b_x_32b(p0_TestBlock__A_op88, p0_TestBlock__B_op80);
  assign p1_smul_90384_comb = smul32b_32b_x_32b(p0_TestBlock__A_op89, p0_TestBlock__B_op90);
  assign p1_smul_89823_comb = smul32b_32b_x_32b(p0_TestBlock__A_op80, p0_TestBlock__B_op1);
  assign p1_smul_89824_comb = smul32b_32b_x_32b(p0_TestBlock__A_op81, p0_TestBlock__B_op11);
  assign p1_smul_89825_comb = smul32b_32b_x_32b(p0_TestBlock__A_op82, p0_TestBlock__B_op21);
  assign p1_smul_89826_comb = smul32b_32b_x_32b(p0_TestBlock__A_op83, p0_TestBlock__B_op31);
  assign p1_smul_90385_comb = smul32b_32b_x_32b(p0_TestBlock__A_op84, p0_TestBlock__B_op41);
  assign p1_smul_90386_comb = smul32b_32b_x_32b(p0_TestBlock__A_op85, p0_TestBlock__B_op51);
  assign p1_smul_90387_comb = smul32b_32b_x_32b(p0_TestBlock__A_op86, p0_TestBlock__B_op61);
  assign p1_smul_90388_comb = smul32b_32b_x_32b(p0_TestBlock__A_op87, p0_TestBlock__B_op71);
  assign p1_smul_90389_comb = smul32b_32b_x_32b(p0_TestBlock__A_op88, p0_TestBlock__B_op81);
  assign p1_smul_90390_comb = smul32b_32b_x_32b(p0_TestBlock__A_op89, p0_TestBlock__B_op91);
  assign p1_smul_89827_comb = smul32b_32b_x_32b(p0_TestBlock__A_op80, p0_TestBlock__B_op2);
  assign p1_smul_89828_comb = smul32b_32b_x_32b(p0_TestBlock__A_op81, p0_TestBlock__B_op12);
  assign p1_smul_89829_comb = smul32b_32b_x_32b(p0_TestBlock__A_op82, p0_TestBlock__B_op22);
  assign p1_smul_89830_comb = smul32b_32b_x_32b(p0_TestBlock__A_op83, p0_TestBlock__B_op32);
  assign p1_smul_90391_comb = smul32b_32b_x_32b(p0_TestBlock__A_op84, p0_TestBlock__B_op42);
  assign p1_smul_90392_comb = smul32b_32b_x_32b(p0_TestBlock__A_op85, p0_TestBlock__B_op52);
  assign p1_smul_90393_comb = smul32b_32b_x_32b(p0_TestBlock__A_op86, p0_TestBlock__B_op62);
  assign p1_smul_90394_comb = smul32b_32b_x_32b(p0_TestBlock__A_op87, p0_TestBlock__B_op72);
  assign p1_smul_90395_comb = smul32b_32b_x_32b(p0_TestBlock__A_op88, p0_TestBlock__B_op82);
  assign p1_smul_90396_comb = smul32b_32b_x_32b(p0_TestBlock__A_op89, p0_TestBlock__B_op92);
  assign p1_smul_89831_comb = smul32b_32b_x_32b(p0_TestBlock__A_op80, p0_TestBlock__B_op3);
  assign p1_smul_89832_comb = smul32b_32b_x_32b(p0_TestBlock__A_op81, p0_TestBlock__B_op13);
  assign p1_smul_89833_comb = smul32b_32b_x_32b(p0_TestBlock__A_op82, p0_TestBlock__B_op23);
  assign p1_smul_89834_comb = smul32b_32b_x_32b(p0_TestBlock__A_op83, p0_TestBlock__B_op33);
  assign p1_smul_90397_comb = smul32b_32b_x_32b(p0_TestBlock__A_op84, p0_TestBlock__B_op43);
  assign p1_smul_90398_comb = smul32b_32b_x_32b(p0_TestBlock__A_op85, p0_TestBlock__B_op53);
  assign p1_smul_90399_comb = smul32b_32b_x_32b(p0_TestBlock__A_op86, p0_TestBlock__B_op63);
  assign p1_smul_90400_comb = smul32b_32b_x_32b(p0_TestBlock__A_op87, p0_TestBlock__B_op73);
  assign p1_smul_90401_comb = smul32b_32b_x_32b(p0_TestBlock__A_op88, p0_TestBlock__B_op83);
  assign p1_smul_90402_comb = smul32b_32b_x_32b(p0_TestBlock__A_op89, p0_TestBlock__B_op93);
  assign p1_smul_89835_comb = smul32b_32b_x_32b(p0_TestBlock__A_op80, p0_TestBlock__B_op4);
  assign p1_smul_89836_comb = smul32b_32b_x_32b(p0_TestBlock__A_op81, p0_TestBlock__B_op14);
  assign p1_smul_89837_comb = smul32b_32b_x_32b(p0_TestBlock__A_op82, p0_TestBlock__B_op24);
  assign p1_smul_89838_comb = smul32b_32b_x_32b(p0_TestBlock__A_op83, p0_TestBlock__B_op34);
  assign p1_smul_90403_comb = smul32b_32b_x_32b(p0_TestBlock__A_op84, p0_TestBlock__B_op44);
  assign p1_smul_90404_comb = smul32b_32b_x_32b(p0_TestBlock__A_op85, p0_TestBlock__B_op54);
  assign p1_smul_90405_comb = smul32b_32b_x_32b(p0_TestBlock__A_op86, p0_TestBlock__B_op64);
  assign p1_smul_90406_comb = smul32b_32b_x_32b(p0_TestBlock__A_op87, p0_TestBlock__B_op74);
  assign p1_smul_90407_comb = smul32b_32b_x_32b(p0_TestBlock__A_op88, p0_TestBlock__B_op84);
  assign p1_smul_90408_comb = smul32b_32b_x_32b(p0_TestBlock__A_op89, p0_TestBlock__B_op94);
  assign p1_smul_89839_comb = smul32b_32b_x_32b(p0_TestBlock__A_op80, p0_TestBlock__B_op5);
  assign p1_smul_89840_comb = smul32b_32b_x_32b(p0_TestBlock__A_op81, p0_TestBlock__B_op15);
  assign p1_smul_89841_comb = smul32b_32b_x_32b(p0_TestBlock__A_op82, p0_TestBlock__B_op25);
  assign p1_smul_89842_comb = smul32b_32b_x_32b(p0_TestBlock__A_op83, p0_TestBlock__B_op35);
  assign p1_smul_90409_comb = smul32b_32b_x_32b(p0_TestBlock__A_op84, p0_TestBlock__B_op45);
  assign p1_smul_90410_comb = smul32b_32b_x_32b(p0_TestBlock__A_op85, p0_TestBlock__B_op55);
  assign p1_smul_90411_comb = smul32b_32b_x_32b(p0_TestBlock__A_op86, p0_TestBlock__B_op65);
  assign p1_smul_90412_comb = smul32b_32b_x_32b(p0_TestBlock__A_op87, p0_TestBlock__B_op75);
  assign p1_smul_90413_comb = smul32b_32b_x_32b(p0_TestBlock__A_op88, p0_TestBlock__B_op85);
  assign p1_smul_90414_comb = smul32b_32b_x_32b(p0_TestBlock__A_op89, p0_TestBlock__B_op95);
  assign p1_smul_89843_comb = smul32b_32b_x_32b(p0_TestBlock__A_op80, p0_TestBlock__B_op6);
  assign p1_smul_89844_comb = smul32b_32b_x_32b(p0_TestBlock__A_op81, p0_TestBlock__B_op16);
  assign p1_smul_89845_comb = smul32b_32b_x_32b(p0_TestBlock__A_op82, p0_TestBlock__B_op26);
  assign p1_smul_89846_comb = smul32b_32b_x_32b(p0_TestBlock__A_op83, p0_TestBlock__B_op36);
  assign p1_smul_90415_comb = smul32b_32b_x_32b(p0_TestBlock__A_op84, p0_TestBlock__B_op46);
  assign p1_smul_90416_comb = smul32b_32b_x_32b(p0_TestBlock__A_op85, p0_TestBlock__B_op56);
  assign p1_smul_90417_comb = smul32b_32b_x_32b(p0_TestBlock__A_op86, p0_TestBlock__B_op66);
  assign p1_smul_90418_comb = smul32b_32b_x_32b(p0_TestBlock__A_op87, p0_TestBlock__B_op76);
  assign p1_smul_90419_comb = smul32b_32b_x_32b(p0_TestBlock__A_op88, p0_TestBlock__B_op86);
  assign p1_smul_90420_comb = smul32b_32b_x_32b(p0_TestBlock__A_op89, p0_TestBlock__B_op96);
  assign p1_smul_89847_comb = smul32b_32b_x_32b(p0_TestBlock__A_op80, p0_TestBlock__B_op7);
  assign p1_smul_89848_comb = smul32b_32b_x_32b(p0_TestBlock__A_op81, p0_TestBlock__B_op17);
  assign p1_smul_89849_comb = smul32b_32b_x_32b(p0_TestBlock__A_op82, p0_TestBlock__B_op27);
  assign p1_smul_89850_comb = smul32b_32b_x_32b(p0_TestBlock__A_op83, p0_TestBlock__B_op37);
  assign p1_smul_90421_comb = smul32b_32b_x_32b(p0_TestBlock__A_op84, p0_TestBlock__B_op47);
  assign p1_smul_90422_comb = smul32b_32b_x_32b(p0_TestBlock__A_op85, p0_TestBlock__B_op57);
  assign p1_smul_90423_comb = smul32b_32b_x_32b(p0_TestBlock__A_op86, p0_TestBlock__B_op67);
  assign p1_smul_90424_comb = smul32b_32b_x_32b(p0_TestBlock__A_op87, p0_TestBlock__B_op77);
  assign p1_smul_90425_comb = smul32b_32b_x_32b(p0_TestBlock__A_op88, p0_TestBlock__B_op87);
  assign p1_smul_90426_comb = smul32b_32b_x_32b(p0_TestBlock__A_op89, p0_TestBlock__B_op97);
  assign p1_smul_89851_comb = smul32b_32b_x_32b(p0_TestBlock__A_op80, p0_TestBlock__B_op8);
  assign p1_smul_89852_comb = smul32b_32b_x_32b(p0_TestBlock__A_op81, p0_TestBlock__B_op18);
  assign p1_smul_89853_comb = smul32b_32b_x_32b(p0_TestBlock__A_op82, p0_TestBlock__B_op28);
  assign p1_smul_89854_comb = smul32b_32b_x_32b(p0_TestBlock__A_op83, p0_TestBlock__B_op38);
  assign p1_smul_90427_comb = smul32b_32b_x_32b(p0_TestBlock__A_op84, p0_TestBlock__B_op48);
  assign p1_smul_90428_comb = smul32b_32b_x_32b(p0_TestBlock__A_op85, p0_TestBlock__B_op58);
  assign p1_smul_90429_comb = smul32b_32b_x_32b(p0_TestBlock__A_op86, p0_TestBlock__B_op68);
  assign p1_smul_90430_comb = smul32b_32b_x_32b(p0_TestBlock__A_op87, p0_TestBlock__B_op78);
  assign p1_smul_90431_comb = smul32b_32b_x_32b(p0_TestBlock__A_op88, p0_TestBlock__B_op88);
  assign p1_smul_90432_comb = smul32b_32b_x_32b(p0_TestBlock__A_op89, p0_TestBlock__B_op98);
  assign p1_smul_89855_comb = smul32b_32b_x_32b(p0_TestBlock__A_op80, p0_TestBlock__B_op9);
  assign p1_smul_89856_comb = smul32b_32b_x_32b(p0_TestBlock__A_op81, p0_TestBlock__B_op19);
  assign p1_smul_89857_comb = smul32b_32b_x_32b(p0_TestBlock__A_op82, p0_TestBlock__B_op29);
  assign p1_smul_89858_comb = smul32b_32b_x_32b(p0_TestBlock__A_op83, p0_TestBlock__B_op39);
  assign p1_smul_90433_comb = smul32b_32b_x_32b(p0_TestBlock__A_op84, p0_TestBlock__B_op49);
  assign p1_smul_90434_comb = smul32b_32b_x_32b(p0_TestBlock__A_op85, p0_TestBlock__B_op59);
  assign p1_smul_90435_comb = smul32b_32b_x_32b(p0_TestBlock__A_op86, p0_TestBlock__B_op69);
  assign p1_smul_90436_comb = smul32b_32b_x_32b(p0_TestBlock__A_op87, p0_TestBlock__B_op79);
  assign p1_smul_90437_comb = smul32b_32b_x_32b(p0_TestBlock__A_op88, p0_TestBlock__B_op89);
  assign p1_smul_90438_comb = smul32b_32b_x_32b(p0_TestBlock__A_op89, p0_TestBlock__B_op99);
  assign p1_smul_89859_comb = smul32b_32b_x_32b(p0_TestBlock__A_op90, p0_TestBlock__B_op0);
  assign p1_smul_89860_comb = smul32b_32b_x_32b(p0_TestBlock__A_op91, p0_TestBlock__B_op10);
  assign p1_smul_89861_comb = smul32b_32b_x_32b(p0_TestBlock__A_op92, p0_TestBlock__B_op20);
  assign p1_smul_89862_comb = smul32b_32b_x_32b(p0_TestBlock__A_op93, p0_TestBlock__B_op30);
  assign p1_smul_90439_comb = smul32b_32b_x_32b(p0_TestBlock__A_op94, p0_TestBlock__B_op40);
  assign p1_smul_90440_comb = smul32b_32b_x_32b(p0_TestBlock__A_op95, p0_TestBlock__B_op50);
  assign p1_smul_90441_comb = smul32b_32b_x_32b(p0_TestBlock__A_op96, p0_TestBlock__B_op60);
  assign p1_smul_90442_comb = smul32b_32b_x_32b(p0_TestBlock__A_op97, p0_TestBlock__B_op70);
  assign p1_smul_90443_comb = smul32b_32b_x_32b(p0_TestBlock__A_op98, p0_TestBlock__B_op80);
  assign p1_smul_90444_comb = smul32b_32b_x_32b(p0_TestBlock__A_op99, p0_TestBlock__B_op90);
  assign p1_smul_89863_comb = smul32b_32b_x_32b(p0_TestBlock__A_op90, p0_TestBlock__B_op1);
  assign p1_smul_89864_comb = smul32b_32b_x_32b(p0_TestBlock__A_op91, p0_TestBlock__B_op11);
  assign p1_smul_89865_comb = smul32b_32b_x_32b(p0_TestBlock__A_op92, p0_TestBlock__B_op21);
  assign p1_smul_89866_comb = smul32b_32b_x_32b(p0_TestBlock__A_op93, p0_TestBlock__B_op31);
  assign p1_smul_90445_comb = smul32b_32b_x_32b(p0_TestBlock__A_op94, p0_TestBlock__B_op41);
  assign p1_smul_90446_comb = smul32b_32b_x_32b(p0_TestBlock__A_op95, p0_TestBlock__B_op51);
  assign p1_smul_90447_comb = smul32b_32b_x_32b(p0_TestBlock__A_op96, p0_TestBlock__B_op61);
  assign p1_smul_90448_comb = smul32b_32b_x_32b(p0_TestBlock__A_op97, p0_TestBlock__B_op71);
  assign p1_smul_90449_comb = smul32b_32b_x_32b(p0_TestBlock__A_op98, p0_TestBlock__B_op81);
  assign p1_smul_90450_comb = smul32b_32b_x_32b(p0_TestBlock__A_op99, p0_TestBlock__B_op91);
  assign p1_smul_89867_comb = smul32b_32b_x_32b(p0_TestBlock__A_op90, p0_TestBlock__B_op2);
  assign p1_smul_89868_comb = smul32b_32b_x_32b(p0_TestBlock__A_op91, p0_TestBlock__B_op12);
  assign p1_smul_89869_comb = smul32b_32b_x_32b(p0_TestBlock__A_op92, p0_TestBlock__B_op22);
  assign p1_smul_89870_comb = smul32b_32b_x_32b(p0_TestBlock__A_op93, p0_TestBlock__B_op32);
  assign p1_smul_90451_comb = smul32b_32b_x_32b(p0_TestBlock__A_op94, p0_TestBlock__B_op42);
  assign p1_smul_90452_comb = smul32b_32b_x_32b(p0_TestBlock__A_op95, p0_TestBlock__B_op52);
  assign p1_smul_90453_comb = smul32b_32b_x_32b(p0_TestBlock__A_op96, p0_TestBlock__B_op62);
  assign p1_smul_90454_comb = smul32b_32b_x_32b(p0_TestBlock__A_op97, p0_TestBlock__B_op72);
  assign p1_smul_90455_comb = smul32b_32b_x_32b(p0_TestBlock__A_op98, p0_TestBlock__B_op82);
  assign p1_smul_90456_comb = smul32b_32b_x_32b(p0_TestBlock__A_op99, p0_TestBlock__B_op92);
  assign p1_smul_89871_comb = smul32b_32b_x_32b(p0_TestBlock__A_op90, p0_TestBlock__B_op3);
  assign p1_smul_89872_comb = smul32b_32b_x_32b(p0_TestBlock__A_op91, p0_TestBlock__B_op13);
  assign p1_smul_89873_comb = smul32b_32b_x_32b(p0_TestBlock__A_op92, p0_TestBlock__B_op23);
  assign p1_smul_89874_comb = smul32b_32b_x_32b(p0_TestBlock__A_op93, p0_TestBlock__B_op33);
  assign p1_smul_90457_comb = smul32b_32b_x_32b(p0_TestBlock__A_op94, p0_TestBlock__B_op43);
  assign p1_smul_90458_comb = smul32b_32b_x_32b(p0_TestBlock__A_op95, p0_TestBlock__B_op53);
  assign p1_smul_90459_comb = smul32b_32b_x_32b(p0_TestBlock__A_op96, p0_TestBlock__B_op63);
  assign p1_smul_90460_comb = smul32b_32b_x_32b(p0_TestBlock__A_op97, p0_TestBlock__B_op73);
  assign p1_smul_90461_comb = smul32b_32b_x_32b(p0_TestBlock__A_op98, p0_TestBlock__B_op83);
  assign p1_smul_90462_comb = smul32b_32b_x_32b(p0_TestBlock__A_op99, p0_TestBlock__B_op93);
  assign p1_smul_89875_comb = smul32b_32b_x_32b(p0_TestBlock__A_op90, p0_TestBlock__B_op4);
  assign p1_smul_89876_comb = smul32b_32b_x_32b(p0_TestBlock__A_op91, p0_TestBlock__B_op14);
  assign p1_smul_89877_comb = smul32b_32b_x_32b(p0_TestBlock__A_op92, p0_TestBlock__B_op24);
  assign p1_smul_89878_comb = smul32b_32b_x_32b(p0_TestBlock__A_op93, p0_TestBlock__B_op34);
  assign p1_smul_90463_comb = smul32b_32b_x_32b(p0_TestBlock__A_op94, p0_TestBlock__B_op44);
  assign p1_smul_90464_comb = smul32b_32b_x_32b(p0_TestBlock__A_op95, p0_TestBlock__B_op54);
  assign p1_smul_90465_comb = smul32b_32b_x_32b(p0_TestBlock__A_op96, p0_TestBlock__B_op64);
  assign p1_smul_90466_comb = smul32b_32b_x_32b(p0_TestBlock__A_op97, p0_TestBlock__B_op74);
  assign p1_smul_90467_comb = smul32b_32b_x_32b(p0_TestBlock__A_op98, p0_TestBlock__B_op84);
  assign p1_smul_90468_comb = smul32b_32b_x_32b(p0_TestBlock__A_op99, p0_TestBlock__B_op94);
  assign p1_smul_89879_comb = smul32b_32b_x_32b(p0_TestBlock__A_op90, p0_TestBlock__B_op5);
  assign p1_smul_89880_comb = smul32b_32b_x_32b(p0_TestBlock__A_op91, p0_TestBlock__B_op15);
  assign p1_smul_89881_comb = smul32b_32b_x_32b(p0_TestBlock__A_op92, p0_TestBlock__B_op25);
  assign p1_smul_89882_comb = smul32b_32b_x_32b(p0_TestBlock__A_op93, p0_TestBlock__B_op35);
  assign p1_smul_90469_comb = smul32b_32b_x_32b(p0_TestBlock__A_op94, p0_TestBlock__B_op45);
  assign p1_smul_90470_comb = smul32b_32b_x_32b(p0_TestBlock__A_op95, p0_TestBlock__B_op55);
  assign p1_smul_90471_comb = smul32b_32b_x_32b(p0_TestBlock__A_op96, p0_TestBlock__B_op65);
  assign p1_smul_90472_comb = smul32b_32b_x_32b(p0_TestBlock__A_op97, p0_TestBlock__B_op75);
  assign p1_smul_90473_comb = smul32b_32b_x_32b(p0_TestBlock__A_op98, p0_TestBlock__B_op85);
  assign p1_smul_90474_comb = smul32b_32b_x_32b(p0_TestBlock__A_op99, p0_TestBlock__B_op95);
  assign p1_smul_89883_comb = smul32b_32b_x_32b(p0_TestBlock__A_op90, p0_TestBlock__B_op6);
  assign p1_smul_89884_comb = smul32b_32b_x_32b(p0_TestBlock__A_op91, p0_TestBlock__B_op16);
  assign p1_smul_89885_comb = smul32b_32b_x_32b(p0_TestBlock__A_op92, p0_TestBlock__B_op26);
  assign p1_smul_89886_comb = smul32b_32b_x_32b(p0_TestBlock__A_op93, p0_TestBlock__B_op36);
  assign p1_smul_90475_comb = smul32b_32b_x_32b(p0_TestBlock__A_op94, p0_TestBlock__B_op46);
  assign p1_smul_90476_comb = smul32b_32b_x_32b(p0_TestBlock__A_op95, p0_TestBlock__B_op56);
  assign p1_smul_90477_comb = smul32b_32b_x_32b(p0_TestBlock__A_op96, p0_TestBlock__B_op66);
  assign p1_smul_90478_comb = smul32b_32b_x_32b(p0_TestBlock__A_op97, p0_TestBlock__B_op76);
  assign p1_smul_90479_comb = smul32b_32b_x_32b(p0_TestBlock__A_op98, p0_TestBlock__B_op86);
  assign p1_smul_90480_comb = smul32b_32b_x_32b(p0_TestBlock__A_op99, p0_TestBlock__B_op96);
  assign p1_smul_89887_comb = smul32b_32b_x_32b(p0_TestBlock__A_op90, p0_TestBlock__B_op7);
  assign p1_smul_89888_comb = smul32b_32b_x_32b(p0_TestBlock__A_op91, p0_TestBlock__B_op17);
  assign p1_smul_89889_comb = smul32b_32b_x_32b(p0_TestBlock__A_op92, p0_TestBlock__B_op27);
  assign p1_smul_89890_comb = smul32b_32b_x_32b(p0_TestBlock__A_op93, p0_TestBlock__B_op37);
  assign p1_smul_90481_comb = smul32b_32b_x_32b(p0_TestBlock__A_op94, p0_TestBlock__B_op47);
  assign p1_smul_90482_comb = smul32b_32b_x_32b(p0_TestBlock__A_op95, p0_TestBlock__B_op57);
  assign p1_smul_90483_comb = smul32b_32b_x_32b(p0_TestBlock__A_op96, p0_TestBlock__B_op67);
  assign p1_smul_90484_comb = smul32b_32b_x_32b(p0_TestBlock__A_op97, p0_TestBlock__B_op77);
  assign p1_smul_90485_comb = smul32b_32b_x_32b(p0_TestBlock__A_op98, p0_TestBlock__B_op87);
  assign p1_smul_90486_comb = smul32b_32b_x_32b(p0_TestBlock__A_op99, p0_TestBlock__B_op97);
  assign p1_smul_89891_comb = smul32b_32b_x_32b(p0_TestBlock__A_op90, p0_TestBlock__B_op8);
  assign p1_smul_89892_comb = smul32b_32b_x_32b(p0_TestBlock__A_op91, p0_TestBlock__B_op18);
  assign p1_smul_89893_comb = smul32b_32b_x_32b(p0_TestBlock__A_op92, p0_TestBlock__B_op28);
  assign p1_smul_89894_comb = smul32b_32b_x_32b(p0_TestBlock__A_op93, p0_TestBlock__B_op38);
  assign p1_smul_90487_comb = smul32b_32b_x_32b(p0_TestBlock__A_op94, p0_TestBlock__B_op48);
  assign p1_smul_90488_comb = smul32b_32b_x_32b(p0_TestBlock__A_op95, p0_TestBlock__B_op58);
  assign p1_smul_90489_comb = smul32b_32b_x_32b(p0_TestBlock__A_op96, p0_TestBlock__B_op68);
  assign p1_smul_90490_comb = smul32b_32b_x_32b(p0_TestBlock__A_op97, p0_TestBlock__B_op78);
  assign p1_smul_90491_comb = smul32b_32b_x_32b(p0_TestBlock__A_op98, p0_TestBlock__B_op88);
  assign p1_smul_90492_comb = smul32b_32b_x_32b(p0_TestBlock__A_op99, p0_TestBlock__B_op98);
  assign p1_smul_89895_comb = smul32b_32b_x_32b(p0_TestBlock__A_op90, p0_TestBlock__B_op9);
  assign p1_smul_89896_comb = smul32b_32b_x_32b(p0_TestBlock__A_op91, p0_TestBlock__B_op19);
  assign p1_smul_89897_comb = smul32b_32b_x_32b(p0_TestBlock__A_op92, p0_TestBlock__B_op29);
  assign p1_smul_89898_comb = smul32b_32b_x_32b(p0_TestBlock__A_op93, p0_TestBlock__B_op39);
  assign p1_smul_90493_comb = smul32b_32b_x_32b(p0_TestBlock__A_op94, p0_TestBlock__B_op49);
  assign p1_smul_90494_comb = smul32b_32b_x_32b(p0_TestBlock__A_op95, p0_TestBlock__B_op59);
  assign p1_smul_90495_comb = smul32b_32b_x_32b(p0_TestBlock__A_op96, p0_TestBlock__B_op69);
  assign p1_smul_90496_comb = smul32b_32b_x_32b(p0_TestBlock__A_op97, p0_TestBlock__B_op79);
  assign p1_smul_90497_comb = smul32b_32b_x_32b(p0_TestBlock__A_op98, p0_TestBlock__B_op89);
  assign p1_smul_90498_comb = smul32b_32b_x_32b(p0_TestBlock__A_op99, p0_TestBlock__B_op99);

  // Registers for pipe stage 1:
  reg [31:0] p1_smul_89499;
  reg [31:0] p1_smul_89500;
  reg [31:0] p1_smul_89501;
  reg [31:0] p1_smul_89502;
  reg [31:0] p1_smul_89899;
  reg [31:0] p1_smul_89900;
  reg [31:0] p1_smul_89901;
  reg [31:0] p1_smul_89902;
  reg [31:0] p1_smul_89903;
  reg [31:0] p1_smul_89904;
  reg [31:0] p1_smul_89503;
  reg [31:0] p1_smul_89504;
  reg [31:0] p1_smul_89505;
  reg [31:0] p1_smul_89506;
  reg [31:0] p1_smul_89905;
  reg [31:0] p1_smul_89906;
  reg [31:0] p1_smul_89907;
  reg [31:0] p1_smul_89908;
  reg [31:0] p1_smul_89909;
  reg [31:0] p1_smul_89910;
  reg [31:0] p1_smul_89507;
  reg [31:0] p1_smul_89508;
  reg [31:0] p1_smul_89509;
  reg [31:0] p1_smul_89510;
  reg [31:0] p1_smul_89911;
  reg [31:0] p1_smul_89912;
  reg [31:0] p1_smul_89913;
  reg [31:0] p1_smul_89914;
  reg [31:0] p1_smul_89915;
  reg [31:0] p1_smul_89916;
  reg [31:0] p1_smul_89511;
  reg [31:0] p1_smul_89512;
  reg [31:0] p1_smul_89513;
  reg [31:0] p1_smul_89514;
  reg [31:0] p1_smul_89917;
  reg [31:0] p1_smul_89918;
  reg [31:0] p1_smul_89919;
  reg [31:0] p1_smul_89920;
  reg [31:0] p1_smul_89921;
  reg [31:0] p1_smul_89922;
  reg [31:0] p1_smul_89515;
  reg [31:0] p1_smul_89516;
  reg [31:0] p1_smul_89517;
  reg [31:0] p1_smul_89518;
  reg [31:0] p1_smul_89923;
  reg [31:0] p1_smul_89924;
  reg [31:0] p1_smul_89925;
  reg [31:0] p1_smul_89926;
  reg [31:0] p1_smul_89927;
  reg [31:0] p1_smul_89928;
  reg [31:0] p1_smul_89519;
  reg [31:0] p1_smul_89520;
  reg [31:0] p1_smul_89521;
  reg [31:0] p1_smul_89522;
  reg [31:0] p1_smul_89929;
  reg [31:0] p1_smul_89930;
  reg [31:0] p1_smul_89931;
  reg [31:0] p1_smul_89932;
  reg [31:0] p1_smul_89933;
  reg [31:0] p1_smul_89934;
  reg [31:0] p1_smul_89523;
  reg [31:0] p1_smul_89524;
  reg [31:0] p1_smul_89525;
  reg [31:0] p1_smul_89526;
  reg [31:0] p1_smul_89935;
  reg [31:0] p1_smul_89936;
  reg [31:0] p1_smul_89937;
  reg [31:0] p1_smul_89938;
  reg [31:0] p1_smul_89939;
  reg [31:0] p1_smul_89940;
  reg [31:0] p1_smul_89527;
  reg [31:0] p1_smul_89528;
  reg [31:0] p1_smul_89529;
  reg [31:0] p1_smul_89530;
  reg [31:0] p1_smul_89941;
  reg [31:0] p1_smul_89942;
  reg [31:0] p1_smul_89943;
  reg [31:0] p1_smul_89944;
  reg [31:0] p1_smul_89945;
  reg [31:0] p1_smul_89946;
  reg [31:0] p1_smul_89531;
  reg [31:0] p1_smul_89532;
  reg [31:0] p1_smul_89533;
  reg [31:0] p1_smul_89534;
  reg [31:0] p1_smul_89947;
  reg [31:0] p1_smul_89948;
  reg [31:0] p1_smul_89949;
  reg [31:0] p1_smul_89950;
  reg [31:0] p1_smul_89951;
  reg [31:0] p1_smul_89952;
  reg [31:0] p1_smul_89535;
  reg [31:0] p1_smul_89536;
  reg [31:0] p1_smul_89537;
  reg [31:0] p1_smul_89538;
  reg [31:0] p1_smul_89953;
  reg [31:0] p1_smul_89954;
  reg [31:0] p1_smul_89955;
  reg [31:0] p1_smul_89956;
  reg [31:0] p1_smul_89957;
  reg [31:0] p1_smul_89958;
  reg [31:0] p1_smul_89539;
  reg [31:0] p1_smul_89540;
  reg [31:0] p1_smul_89541;
  reg [31:0] p1_smul_89542;
  reg [31:0] p1_smul_89959;
  reg [31:0] p1_smul_89960;
  reg [31:0] p1_smul_89961;
  reg [31:0] p1_smul_89962;
  reg [31:0] p1_smul_89963;
  reg [31:0] p1_smul_89964;
  reg [31:0] p1_smul_89543;
  reg [31:0] p1_smul_89544;
  reg [31:0] p1_smul_89545;
  reg [31:0] p1_smul_89546;
  reg [31:0] p1_smul_89965;
  reg [31:0] p1_smul_89966;
  reg [31:0] p1_smul_89967;
  reg [31:0] p1_smul_89968;
  reg [31:0] p1_smul_89969;
  reg [31:0] p1_smul_89970;
  reg [31:0] p1_smul_89547;
  reg [31:0] p1_smul_89548;
  reg [31:0] p1_smul_89549;
  reg [31:0] p1_smul_89550;
  reg [31:0] p1_smul_89971;
  reg [31:0] p1_smul_89972;
  reg [31:0] p1_smul_89973;
  reg [31:0] p1_smul_89974;
  reg [31:0] p1_smul_89975;
  reg [31:0] p1_smul_89976;
  reg [31:0] p1_smul_89551;
  reg [31:0] p1_smul_89552;
  reg [31:0] p1_smul_89553;
  reg [31:0] p1_smul_89554;
  reg [31:0] p1_smul_89977;
  reg [31:0] p1_smul_89978;
  reg [31:0] p1_smul_89979;
  reg [31:0] p1_smul_89980;
  reg [31:0] p1_smul_89981;
  reg [31:0] p1_smul_89982;
  reg [31:0] p1_smul_89555;
  reg [31:0] p1_smul_89556;
  reg [31:0] p1_smul_89557;
  reg [31:0] p1_smul_89558;
  reg [31:0] p1_smul_89983;
  reg [31:0] p1_smul_89984;
  reg [31:0] p1_smul_89985;
  reg [31:0] p1_smul_89986;
  reg [31:0] p1_smul_89987;
  reg [31:0] p1_smul_89988;
  reg [31:0] p1_smul_89559;
  reg [31:0] p1_smul_89560;
  reg [31:0] p1_smul_89561;
  reg [31:0] p1_smul_89562;
  reg [31:0] p1_smul_89989;
  reg [31:0] p1_smul_89990;
  reg [31:0] p1_smul_89991;
  reg [31:0] p1_smul_89992;
  reg [31:0] p1_smul_89993;
  reg [31:0] p1_smul_89994;
  reg [31:0] p1_smul_89563;
  reg [31:0] p1_smul_89564;
  reg [31:0] p1_smul_89565;
  reg [31:0] p1_smul_89566;
  reg [31:0] p1_smul_89995;
  reg [31:0] p1_smul_89996;
  reg [31:0] p1_smul_89997;
  reg [31:0] p1_smul_89998;
  reg [31:0] p1_smul_89999;
  reg [31:0] p1_smul_90000;
  reg [31:0] p1_smul_89567;
  reg [31:0] p1_smul_89568;
  reg [31:0] p1_smul_89569;
  reg [31:0] p1_smul_89570;
  reg [31:0] p1_smul_90001;
  reg [31:0] p1_smul_90002;
  reg [31:0] p1_smul_90003;
  reg [31:0] p1_smul_90004;
  reg [31:0] p1_smul_90005;
  reg [31:0] p1_smul_90006;
  reg [31:0] p1_smul_89571;
  reg [31:0] p1_smul_89572;
  reg [31:0] p1_smul_89573;
  reg [31:0] p1_smul_89574;
  reg [31:0] p1_smul_90007;
  reg [31:0] p1_smul_90008;
  reg [31:0] p1_smul_90009;
  reg [31:0] p1_smul_90010;
  reg [31:0] p1_smul_90011;
  reg [31:0] p1_smul_90012;
  reg [31:0] p1_smul_89575;
  reg [31:0] p1_smul_89576;
  reg [31:0] p1_smul_89577;
  reg [31:0] p1_smul_89578;
  reg [31:0] p1_smul_90013;
  reg [31:0] p1_smul_90014;
  reg [31:0] p1_smul_90015;
  reg [31:0] p1_smul_90016;
  reg [31:0] p1_smul_90017;
  reg [31:0] p1_smul_90018;
  reg [31:0] p1_smul_89579;
  reg [31:0] p1_smul_89580;
  reg [31:0] p1_smul_89581;
  reg [31:0] p1_smul_89582;
  reg [31:0] p1_smul_90019;
  reg [31:0] p1_smul_90020;
  reg [31:0] p1_smul_90021;
  reg [31:0] p1_smul_90022;
  reg [31:0] p1_smul_90023;
  reg [31:0] p1_smul_90024;
  reg [31:0] p1_smul_89583;
  reg [31:0] p1_smul_89584;
  reg [31:0] p1_smul_89585;
  reg [31:0] p1_smul_89586;
  reg [31:0] p1_smul_90025;
  reg [31:0] p1_smul_90026;
  reg [31:0] p1_smul_90027;
  reg [31:0] p1_smul_90028;
  reg [31:0] p1_smul_90029;
  reg [31:0] p1_smul_90030;
  reg [31:0] p1_smul_89587;
  reg [31:0] p1_smul_89588;
  reg [31:0] p1_smul_89589;
  reg [31:0] p1_smul_89590;
  reg [31:0] p1_smul_90031;
  reg [31:0] p1_smul_90032;
  reg [31:0] p1_smul_90033;
  reg [31:0] p1_smul_90034;
  reg [31:0] p1_smul_90035;
  reg [31:0] p1_smul_90036;
  reg [31:0] p1_smul_89591;
  reg [31:0] p1_smul_89592;
  reg [31:0] p1_smul_89593;
  reg [31:0] p1_smul_89594;
  reg [31:0] p1_smul_90037;
  reg [31:0] p1_smul_90038;
  reg [31:0] p1_smul_90039;
  reg [31:0] p1_smul_90040;
  reg [31:0] p1_smul_90041;
  reg [31:0] p1_smul_90042;
  reg [31:0] p1_smul_89595;
  reg [31:0] p1_smul_89596;
  reg [31:0] p1_smul_89597;
  reg [31:0] p1_smul_89598;
  reg [31:0] p1_smul_90043;
  reg [31:0] p1_smul_90044;
  reg [31:0] p1_smul_90045;
  reg [31:0] p1_smul_90046;
  reg [31:0] p1_smul_90047;
  reg [31:0] p1_smul_90048;
  reg [31:0] p1_smul_89599;
  reg [31:0] p1_smul_89600;
  reg [31:0] p1_smul_89601;
  reg [31:0] p1_smul_89602;
  reg [31:0] p1_smul_90049;
  reg [31:0] p1_smul_90050;
  reg [31:0] p1_smul_90051;
  reg [31:0] p1_smul_90052;
  reg [31:0] p1_smul_90053;
  reg [31:0] p1_smul_90054;
  reg [31:0] p1_smul_89603;
  reg [31:0] p1_smul_89604;
  reg [31:0] p1_smul_89605;
  reg [31:0] p1_smul_89606;
  reg [31:0] p1_smul_90055;
  reg [31:0] p1_smul_90056;
  reg [31:0] p1_smul_90057;
  reg [31:0] p1_smul_90058;
  reg [31:0] p1_smul_90059;
  reg [31:0] p1_smul_90060;
  reg [31:0] p1_smul_89607;
  reg [31:0] p1_smul_89608;
  reg [31:0] p1_smul_89609;
  reg [31:0] p1_smul_89610;
  reg [31:0] p1_smul_90061;
  reg [31:0] p1_smul_90062;
  reg [31:0] p1_smul_90063;
  reg [31:0] p1_smul_90064;
  reg [31:0] p1_smul_90065;
  reg [31:0] p1_smul_90066;
  reg [31:0] p1_smul_89611;
  reg [31:0] p1_smul_89612;
  reg [31:0] p1_smul_89613;
  reg [31:0] p1_smul_89614;
  reg [31:0] p1_smul_90067;
  reg [31:0] p1_smul_90068;
  reg [31:0] p1_smul_90069;
  reg [31:0] p1_smul_90070;
  reg [31:0] p1_smul_90071;
  reg [31:0] p1_smul_90072;
  reg [31:0] p1_smul_89615;
  reg [31:0] p1_smul_89616;
  reg [31:0] p1_smul_89617;
  reg [31:0] p1_smul_89618;
  reg [31:0] p1_smul_90073;
  reg [31:0] p1_smul_90074;
  reg [31:0] p1_smul_90075;
  reg [31:0] p1_smul_90076;
  reg [31:0] p1_smul_90077;
  reg [31:0] p1_smul_90078;
  reg [31:0] p1_smul_89619;
  reg [31:0] p1_smul_89620;
  reg [31:0] p1_smul_89621;
  reg [31:0] p1_smul_89622;
  reg [31:0] p1_smul_90079;
  reg [31:0] p1_smul_90080;
  reg [31:0] p1_smul_90081;
  reg [31:0] p1_smul_90082;
  reg [31:0] p1_smul_90083;
  reg [31:0] p1_smul_90084;
  reg [31:0] p1_smul_89623;
  reg [31:0] p1_smul_89624;
  reg [31:0] p1_smul_89625;
  reg [31:0] p1_smul_89626;
  reg [31:0] p1_smul_90085;
  reg [31:0] p1_smul_90086;
  reg [31:0] p1_smul_90087;
  reg [31:0] p1_smul_90088;
  reg [31:0] p1_smul_90089;
  reg [31:0] p1_smul_90090;
  reg [31:0] p1_smul_89627;
  reg [31:0] p1_smul_89628;
  reg [31:0] p1_smul_89629;
  reg [31:0] p1_smul_89630;
  reg [31:0] p1_smul_90091;
  reg [31:0] p1_smul_90092;
  reg [31:0] p1_smul_90093;
  reg [31:0] p1_smul_90094;
  reg [31:0] p1_smul_90095;
  reg [31:0] p1_smul_90096;
  reg [31:0] p1_smul_89631;
  reg [31:0] p1_smul_89632;
  reg [31:0] p1_smul_89633;
  reg [31:0] p1_smul_89634;
  reg [31:0] p1_smul_90097;
  reg [31:0] p1_smul_90098;
  reg [31:0] p1_smul_90099;
  reg [31:0] p1_smul_90100;
  reg [31:0] p1_smul_90101;
  reg [31:0] p1_smul_90102;
  reg [31:0] p1_smul_89635;
  reg [31:0] p1_smul_89636;
  reg [31:0] p1_smul_89637;
  reg [31:0] p1_smul_89638;
  reg [31:0] p1_smul_90103;
  reg [31:0] p1_smul_90104;
  reg [31:0] p1_smul_90105;
  reg [31:0] p1_smul_90106;
  reg [31:0] p1_smul_90107;
  reg [31:0] p1_smul_90108;
  reg [31:0] p1_smul_89639;
  reg [31:0] p1_smul_89640;
  reg [31:0] p1_smul_89641;
  reg [31:0] p1_smul_89642;
  reg [31:0] p1_smul_90109;
  reg [31:0] p1_smul_90110;
  reg [31:0] p1_smul_90111;
  reg [31:0] p1_smul_90112;
  reg [31:0] p1_smul_90113;
  reg [31:0] p1_smul_90114;
  reg [31:0] p1_smul_89643;
  reg [31:0] p1_smul_89644;
  reg [31:0] p1_smul_89645;
  reg [31:0] p1_smul_89646;
  reg [31:0] p1_smul_90115;
  reg [31:0] p1_smul_90116;
  reg [31:0] p1_smul_90117;
  reg [31:0] p1_smul_90118;
  reg [31:0] p1_smul_90119;
  reg [31:0] p1_smul_90120;
  reg [31:0] p1_smul_89647;
  reg [31:0] p1_smul_89648;
  reg [31:0] p1_smul_89649;
  reg [31:0] p1_smul_89650;
  reg [31:0] p1_smul_90121;
  reg [31:0] p1_smul_90122;
  reg [31:0] p1_smul_90123;
  reg [31:0] p1_smul_90124;
  reg [31:0] p1_smul_90125;
  reg [31:0] p1_smul_90126;
  reg [31:0] p1_smul_89651;
  reg [31:0] p1_smul_89652;
  reg [31:0] p1_smul_89653;
  reg [31:0] p1_smul_89654;
  reg [31:0] p1_smul_90127;
  reg [31:0] p1_smul_90128;
  reg [31:0] p1_smul_90129;
  reg [31:0] p1_smul_90130;
  reg [31:0] p1_smul_90131;
  reg [31:0] p1_smul_90132;
  reg [31:0] p1_smul_89655;
  reg [31:0] p1_smul_89656;
  reg [31:0] p1_smul_89657;
  reg [31:0] p1_smul_89658;
  reg [31:0] p1_smul_90133;
  reg [31:0] p1_smul_90134;
  reg [31:0] p1_smul_90135;
  reg [31:0] p1_smul_90136;
  reg [31:0] p1_smul_90137;
  reg [31:0] p1_smul_90138;
  reg [31:0] p1_smul_89659;
  reg [31:0] p1_smul_89660;
  reg [31:0] p1_smul_89661;
  reg [31:0] p1_smul_89662;
  reg [31:0] p1_smul_90139;
  reg [31:0] p1_smul_90140;
  reg [31:0] p1_smul_90141;
  reg [31:0] p1_smul_90142;
  reg [31:0] p1_smul_90143;
  reg [31:0] p1_smul_90144;
  reg [31:0] p1_smul_89663;
  reg [31:0] p1_smul_89664;
  reg [31:0] p1_smul_89665;
  reg [31:0] p1_smul_89666;
  reg [31:0] p1_smul_90145;
  reg [31:0] p1_smul_90146;
  reg [31:0] p1_smul_90147;
  reg [31:0] p1_smul_90148;
  reg [31:0] p1_smul_90149;
  reg [31:0] p1_smul_90150;
  reg [31:0] p1_smul_89667;
  reg [31:0] p1_smul_89668;
  reg [31:0] p1_smul_89669;
  reg [31:0] p1_smul_89670;
  reg [31:0] p1_smul_90151;
  reg [31:0] p1_smul_90152;
  reg [31:0] p1_smul_90153;
  reg [31:0] p1_smul_90154;
  reg [31:0] p1_smul_90155;
  reg [31:0] p1_smul_90156;
  reg [31:0] p1_smul_89671;
  reg [31:0] p1_smul_89672;
  reg [31:0] p1_smul_89673;
  reg [31:0] p1_smul_89674;
  reg [31:0] p1_smul_90157;
  reg [31:0] p1_smul_90158;
  reg [31:0] p1_smul_90159;
  reg [31:0] p1_smul_90160;
  reg [31:0] p1_smul_90161;
  reg [31:0] p1_smul_90162;
  reg [31:0] p1_smul_89675;
  reg [31:0] p1_smul_89676;
  reg [31:0] p1_smul_89677;
  reg [31:0] p1_smul_89678;
  reg [31:0] p1_smul_90163;
  reg [31:0] p1_smul_90164;
  reg [31:0] p1_smul_90165;
  reg [31:0] p1_smul_90166;
  reg [31:0] p1_smul_90167;
  reg [31:0] p1_smul_90168;
  reg [31:0] p1_smul_89679;
  reg [31:0] p1_smul_89680;
  reg [31:0] p1_smul_89681;
  reg [31:0] p1_smul_89682;
  reg [31:0] p1_smul_90169;
  reg [31:0] p1_smul_90170;
  reg [31:0] p1_smul_90171;
  reg [31:0] p1_smul_90172;
  reg [31:0] p1_smul_90173;
  reg [31:0] p1_smul_90174;
  reg [31:0] p1_smul_89683;
  reg [31:0] p1_smul_89684;
  reg [31:0] p1_smul_89685;
  reg [31:0] p1_smul_89686;
  reg [31:0] p1_smul_90175;
  reg [31:0] p1_smul_90176;
  reg [31:0] p1_smul_90177;
  reg [31:0] p1_smul_90178;
  reg [31:0] p1_smul_90179;
  reg [31:0] p1_smul_90180;
  reg [31:0] p1_smul_89687;
  reg [31:0] p1_smul_89688;
  reg [31:0] p1_smul_89689;
  reg [31:0] p1_smul_89690;
  reg [31:0] p1_smul_90181;
  reg [31:0] p1_smul_90182;
  reg [31:0] p1_smul_90183;
  reg [31:0] p1_smul_90184;
  reg [31:0] p1_smul_90185;
  reg [31:0] p1_smul_90186;
  reg [31:0] p1_smul_89691;
  reg [31:0] p1_smul_89692;
  reg [31:0] p1_smul_89693;
  reg [31:0] p1_smul_89694;
  reg [31:0] p1_smul_90187;
  reg [31:0] p1_smul_90188;
  reg [31:0] p1_smul_90189;
  reg [31:0] p1_smul_90190;
  reg [31:0] p1_smul_90191;
  reg [31:0] p1_smul_90192;
  reg [31:0] p1_smul_89695;
  reg [31:0] p1_smul_89696;
  reg [31:0] p1_smul_89697;
  reg [31:0] p1_smul_89698;
  reg [31:0] p1_smul_90193;
  reg [31:0] p1_smul_90194;
  reg [31:0] p1_smul_90195;
  reg [31:0] p1_smul_90196;
  reg [31:0] p1_smul_90197;
  reg [31:0] p1_smul_90198;
  reg [31:0] p1_smul_89699;
  reg [31:0] p1_smul_89700;
  reg [31:0] p1_smul_89701;
  reg [31:0] p1_smul_89702;
  reg [31:0] p1_smul_90199;
  reg [31:0] p1_smul_90200;
  reg [31:0] p1_smul_90201;
  reg [31:0] p1_smul_90202;
  reg [31:0] p1_smul_90203;
  reg [31:0] p1_smul_90204;
  reg [31:0] p1_smul_89703;
  reg [31:0] p1_smul_89704;
  reg [31:0] p1_smul_89705;
  reg [31:0] p1_smul_89706;
  reg [31:0] p1_smul_90205;
  reg [31:0] p1_smul_90206;
  reg [31:0] p1_smul_90207;
  reg [31:0] p1_smul_90208;
  reg [31:0] p1_smul_90209;
  reg [31:0] p1_smul_90210;
  reg [31:0] p1_smul_89707;
  reg [31:0] p1_smul_89708;
  reg [31:0] p1_smul_89709;
  reg [31:0] p1_smul_89710;
  reg [31:0] p1_smul_90211;
  reg [31:0] p1_smul_90212;
  reg [31:0] p1_smul_90213;
  reg [31:0] p1_smul_90214;
  reg [31:0] p1_smul_90215;
  reg [31:0] p1_smul_90216;
  reg [31:0] p1_smul_89711;
  reg [31:0] p1_smul_89712;
  reg [31:0] p1_smul_89713;
  reg [31:0] p1_smul_89714;
  reg [31:0] p1_smul_90217;
  reg [31:0] p1_smul_90218;
  reg [31:0] p1_smul_90219;
  reg [31:0] p1_smul_90220;
  reg [31:0] p1_smul_90221;
  reg [31:0] p1_smul_90222;
  reg [31:0] p1_smul_89715;
  reg [31:0] p1_smul_89716;
  reg [31:0] p1_smul_89717;
  reg [31:0] p1_smul_89718;
  reg [31:0] p1_smul_90223;
  reg [31:0] p1_smul_90224;
  reg [31:0] p1_smul_90225;
  reg [31:0] p1_smul_90226;
  reg [31:0] p1_smul_90227;
  reg [31:0] p1_smul_90228;
  reg [31:0] p1_smul_89719;
  reg [31:0] p1_smul_89720;
  reg [31:0] p1_smul_89721;
  reg [31:0] p1_smul_89722;
  reg [31:0] p1_smul_90229;
  reg [31:0] p1_smul_90230;
  reg [31:0] p1_smul_90231;
  reg [31:0] p1_smul_90232;
  reg [31:0] p1_smul_90233;
  reg [31:0] p1_smul_90234;
  reg [31:0] p1_smul_89723;
  reg [31:0] p1_smul_89724;
  reg [31:0] p1_smul_89725;
  reg [31:0] p1_smul_89726;
  reg [31:0] p1_smul_90235;
  reg [31:0] p1_smul_90236;
  reg [31:0] p1_smul_90237;
  reg [31:0] p1_smul_90238;
  reg [31:0] p1_smul_90239;
  reg [31:0] p1_smul_90240;
  reg [31:0] p1_smul_89727;
  reg [31:0] p1_smul_89728;
  reg [31:0] p1_smul_89729;
  reg [31:0] p1_smul_89730;
  reg [31:0] p1_smul_90241;
  reg [31:0] p1_smul_90242;
  reg [31:0] p1_smul_90243;
  reg [31:0] p1_smul_90244;
  reg [31:0] p1_smul_90245;
  reg [31:0] p1_smul_90246;
  reg [31:0] p1_smul_89731;
  reg [31:0] p1_smul_89732;
  reg [31:0] p1_smul_89733;
  reg [31:0] p1_smul_89734;
  reg [31:0] p1_smul_90247;
  reg [31:0] p1_smul_90248;
  reg [31:0] p1_smul_90249;
  reg [31:0] p1_smul_90250;
  reg [31:0] p1_smul_90251;
  reg [31:0] p1_smul_90252;
  reg [31:0] p1_smul_89735;
  reg [31:0] p1_smul_89736;
  reg [31:0] p1_smul_89737;
  reg [31:0] p1_smul_89738;
  reg [31:0] p1_smul_90253;
  reg [31:0] p1_smul_90254;
  reg [31:0] p1_smul_90255;
  reg [31:0] p1_smul_90256;
  reg [31:0] p1_smul_90257;
  reg [31:0] p1_smul_90258;
  reg [31:0] p1_smul_89739;
  reg [31:0] p1_smul_89740;
  reg [31:0] p1_smul_89741;
  reg [31:0] p1_smul_89742;
  reg [31:0] p1_smul_90259;
  reg [31:0] p1_smul_90260;
  reg [31:0] p1_smul_90261;
  reg [31:0] p1_smul_90262;
  reg [31:0] p1_smul_90263;
  reg [31:0] p1_smul_90264;
  reg [31:0] p1_smul_89743;
  reg [31:0] p1_smul_89744;
  reg [31:0] p1_smul_89745;
  reg [31:0] p1_smul_89746;
  reg [31:0] p1_smul_90265;
  reg [31:0] p1_smul_90266;
  reg [31:0] p1_smul_90267;
  reg [31:0] p1_smul_90268;
  reg [31:0] p1_smul_90269;
  reg [31:0] p1_smul_90270;
  reg [31:0] p1_smul_89747;
  reg [31:0] p1_smul_89748;
  reg [31:0] p1_smul_89749;
  reg [31:0] p1_smul_89750;
  reg [31:0] p1_smul_90271;
  reg [31:0] p1_smul_90272;
  reg [31:0] p1_smul_90273;
  reg [31:0] p1_smul_90274;
  reg [31:0] p1_smul_90275;
  reg [31:0] p1_smul_90276;
  reg [31:0] p1_smul_89751;
  reg [31:0] p1_smul_89752;
  reg [31:0] p1_smul_89753;
  reg [31:0] p1_smul_89754;
  reg [31:0] p1_smul_90277;
  reg [31:0] p1_smul_90278;
  reg [31:0] p1_smul_90279;
  reg [31:0] p1_smul_90280;
  reg [31:0] p1_smul_90281;
  reg [31:0] p1_smul_90282;
  reg [31:0] p1_smul_89755;
  reg [31:0] p1_smul_89756;
  reg [31:0] p1_smul_89757;
  reg [31:0] p1_smul_89758;
  reg [31:0] p1_smul_90283;
  reg [31:0] p1_smul_90284;
  reg [31:0] p1_smul_90285;
  reg [31:0] p1_smul_90286;
  reg [31:0] p1_smul_90287;
  reg [31:0] p1_smul_90288;
  reg [31:0] p1_smul_89759;
  reg [31:0] p1_smul_89760;
  reg [31:0] p1_smul_89761;
  reg [31:0] p1_smul_89762;
  reg [31:0] p1_smul_90289;
  reg [31:0] p1_smul_90290;
  reg [31:0] p1_smul_90291;
  reg [31:0] p1_smul_90292;
  reg [31:0] p1_smul_90293;
  reg [31:0] p1_smul_90294;
  reg [31:0] p1_smul_89763;
  reg [31:0] p1_smul_89764;
  reg [31:0] p1_smul_89765;
  reg [31:0] p1_smul_89766;
  reg [31:0] p1_smul_90295;
  reg [31:0] p1_smul_90296;
  reg [31:0] p1_smul_90297;
  reg [31:0] p1_smul_90298;
  reg [31:0] p1_smul_90299;
  reg [31:0] p1_smul_90300;
  reg [31:0] p1_smul_89767;
  reg [31:0] p1_smul_89768;
  reg [31:0] p1_smul_89769;
  reg [31:0] p1_smul_89770;
  reg [31:0] p1_smul_90301;
  reg [31:0] p1_smul_90302;
  reg [31:0] p1_smul_90303;
  reg [31:0] p1_smul_90304;
  reg [31:0] p1_smul_90305;
  reg [31:0] p1_smul_90306;
  reg [31:0] p1_smul_89771;
  reg [31:0] p1_smul_89772;
  reg [31:0] p1_smul_89773;
  reg [31:0] p1_smul_89774;
  reg [31:0] p1_smul_90307;
  reg [31:0] p1_smul_90308;
  reg [31:0] p1_smul_90309;
  reg [31:0] p1_smul_90310;
  reg [31:0] p1_smul_90311;
  reg [31:0] p1_smul_90312;
  reg [31:0] p1_smul_89775;
  reg [31:0] p1_smul_89776;
  reg [31:0] p1_smul_89777;
  reg [31:0] p1_smul_89778;
  reg [31:0] p1_smul_90313;
  reg [31:0] p1_smul_90314;
  reg [31:0] p1_smul_90315;
  reg [31:0] p1_smul_90316;
  reg [31:0] p1_smul_90317;
  reg [31:0] p1_smul_90318;
  reg [31:0] p1_smul_89779;
  reg [31:0] p1_smul_89780;
  reg [31:0] p1_smul_89781;
  reg [31:0] p1_smul_89782;
  reg [31:0] p1_smul_90319;
  reg [31:0] p1_smul_90320;
  reg [31:0] p1_smul_90321;
  reg [31:0] p1_smul_90322;
  reg [31:0] p1_smul_90323;
  reg [31:0] p1_smul_90324;
  reg [31:0] p1_smul_89783;
  reg [31:0] p1_smul_89784;
  reg [31:0] p1_smul_89785;
  reg [31:0] p1_smul_89786;
  reg [31:0] p1_smul_90325;
  reg [31:0] p1_smul_90326;
  reg [31:0] p1_smul_90327;
  reg [31:0] p1_smul_90328;
  reg [31:0] p1_smul_90329;
  reg [31:0] p1_smul_90330;
  reg [31:0] p1_smul_89787;
  reg [31:0] p1_smul_89788;
  reg [31:0] p1_smul_89789;
  reg [31:0] p1_smul_89790;
  reg [31:0] p1_smul_90331;
  reg [31:0] p1_smul_90332;
  reg [31:0] p1_smul_90333;
  reg [31:0] p1_smul_90334;
  reg [31:0] p1_smul_90335;
  reg [31:0] p1_smul_90336;
  reg [31:0] p1_smul_89791;
  reg [31:0] p1_smul_89792;
  reg [31:0] p1_smul_89793;
  reg [31:0] p1_smul_89794;
  reg [31:0] p1_smul_90337;
  reg [31:0] p1_smul_90338;
  reg [31:0] p1_smul_90339;
  reg [31:0] p1_smul_90340;
  reg [31:0] p1_smul_90341;
  reg [31:0] p1_smul_90342;
  reg [31:0] p1_smul_89795;
  reg [31:0] p1_smul_89796;
  reg [31:0] p1_smul_89797;
  reg [31:0] p1_smul_89798;
  reg [31:0] p1_smul_90343;
  reg [31:0] p1_smul_90344;
  reg [31:0] p1_smul_90345;
  reg [31:0] p1_smul_90346;
  reg [31:0] p1_smul_90347;
  reg [31:0] p1_smul_90348;
  reg [31:0] p1_smul_89799;
  reg [31:0] p1_smul_89800;
  reg [31:0] p1_smul_89801;
  reg [31:0] p1_smul_89802;
  reg [31:0] p1_smul_90349;
  reg [31:0] p1_smul_90350;
  reg [31:0] p1_smul_90351;
  reg [31:0] p1_smul_90352;
  reg [31:0] p1_smul_90353;
  reg [31:0] p1_smul_90354;
  reg [31:0] p1_smul_89803;
  reg [31:0] p1_smul_89804;
  reg [31:0] p1_smul_89805;
  reg [31:0] p1_smul_89806;
  reg [31:0] p1_smul_90355;
  reg [31:0] p1_smul_90356;
  reg [31:0] p1_smul_90357;
  reg [31:0] p1_smul_90358;
  reg [31:0] p1_smul_90359;
  reg [31:0] p1_smul_90360;
  reg [31:0] p1_smul_89807;
  reg [31:0] p1_smul_89808;
  reg [31:0] p1_smul_89809;
  reg [31:0] p1_smul_89810;
  reg [31:0] p1_smul_90361;
  reg [31:0] p1_smul_90362;
  reg [31:0] p1_smul_90363;
  reg [31:0] p1_smul_90364;
  reg [31:0] p1_smul_90365;
  reg [31:0] p1_smul_90366;
  reg [31:0] p1_smul_89811;
  reg [31:0] p1_smul_89812;
  reg [31:0] p1_smul_89813;
  reg [31:0] p1_smul_89814;
  reg [31:0] p1_smul_90367;
  reg [31:0] p1_smul_90368;
  reg [31:0] p1_smul_90369;
  reg [31:0] p1_smul_90370;
  reg [31:0] p1_smul_90371;
  reg [31:0] p1_smul_90372;
  reg [31:0] p1_smul_89815;
  reg [31:0] p1_smul_89816;
  reg [31:0] p1_smul_89817;
  reg [31:0] p1_smul_89818;
  reg [31:0] p1_smul_90373;
  reg [31:0] p1_smul_90374;
  reg [31:0] p1_smul_90375;
  reg [31:0] p1_smul_90376;
  reg [31:0] p1_smul_90377;
  reg [31:0] p1_smul_90378;
  reg [31:0] p1_smul_89819;
  reg [31:0] p1_smul_89820;
  reg [31:0] p1_smul_89821;
  reg [31:0] p1_smul_89822;
  reg [31:0] p1_smul_90379;
  reg [31:0] p1_smul_90380;
  reg [31:0] p1_smul_90381;
  reg [31:0] p1_smul_90382;
  reg [31:0] p1_smul_90383;
  reg [31:0] p1_smul_90384;
  reg [31:0] p1_smul_89823;
  reg [31:0] p1_smul_89824;
  reg [31:0] p1_smul_89825;
  reg [31:0] p1_smul_89826;
  reg [31:0] p1_smul_90385;
  reg [31:0] p1_smul_90386;
  reg [31:0] p1_smul_90387;
  reg [31:0] p1_smul_90388;
  reg [31:0] p1_smul_90389;
  reg [31:0] p1_smul_90390;
  reg [31:0] p1_smul_89827;
  reg [31:0] p1_smul_89828;
  reg [31:0] p1_smul_89829;
  reg [31:0] p1_smul_89830;
  reg [31:0] p1_smul_90391;
  reg [31:0] p1_smul_90392;
  reg [31:0] p1_smul_90393;
  reg [31:0] p1_smul_90394;
  reg [31:0] p1_smul_90395;
  reg [31:0] p1_smul_90396;
  reg [31:0] p1_smul_89831;
  reg [31:0] p1_smul_89832;
  reg [31:0] p1_smul_89833;
  reg [31:0] p1_smul_89834;
  reg [31:0] p1_smul_90397;
  reg [31:0] p1_smul_90398;
  reg [31:0] p1_smul_90399;
  reg [31:0] p1_smul_90400;
  reg [31:0] p1_smul_90401;
  reg [31:0] p1_smul_90402;
  reg [31:0] p1_smul_89835;
  reg [31:0] p1_smul_89836;
  reg [31:0] p1_smul_89837;
  reg [31:0] p1_smul_89838;
  reg [31:0] p1_smul_90403;
  reg [31:0] p1_smul_90404;
  reg [31:0] p1_smul_90405;
  reg [31:0] p1_smul_90406;
  reg [31:0] p1_smul_90407;
  reg [31:0] p1_smul_90408;
  reg [31:0] p1_smul_89839;
  reg [31:0] p1_smul_89840;
  reg [31:0] p1_smul_89841;
  reg [31:0] p1_smul_89842;
  reg [31:0] p1_smul_90409;
  reg [31:0] p1_smul_90410;
  reg [31:0] p1_smul_90411;
  reg [31:0] p1_smul_90412;
  reg [31:0] p1_smul_90413;
  reg [31:0] p1_smul_90414;
  reg [31:0] p1_smul_89843;
  reg [31:0] p1_smul_89844;
  reg [31:0] p1_smul_89845;
  reg [31:0] p1_smul_89846;
  reg [31:0] p1_smul_90415;
  reg [31:0] p1_smul_90416;
  reg [31:0] p1_smul_90417;
  reg [31:0] p1_smul_90418;
  reg [31:0] p1_smul_90419;
  reg [31:0] p1_smul_90420;
  reg [31:0] p1_smul_89847;
  reg [31:0] p1_smul_89848;
  reg [31:0] p1_smul_89849;
  reg [31:0] p1_smul_89850;
  reg [31:0] p1_smul_90421;
  reg [31:0] p1_smul_90422;
  reg [31:0] p1_smul_90423;
  reg [31:0] p1_smul_90424;
  reg [31:0] p1_smul_90425;
  reg [31:0] p1_smul_90426;
  reg [31:0] p1_smul_89851;
  reg [31:0] p1_smul_89852;
  reg [31:0] p1_smul_89853;
  reg [31:0] p1_smul_89854;
  reg [31:0] p1_smul_90427;
  reg [31:0] p1_smul_90428;
  reg [31:0] p1_smul_90429;
  reg [31:0] p1_smul_90430;
  reg [31:0] p1_smul_90431;
  reg [31:0] p1_smul_90432;
  reg [31:0] p1_smul_89855;
  reg [31:0] p1_smul_89856;
  reg [31:0] p1_smul_89857;
  reg [31:0] p1_smul_89858;
  reg [31:0] p1_smul_90433;
  reg [31:0] p1_smul_90434;
  reg [31:0] p1_smul_90435;
  reg [31:0] p1_smul_90436;
  reg [31:0] p1_smul_90437;
  reg [31:0] p1_smul_90438;
  reg [31:0] p1_smul_89859;
  reg [31:0] p1_smul_89860;
  reg [31:0] p1_smul_89861;
  reg [31:0] p1_smul_89862;
  reg [31:0] p1_smul_90439;
  reg [31:0] p1_smul_90440;
  reg [31:0] p1_smul_90441;
  reg [31:0] p1_smul_90442;
  reg [31:0] p1_smul_90443;
  reg [31:0] p1_smul_90444;
  reg [31:0] p1_smul_89863;
  reg [31:0] p1_smul_89864;
  reg [31:0] p1_smul_89865;
  reg [31:0] p1_smul_89866;
  reg [31:0] p1_smul_90445;
  reg [31:0] p1_smul_90446;
  reg [31:0] p1_smul_90447;
  reg [31:0] p1_smul_90448;
  reg [31:0] p1_smul_90449;
  reg [31:0] p1_smul_90450;
  reg [31:0] p1_smul_89867;
  reg [31:0] p1_smul_89868;
  reg [31:0] p1_smul_89869;
  reg [31:0] p1_smul_89870;
  reg [31:0] p1_smul_90451;
  reg [31:0] p1_smul_90452;
  reg [31:0] p1_smul_90453;
  reg [31:0] p1_smul_90454;
  reg [31:0] p1_smul_90455;
  reg [31:0] p1_smul_90456;
  reg [31:0] p1_smul_89871;
  reg [31:0] p1_smul_89872;
  reg [31:0] p1_smul_89873;
  reg [31:0] p1_smul_89874;
  reg [31:0] p1_smul_90457;
  reg [31:0] p1_smul_90458;
  reg [31:0] p1_smul_90459;
  reg [31:0] p1_smul_90460;
  reg [31:0] p1_smul_90461;
  reg [31:0] p1_smul_90462;
  reg [31:0] p1_smul_89875;
  reg [31:0] p1_smul_89876;
  reg [31:0] p1_smul_89877;
  reg [31:0] p1_smul_89878;
  reg [31:0] p1_smul_90463;
  reg [31:0] p1_smul_90464;
  reg [31:0] p1_smul_90465;
  reg [31:0] p1_smul_90466;
  reg [31:0] p1_smul_90467;
  reg [31:0] p1_smul_90468;
  reg [31:0] p1_smul_89879;
  reg [31:0] p1_smul_89880;
  reg [31:0] p1_smul_89881;
  reg [31:0] p1_smul_89882;
  reg [31:0] p1_smul_90469;
  reg [31:0] p1_smul_90470;
  reg [31:0] p1_smul_90471;
  reg [31:0] p1_smul_90472;
  reg [31:0] p1_smul_90473;
  reg [31:0] p1_smul_90474;
  reg [31:0] p1_smul_89883;
  reg [31:0] p1_smul_89884;
  reg [31:0] p1_smul_89885;
  reg [31:0] p1_smul_89886;
  reg [31:0] p1_smul_90475;
  reg [31:0] p1_smul_90476;
  reg [31:0] p1_smul_90477;
  reg [31:0] p1_smul_90478;
  reg [31:0] p1_smul_90479;
  reg [31:0] p1_smul_90480;
  reg [31:0] p1_smul_89887;
  reg [31:0] p1_smul_89888;
  reg [31:0] p1_smul_89889;
  reg [31:0] p1_smul_89890;
  reg [31:0] p1_smul_90481;
  reg [31:0] p1_smul_90482;
  reg [31:0] p1_smul_90483;
  reg [31:0] p1_smul_90484;
  reg [31:0] p1_smul_90485;
  reg [31:0] p1_smul_90486;
  reg [31:0] p1_smul_89891;
  reg [31:0] p1_smul_89892;
  reg [31:0] p1_smul_89893;
  reg [31:0] p1_smul_89894;
  reg [31:0] p1_smul_90487;
  reg [31:0] p1_smul_90488;
  reg [31:0] p1_smul_90489;
  reg [31:0] p1_smul_90490;
  reg [31:0] p1_smul_90491;
  reg [31:0] p1_smul_90492;
  reg [31:0] p1_smul_89895;
  reg [31:0] p1_smul_89896;
  reg [31:0] p1_smul_89897;
  reg [31:0] p1_smul_89898;
  reg [31:0] p1_smul_90493;
  reg [31:0] p1_smul_90494;
  reg [31:0] p1_smul_90495;
  reg [31:0] p1_smul_90496;
  reg [31:0] p1_smul_90497;
  reg [31:0] p1_smul_90498;
  always_ff @ (posedge clk) begin
    p1_smul_89499 <= p1_smul_89499_comb;
    p1_smul_89500 <= p1_smul_89500_comb;
    p1_smul_89501 <= p1_smul_89501_comb;
    p1_smul_89502 <= p1_smul_89502_comb;
    p1_smul_89899 <= p1_smul_89899_comb;
    p1_smul_89900 <= p1_smul_89900_comb;
    p1_smul_89901 <= p1_smul_89901_comb;
    p1_smul_89902 <= p1_smul_89902_comb;
    p1_smul_89903 <= p1_smul_89903_comb;
    p1_smul_89904 <= p1_smul_89904_comb;
    p1_smul_89503 <= p1_smul_89503_comb;
    p1_smul_89504 <= p1_smul_89504_comb;
    p1_smul_89505 <= p1_smul_89505_comb;
    p1_smul_89506 <= p1_smul_89506_comb;
    p1_smul_89905 <= p1_smul_89905_comb;
    p1_smul_89906 <= p1_smul_89906_comb;
    p1_smul_89907 <= p1_smul_89907_comb;
    p1_smul_89908 <= p1_smul_89908_comb;
    p1_smul_89909 <= p1_smul_89909_comb;
    p1_smul_89910 <= p1_smul_89910_comb;
    p1_smul_89507 <= p1_smul_89507_comb;
    p1_smul_89508 <= p1_smul_89508_comb;
    p1_smul_89509 <= p1_smul_89509_comb;
    p1_smul_89510 <= p1_smul_89510_comb;
    p1_smul_89911 <= p1_smul_89911_comb;
    p1_smul_89912 <= p1_smul_89912_comb;
    p1_smul_89913 <= p1_smul_89913_comb;
    p1_smul_89914 <= p1_smul_89914_comb;
    p1_smul_89915 <= p1_smul_89915_comb;
    p1_smul_89916 <= p1_smul_89916_comb;
    p1_smul_89511 <= p1_smul_89511_comb;
    p1_smul_89512 <= p1_smul_89512_comb;
    p1_smul_89513 <= p1_smul_89513_comb;
    p1_smul_89514 <= p1_smul_89514_comb;
    p1_smul_89917 <= p1_smul_89917_comb;
    p1_smul_89918 <= p1_smul_89918_comb;
    p1_smul_89919 <= p1_smul_89919_comb;
    p1_smul_89920 <= p1_smul_89920_comb;
    p1_smul_89921 <= p1_smul_89921_comb;
    p1_smul_89922 <= p1_smul_89922_comb;
    p1_smul_89515 <= p1_smul_89515_comb;
    p1_smul_89516 <= p1_smul_89516_comb;
    p1_smul_89517 <= p1_smul_89517_comb;
    p1_smul_89518 <= p1_smul_89518_comb;
    p1_smul_89923 <= p1_smul_89923_comb;
    p1_smul_89924 <= p1_smul_89924_comb;
    p1_smul_89925 <= p1_smul_89925_comb;
    p1_smul_89926 <= p1_smul_89926_comb;
    p1_smul_89927 <= p1_smul_89927_comb;
    p1_smul_89928 <= p1_smul_89928_comb;
    p1_smul_89519 <= p1_smul_89519_comb;
    p1_smul_89520 <= p1_smul_89520_comb;
    p1_smul_89521 <= p1_smul_89521_comb;
    p1_smul_89522 <= p1_smul_89522_comb;
    p1_smul_89929 <= p1_smul_89929_comb;
    p1_smul_89930 <= p1_smul_89930_comb;
    p1_smul_89931 <= p1_smul_89931_comb;
    p1_smul_89932 <= p1_smul_89932_comb;
    p1_smul_89933 <= p1_smul_89933_comb;
    p1_smul_89934 <= p1_smul_89934_comb;
    p1_smul_89523 <= p1_smul_89523_comb;
    p1_smul_89524 <= p1_smul_89524_comb;
    p1_smul_89525 <= p1_smul_89525_comb;
    p1_smul_89526 <= p1_smul_89526_comb;
    p1_smul_89935 <= p1_smul_89935_comb;
    p1_smul_89936 <= p1_smul_89936_comb;
    p1_smul_89937 <= p1_smul_89937_comb;
    p1_smul_89938 <= p1_smul_89938_comb;
    p1_smul_89939 <= p1_smul_89939_comb;
    p1_smul_89940 <= p1_smul_89940_comb;
    p1_smul_89527 <= p1_smul_89527_comb;
    p1_smul_89528 <= p1_smul_89528_comb;
    p1_smul_89529 <= p1_smul_89529_comb;
    p1_smul_89530 <= p1_smul_89530_comb;
    p1_smul_89941 <= p1_smul_89941_comb;
    p1_smul_89942 <= p1_smul_89942_comb;
    p1_smul_89943 <= p1_smul_89943_comb;
    p1_smul_89944 <= p1_smul_89944_comb;
    p1_smul_89945 <= p1_smul_89945_comb;
    p1_smul_89946 <= p1_smul_89946_comb;
    p1_smul_89531 <= p1_smul_89531_comb;
    p1_smul_89532 <= p1_smul_89532_comb;
    p1_smul_89533 <= p1_smul_89533_comb;
    p1_smul_89534 <= p1_smul_89534_comb;
    p1_smul_89947 <= p1_smul_89947_comb;
    p1_smul_89948 <= p1_smul_89948_comb;
    p1_smul_89949 <= p1_smul_89949_comb;
    p1_smul_89950 <= p1_smul_89950_comb;
    p1_smul_89951 <= p1_smul_89951_comb;
    p1_smul_89952 <= p1_smul_89952_comb;
    p1_smul_89535 <= p1_smul_89535_comb;
    p1_smul_89536 <= p1_smul_89536_comb;
    p1_smul_89537 <= p1_smul_89537_comb;
    p1_smul_89538 <= p1_smul_89538_comb;
    p1_smul_89953 <= p1_smul_89953_comb;
    p1_smul_89954 <= p1_smul_89954_comb;
    p1_smul_89955 <= p1_smul_89955_comb;
    p1_smul_89956 <= p1_smul_89956_comb;
    p1_smul_89957 <= p1_smul_89957_comb;
    p1_smul_89958 <= p1_smul_89958_comb;
    p1_smul_89539 <= p1_smul_89539_comb;
    p1_smul_89540 <= p1_smul_89540_comb;
    p1_smul_89541 <= p1_smul_89541_comb;
    p1_smul_89542 <= p1_smul_89542_comb;
    p1_smul_89959 <= p1_smul_89959_comb;
    p1_smul_89960 <= p1_smul_89960_comb;
    p1_smul_89961 <= p1_smul_89961_comb;
    p1_smul_89962 <= p1_smul_89962_comb;
    p1_smul_89963 <= p1_smul_89963_comb;
    p1_smul_89964 <= p1_smul_89964_comb;
    p1_smul_89543 <= p1_smul_89543_comb;
    p1_smul_89544 <= p1_smul_89544_comb;
    p1_smul_89545 <= p1_smul_89545_comb;
    p1_smul_89546 <= p1_smul_89546_comb;
    p1_smul_89965 <= p1_smul_89965_comb;
    p1_smul_89966 <= p1_smul_89966_comb;
    p1_smul_89967 <= p1_smul_89967_comb;
    p1_smul_89968 <= p1_smul_89968_comb;
    p1_smul_89969 <= p1_smul_89969_comb;
    p1_smul_89970 <= p1_smul_89970_comb;
    p1_smul_89547 <= p1_smul_89547_comb;
    p1_smul_89548 <= p1_smul_89548_comb;
    p1_smul_89549 <= p1_smul_89549_comb;
    p1_smul_89550 <= p1_smul_89550_comb;
    p1_smul_89971 <= p1_smul_89971_comb;
    p1_smul_89972 <= p1_smul_89972_comb;
    p1_smul_89973 <= p1_smul_89973_comb;
    p1_smul_89974 <= p1_smul_89974_comb;
    p1_smul_89975 <= p1_smul_89975_comb;
    p1_smul_89976 <= p1_smul_89976_comb;
    p1_smul_89551 <= p1_smul_89551_comb;
    p1_smul_89552 <= p1_smul_89552_comb;
    p1_smul_89553 <= p1_smul_89553_comb;
    p1_smul_89554 <= p1_smul_89554_comb;
    p1_smul_89977 <= p1_smul_89977_comb;
    p1_smul_89978 <= p1_smul_89978_comb;
    p1_smul_89979 <= p1_smul_89979_comb;
    p1_smul_89980 <= p1_smul_89980_comb;
    p1_smul_89981 <= p1_smul_89981_comb;
    p1_smul_89982 <= p1_smul_89982_comb;
    p1_smul_89555 <= p1_smul_89555_comb;
    p1_smul_89556 <= p1_smul_89556_comb;
    p1_smul_89557 <= p1_smul_89557_comb;
    p1_smul_89558 <= p1_smul_89558_comb;
    p1_smul_89983 <= p1_smul_89983_comb;
    p1_smul_89984 <= p1_smul_89984_comb;
    p1_smul_89985 <= p1_smul_89985_comb;
    p1_smul_89986 <= p1_smul_89986_comb;
    p1_smul_89987 <= p1_smul_89987_comb;
    p1_smul_89988 <= p1_smul_89988_comb;
    p1_smul_89559 <= p1_smul_89559_comb;
    p1_smul_89560 <= p1_smul_89560_comb;
    p1_smul_89561 <= p1_smul_89561_comb;
    p1_smul_89562 <= p1_smul_89562_comb;
    p1_smul_89989 <= p1_smul_89989_comb;
    p1_smul_89990 <= p1_smul_89990_comb;
    p1_smul_89991 <= p1_smul_89991_comb;
    p1_smul_89992 <= p1_smul_89992_comb;
    p1_smul_89993 <= p1_smul_89993_comb;
    p1_smul_89994 <= p1_smul_89994_comb;
    p1_smul_89563 <= p1_smul_89563_comb;
    p1_smul_89564 <= p1_smul_89564_comb;
    p1_smul_89565 <= p1_smul_89565_comb;
    p1_smul_89566 <= p1_smul_89566_comb;
    p1_smul_89995 <= p1_smul_89995_comb;
    p1_smul_89996 <= p1_smul_89996_comb;
    p1_smul_89997 <= p1_smul_89997_comb;
    p1_smul_89998 <= p1_smul_89998_comb;
    p1_smul_89999 <= p1_smul_89999_comb;
    p1_smul_90000 <= p1_smul_90000_comb;
    p1_smul_89567 <= p1_smul_89567_comb;
    p1_smul_89568 <= p1_smul_89568_comb;
    p1_smul_89569 <= p1_smul_89569_comb;
    p1_smul_89570 <= p1_smul_89570_comb;
    p1_smul_90001 <= p1_smul_90001_comb;
    p1_smul_90002 <= p1_smul_90002_comb;
    p1_smul_90003 <= p1_smul_90003_comb;
    p1_smul_90004 <= p1_smul_90004_comb;
    p1_smul_90005 <= p1_smul_90005_comb;
    p1_smul_90006 <= p1_smul_90006_comb;
    p1_smul_89571 <= p1_smul_89571_comb;
    p1_smul_89572 <= p1_smul_89572_comb;
    p1_smul_89573 <= p1_smul_89573_comb;
    p1_smul_89574 <= p1_smul_89574_comb;
    p1_smul_90007 <= p1_smul_90007_comb;
    p1_smul_90008 <= p1_smul_90008_comb;
    p1_smul_90009 <= p1_smul_90009_comb;
    p1_smul_90010 <= p1_smul_90010_comb;
    p1_smul_90011 <= p1_smul_90011_comb;
    p1_smul_90012 <= p1_smul_90012_comb;
    p1_smul_89575 <= p1_smul_89575_comb;
    p1_smul_89576 <= p1_smul_89576_comb;
    p1_smul_89577 <= p1_smul_89577_comb;
    p1_smul_89578 <= p1_smul_89578_comb;
    p1_smul_90013 <= p1_smul_90013_comb;
    p1_smul_90014 <= p1_smul_90014_comb;
    p1_smul_90015 <= p1_smul_90015_comb;
    p1_smul_90016 <= p1_smul_90016_comb;
    p1_smul_90017 <= p1_smul_90017_comb;
    p1_smul_90018 <= p1_smul_90018_comb;
    p1_smul_89579 <= p1_smul_89579_comb;
    p1_smul_89580 <= p1_smul_89580_comb;
    p1_smul_89581 <= p1_smul_89581_comb;
    p1_smul_89582 <= p1_smul_89582_comb;
    p1_smul_90019 <= p1_smul_90019_comb;
    p1_smul_90020 <= p1_smul_90020_comb;
    p1_smul_90021 <= p1_smul_90021_comb;
    p1_smul_90022 <= p1_smul_90022_comb;
    p1_smul_90023 <= p1_smul_90023_comb;
    p1_smul_90024 <= p1_smul_90024_comb;
    p1_smul_89583 <= p1_smul_89583_comb;
    p1_smul_89584 <= p1_smul_89584_comb;
    p1_smul_89585 <= p1_smul_89585_comb;
    p1_smul_89586 <= p1_smul_89586_comb;
    p1_smul_90025 <= p1_smul_90025_comb;
    p1_smul_90026 <= p1_smul_90026_comb;
    p1_smul_90027 <= p1_smul_90027_comb;
    p1_smul_90028 <= p1_smul_90028_comb;
    p1_smul_90029 <= p1_smul_90029_comb;
    p1_smul_90030 <= p1_smul_90030_comb;
    p1_smul_89587 <= p1_smul_89587_comb;
    p1_smul_89588 <= p1_smul_89588_comb;
    p1_smul_89589 <= p1_smul_89589_comb;
    p1_smul_89590 <= p1_smul_89590_comb;
    p1_smul_90031 <= p1_smul_90031_comb;
    p1_smul_90032 <= p1_smul_90032_comb;
    p1_smul_90033 <= p1_smul_90033_comb;
    p1_smul_90034 <= p1_smul_90034_comb;
    p1_smul_90035 <= p1_smul_90035_comb;
    p1_smul_90036 <= p1_smul_90036_comb;
    p1_smul_89591 <= p1_smul_89591_comb;
    p1_smul_89592 <= p1_smul_89592_comb;
    p1_smul_89593 <= p1_smul_89593_comb;
    p1_smul_89594 <= p1_smul_89594_comb;
    p1_smul_90037 <= p1_smul_90037_comb;
    p1_smul_90038 <= p1_smul_90038_comb;
    p1_smul_90039 <= p1_smul_90039_comb;
    p1_smul_90040 <= p1_smul_90040_comb;
    p1_smul_90041 <= p1_smul_90041_comb;
    p1_smul_90042 <= p1_smul_90042_comb;
    p1_smul_89595 <= p1_smul_89595_comb;
    p1_smul_89596 <= p1_smul_89596_comb;
    p1_smul_89597 <= p1_smul_89597_comb;
    p1_smul_89598 <= p1_smul_89598_comb;
    p1_smul_90043 <= p1_smul_90043_comb;
    p1_smul_90044 <= p1_smul_90044_comb;
    p1_smul_90045 <= p1_smul_90045_comb;
    p1_smul_90046 <= p1_smul_90046_comb;
    p1_smul_90047 <= p1_smul_90047_comb;
    p1_smul_90048 <= p1_smul_90048_comb;
    p1_smul_89599 <= p1_smul_89599_comb;
    p1_smul_89600 <= p1_smul_89600_comb;
    p1_smul_89601 <= p1_smul_89601_comb;
    p1_smul_89602 <= p1_smul_89602_comb;
    p1_smul_90049 <= p1_smul_90049_comb;
    p1_smul_90050 <= p1_smul_90050_comb;
    p1_smul_90051 <= p1_smul_90051_comb;
    p1_smul_90052 <= p1_smul_90052_comb;
    p1_smul_90053 <= p1_smul_90053_comb;
    p1_smul_90054 <= p1_smul_90054_comb;
    p1_smul_89603 <= p1_smul_89603_comb;
    p1_smul_89604 <= p1_smul_89604_comb;
    p1_smul_89605 <= p1_smul_89605_comb;
    p1_smul_89606 <= p1_smul_89606_comb;
    p1_smul_90055 <= p1_smul_90055_comb;
    p1_smul_90056 <= p1_smul_90056_comb;
    p1_smul_90057 <= p1_smul_90057_comb;
    p1_smul_90058 <= p1_smul_90058_comb;
    p1_smul_90059 <= p1_smul_90059_comb;
    p1_smul_90060 <= p1_smul_90060_comb;
    p1_smul_89607 <= p1_smul_89607_comb;
    p1_smul_89608 <= p1_smul_89608_comb;
    p1_smul_89609 <= p1_smul_89609_comb;
    p1_smul_89610 <= p1_smul_89610_comb;
    p1_smul_90061 <= p1_smul_90061_comb;
    p1_smul_90062 <= p1_smul_90062_comb;
    p1_smul_90063 <= p1_smul_90063_comb;
    p1_smul_90064 <= p1_smul_90064_comb;
    p1_smul_90065 <= p1_smul_90065_comb;
    p1_smul_90066 <= p1_smul_90066_comb;
    p1_smul_89611 <= p1_smul_89611_comb;
    p1_smul_89612 <= p1_smul_89612_comb;
    p1_smul_89613 <= p1_smul_89613_comb;
    p1_smul_89614 <= p1_smul_89614_comb;
    p1_smul_90067 <= p1_smul_90067_comb;
    p1_smul_90068 <= p1_smul_90068_comb;
    p1_smul_90069 <= p1_smul_90069_comb;
    p1_smul_90070 <= p1_smul_90070_comb;
    p1_smul_90071 <= p1_smul_90071_comb;
    p1_smul_90072 <= p1_smul_90072_comb;
    p1_smul_89615 <= p1_smul_89615_comb;
    p1_smul_89616 <= p1_smul_89616_comb;
    p1_smul_89617 <= p1_smul_89617_comb;
    p1_smul_89618 <= p1_smul_89618_comb;
    p1_smul_90073 <= p1_smul_90073_comb;
    p1_smul_90074 <= p1_smul_90074_comb;
    p1_smul_90075 <= p1_smul_90075_comb;
    p1_smul_90076 <= p1_smul_90076_comb;
    p1_smul_90077 <= p1_smul_90077_comb;
    p1_smul_90078 <= p1_smul_90078_comb;
    p1_smul_89619 <= p1_smul_89619_comb;
    p1_smul_89620 <= p1_smul_89620_comb;
    p1_smul_89621 <= p1_smul_89621_comb;
    p1_smul_89622 <= p1_smul_89622_comb;
    p1_smul_90079 <= p1_smul_90079_comb;
    p1_smul_90080 <= p1_smul_90080_comb;
    p1_smul_90081 <= p1_smul_90081_comb;
    p1_smul_90082 <= p1_smul_90082_comb;
    p1_smul_90083 <= p1_smul_90083_comb;
    p1_smul_90084 <= p1_smul_90084_comb;
    p1_smul_89623 <= p1_smul_89623_comb;
    p1_smul_89624 <= p1_smul_89624_comb;
    p1_smul_89625 <= p1_smul_89625_comb;
    p1_smul_89626 <= p1_smul_89626_comb;
    p1_smul_90085 <= p1_smul_90085_comb;
    p1_smul_90086 <= p1_smul_90086_comb;
    p1_smul_90087 <= p1_smul_90087_comb;
    p1_smul_90088 <= p1_smul_90088_comb;
    p1_smul_90089 <= p1_smul_90089_comb;
    p1_smul_90090 <= p1_smul_90090_comb;
    p1_smul_89627 <= p1_smul_89627_comb;
    p1_smul_89628 <= p1_smul_89628_comb;
    p1_smul_89629 <= p1_smul_89629_comb;
    p1_smul_89630 <= p1_smul_89630_comb;
    p1_smul_90091 <= p1_smul_90091_comb;
    p1_smul_90092 <= p1_smul_90092_comb;
    p1_smul_90093 <= p1_smul_90093_comb;
    p1_smul_90094 <= p1_smul_90094_comb;
    p1_smul_90095 <= p1_smul_90095_comb;
    p1_smul_90096 <= p1_smul_90096_comb;
    p1_smul_89631 <= p1_smul_89631_comb;
    p1_smul_89632 <= p1_smul_89632_comb;
    p1_smul_89633 <= p1_smul_89633_comb;
    p1_smul_89634 <= p1_smul_89634_comb;
    p1_smul_90097 <= p1_smul_90097_comb;
    p1_smul_90098 <= p1_smul_90098_comb;
    p1_smul_90099 <= p1_smul_90099_comb;
    p1_smul_90100 <= p1_smul_90100_comb;
    p1_smul_90101 <= p1_smul_90101_comb;
    p1_smul_90102 <= p1_smul_90102_comb;
    p1_smul_89635 <= p1_smul_89635_comb;
    p1_smul_89636 <= p1_smul_89636_comb;
    p1_smul_89637 <= p1_smul_89637_comb;
    p1_smul_89638 <= p1_smul_89638_comb;
    p1_smul_90103 <= p1_smul_90103_comb;
    p1_smul_90104 <= p1_smul_90104_comb;
    p1_smul_90105 <= p1_smul_90105_comb;
    p1_smul_90106 <= p1_smul_90106_comb;
    p1_smul_90107 <= p1_smul_90107_comb;
    p1_smul_90108 <= p1_smul_90108_comb;
    p1_smul_89639 <= p1_smul_89639_comb;
    p1_smul_89640 <= p1_smul_89640_comb;
    p1_smul_89641 <= p1_smul_89641_comb;
    p1_smul_89642 <= p1_smul_89642_comb;
    p1_smul_90109 <= p1_smul_90109_comb;
    p1_smul_90110 <= p1_smul_90110_comb;
    p1_smul_90111 <= p1_smul_90111_comb;
    p1_smul_90112 <= p1_smul_90112_comb;
    p1_smul_90113 <= p1_smul_90113_comb;
    p1_smul_90114 <= p1_smul_90114_comb;
    p1_smul_89643 <= p1_smul_89643_comb;
    p1_smul_89644 <= p1_smul_89644_comb;
    p1_smul_89645 <= p1_smul_89645_comb;
    p1_smul_89646 <= p1_smul_89646_comb;
    p1_smul_90115 <= p1_smul_90115_comb;
    p1_smul_90116 <= p1_smul_90116_comb;
    p1_smul_90117 <= p1_smul_90117_comb;
    p1_smul_90118 <= p1_smul_90118_comb;
    p1_smul_90119 <= p1_smul_90119_comb;
    p1_smul_90120 <= p1_smul_90120_comb;
    p1_smul_89647 <= p1_smul_89647_comb;
    p1_smul_89648 <= p1_smul_89648_comb;
    p1_smul_89649 <= p1_smul_89649_comb;
    p1_smul_89650 <= p1_smul_89650_comb;
    p1_smul_90121 <= p1_smul_90121_comb;
    p1_smul_90122 <= p1_smul_90122_comb;
    p1_smul_90123 <= p1_smul_90123_comb;
    p1_smul_90124 <= p1_smul_90124_comb;
    p1_smul_90125 <= p1_smul_90125_comb;
    p1_smul_90126 <= p1_smul_90126_comb;
    p1_smul_89651 <= p1_smul_89651_comb;
    p1_smul_89652 <= p1_smul_89652_comb;
    p1_smul_89653 <= p1_smul_89653_comb;
    p1_smul_89654 <= p1_smul_89654_comb;
    p1_smul_90127 <= p1_smul_90127_comb;
    p1_smul_90128 <= p1_smul_90128_comb;
    p1_smul_90129 <= p1_smul_90129_comb;
    p1_smul_90130 <= p1_smul_90130_comb;
    p1_smul_90131 <= p1_smul_90131_comb;
    p1_smul_90132 <= p1_smul_90132_comb;
    p1_smul_89655 <= p1_smul_89655_comb;
    p1_smul_89656 <= p1_smul_89656_comb;
    p1_smul_89657 <= p1_smul_89657_comb;
    p1_smul_89658 <= p1_smul_89658_comb;
    p1_smul_90133 <= p1_smul_90133_comb;
    p1_smul_90134 <= p1_smul_90134_comb;
    p1_smul_90135 <= p1_smul_90135_comb;
    p1_smul_90136 <= p1_smul_90136_comb;
    p1_smul_90137 <= p1_smul_90137_comb;
    p1_smul_90138 <= p1_smul_90138_comb;
    p1_smul_89659 <= p1_smul_89659_comb;
    p1_smul_89660 <= p1_smul_89660_comb;
    p1_smul_89661 <= p1_smul_89661_comb;
    p1_smul_89662 <= p1_smul_89662_comb;
    p1_smul_90139 <= p1_smul_90139_comb;
    p1_smul_90140 <= p1_smul_90140_comb;
    p1_smul_90141 <= p1_smul_90141_comb;
    p1_smul_90142 <= p1_smul_90142_comb;
    p1_smul_90143 <= p1_smul_90143_comb;
    p1_smul_90144 <= p1_smul_90144_comb;
    p1_smul_89663 <= p1_smul_89663_comb;
    p1_smul_89664 <= p1_smul_89664_comb;
    p1_smul_89665 <= p1_smul_89665_comb;
    p1_smul_89666 <= p1_smul_89666_comb;
    p1_smul_90145 <= p1_smul_90145_comb;
    p1_smul_90146 <= p1_smul_90146_comb;
    p1_smul_90147 <= p1_smul_90147_comb;
    p1_smul_90148 <= p1_smul_90148_comb;
    p1_smul_90149 <= p1_smul_90149_comb;
    p1_smul_90150 <= p1_smul_90150_comb;
    p1_smul_89667 <= p1_smul_89667_comb;
    p1_smul_89668 <= p1_smul_89668_comb;
    p1_smul_89669 <= p1_smul_89669_comb;
    p1_smul_89670 <= p1_smul_89670_comb;
    p1_smul_90151 <= p1_smul_90151_comb;
    p1_smul_90152 <= p1_smul_90152_comb;
    p1_smul_90153 <= p1_smul_90153_comb;
    p1_smul_90154 <= p1_smul_90154_comb;
    p1_smul_90155 <= p1_smul_90155_comb;
    p1_smul_90156 <= p1_smul_90156_comb;
    p1_smul_89671 <= p1_smul_89671_comb;
    p1_smul_89672 <= p1_smul_89672_comb;
    p1_smul_89673 <= p1_smul_89673_comb;
    p1_smul_89674 <= p1_smul_89674_comb;
    p1_smul_90157 <= p1_smul_90157_comb;
    p1_smul_90158 <= p1_smul_90158_comb;
    p1_smul_90159 <= p1_smul_90159_comb;
    p1_smul_90160 <= p1_smul_90160_comb;
    p1_smul_90161 <= p1_smul_90161_comb;
    p1_smul_90162 <= p1_smul_90162_comb;
    p1_smul_89675 <= p1_smul_89675_comb;
    p1_smul_89676 <= p1_smul_89676_comb;
    p1_smul_89677 <= p1_smul_89677_comb;
    p1_smul_89678 <= p1_smul_89678_comb;
    p1_smul_90163 <= p1_smul_90163_comb;
    p1_smul_90164 <= p1_smul_90164_comb;
    p1_smul_90165 <= p1_smul_90165_comb;
    p1_smul_90166 <= p1_smul_90166_comb;
    p1_smul_90167 <= p1_smul_90167_comb;
    p1_smul_90168 <= p1_smul_90168_comb;
    p1_smul_89679 <= p1_smul_89679_comb;
    p1_smul_89680 <= p1_smul_89680_comb;
    p1_smul_89681 <= p1_smul_89681_comb;
    p1_smul_89682 <= p1_smul_89682_comb;
    p1_smul_90169 <= p1_smul_90169_comb;
    p1_smul_90170 <= p1_smul_90170_comb;
    p1_smul_90171 <= p1_smul_90171_comb;
    p1_smul_90172 <= p1_smul_90172_comb;
    p1_smul_90173 <= p1_smul_90173_comb;
    p1_smul_90174 <= p1_smul_90174_comb;
    p1_smul_89683 <= p1_smul_89683_comb;
    p1_smul_89684 <= p1_smul_89684_comb;
    p1_smul_89685 <= p1_smul_89685_comb;
    p1_smul_89686 <= p1_smul_89686_comb;
    p1_smul_90175 <= p1_smul_90175_comb;
    p1_smul_90176 <= p1_smul_90176_comb;
    p1_smul_90177 <= p1_smul_90177_comb;
    p1_smul_90178 <= p1_smul_90178_comb;
    p1_smul_90179 <= p1_smul_90179_comb;
    p1_smul_90180 <= p1_smul_90180_comb;
    p1_smul_89687 <= p1_smul_89687_comb;
    p1_smul_89688 <= p1_smul_89688_comb;
    p1_smul_89689 <= p1_smul_89689_comb;
    p1_smul_89690 <= p1_smul_89690_comb;
    p1_smul_90181 <= p1_smul_90181_comb;
    p1_smul_90182 <= p1_smul_90182_comb;
    p1_smul_90183 <= p1_smul_90183_comb;
    p1_smul_90184 <= p1_smul_90184_comb;
    p1_smul_90185 <= p1_smul_90185_comb;
    p1_smul_90186 <= p1_smul_90186_comb;
    p1_smul_89691 <= p1_smul_89691_comb;
    p1_smul_89692 <= p1_smul_89692_comb;
    p1_smul_89693 <= p1_smul_89693_comb;
    p1_smul_89694 <= p1_smul_89694_comb;
    p1_smul_90187 <= p1_smul_90187_comb;
    p1_smul_90188 <= p1_smul_90188_comb;
    p1_smul_90189 <= p1_smul_90189_comb;
    p1_smul_90190 <= p1_smul_90190_comb;
    p1_smul_90191 <= p1_smul_90191_comb;
    p1_smul_90192 <= p1_smul_90192_comb;
    p1_smul_89695 <= p1_smul_89695_comb;
    p1_smul_89696 <= p1_smul_89696_comb;
    p1_smul_89697 <= p1_smul_89697_comb;
    p1_smul_89698 <= p1_smul_89698_comb;
    p1_smul_90193 <= p1_smul_90193_comb;
    p1_smul_90194 <= p1_smul_90194_comb;
    p1_smul_90195 <= p1_smul_90195_comb;
    p1_smul_90196 <= p1_smul_90196_comb;
    p1_smul_90197 <= p1_smul_90197_comb;
    p1_smul_90198 <= p1_smul_90198_comb;
    p1_smul_89699 <= p1_smul_89699_comb;
    p1_smul_89700 <= p1_smul_89700_comb;
    p1_smul_89701 <= p1_smul_89701_comb;
    p1_smul_89702 <= p1_smul_89702_comb;
    p1_smul_90199 <= p1_smul_90199_comb;
    p1_smul_90200 <= p1_smul_90200_comb;
    p1_smul_90201 <= p1_smul_90201_comb;
    p1_smul_90202 <= p1_smul_90202_comb;
    p1_smul_90203 <= p1_smul_90203_comb;
    p1_smul_90204 <= p1_smul_90204_comb;
    p1_smul_89703 <= p1_smul_89703_comb;
    p1_smul_89704 <= p1_smul_89704_comb;
    p1_smul_89705 <= p1_smul_89705_comb;
    p1_smul_89706 <= p1_smul_89706_comb;
    p1_smul_90205 <= p1_smul_90205_comb;
    p1_smul_90206 <= p1_smul_90206_comb;
    p1_smul_90207 <= p1_smul_90207_comb;
    p1_smul_90208 <= p1_smul_90208_comb;
    p1_smul_90209 <= p1_smul_90209_comb;
    p1_smul_90210 <= p1_smul_90210_comb;
    p1_smul_89707 <= p1_smul_89707_comb;
    p1_smul_89708 <= p1_smul_89708_comb;
    p1_smul_89709 <= p1_smul_89709_comb;
    p1_smul_89710 <= p1_smul_89710_comb;
    p1_smul_90211 <= p1_smul_90211_comb;
    p1_smul_90212 <= p1_smul_90212_comb;
    p1_smul_90213 <= p1_smul_90213_comb;
    p1_smul_90214 <= p1_smul_90214_comb;
    p1_smul_90215 <= p1_smul_90215_comb;
    p1_smul_90216 <= p1_smul_90216_comb;
    p1_smul_89711 <= p1_smul_89711_comb;
    p1_smul_89712 <= p1_smul_89712_comb;
    p1_smul_89713 <= p1_smul_89713_comb;
    p1_smul_89714 <= p1_smul_89714_comb;
    p1_smul_90217 <= p1_smul_90217_comb;
    p1_smul_90218 <= p1_smul_90218_comb;
    p1_smul_90219 <= p1_smul_90219_comb;
    p1_smul_90220 <= p1_smul_90220_comb;
    p1_smul_90221 <= p1_smul_90221_comb;
    p1_smul_90222 <= p1_smul_90222_comb;
    p1_smul_89715 <= p1_smul_89715_comb;
    p1_smul_89716 <= p1_smul_89716_comb;
    p1_smul_89717 <= p1_smul_89717_comb;
    p1_smul_89718 <= p1_smul_89718_comb;
    p1_smul_90223 <= p1_smul_90223_comb;
    p1_smul_90224 <= p1_smul_90224_comb;
    p1_smul_90225 <= p1_smul_90225_comb;
    p1_smul_90226 <= p1_smul_90226_comb;
    p1_smul_90227 <= p1_smul_90227_comb;
    p1_smul_90228 <= p1_smul_90228_comb;
    p1_smul_89719 <= p1_smul_89719_comb;
    p1_smul_89720 <= p1_smul_89720_comb;
    p1_smul_89721 <= p1_smul_89721_comb;
    p1_smul_89722 <= p1_smul_89722_comb;
    p1_smul_90229 <= p1_smul_90229_comb;
    p1_smul_90230 <= p1_smul_90230_comb;
    p1_smul_90231 <= p1_smul_90231_comb;
    p1_smul_90232 <= p1_smul_90232_comb;
    p1_smul_90233 <= p1_smul_90233_comb;
    p1_smul_90234 <= p1_smul_90234_comb;
    p1_smul_89723 <= p1_smul_89723_comb;
    p1_smul_89724 <= p1_smul_89724_comb;
    p1_smul_89725 <= p1_smul_89725_comb;
    p1_smul_89726 <= p1_smul_89726_comb;
    p1_smul_90235 <= p1_smul_90235_comb;
    p1_smul_90236 <= p1_smul_90236_comb;
    p1_smul_90237 <= p1_smul_90237_comb;
    p1_smul_90238 <= p1_smul_90238_comb;
    p1_smul_90239 <= p1_smul_90239_comb;
    p1_smul_90240 <= p1_smul_90240_comb;
    p1_smul_89727 <= p1_smul_89727_comb;
    p1_smul_89728 <= p1_smul_89728_comb;
    p1_smul_89729 <= p1_smul_89729_comb;
    p1_smul_89730 <= p1_smul_89730_comb;
    p1_smul_90241 <= p1_smul_90241_comb;
    p1_smul_90242 <= p1_smul_90242_comb;
    p1_smul_90243 <= p1_smul_90243_comb;
    p1_smul_90244 <= p1_smul_90244_comb;
    p1_smul_90245 <= p1_smul_90245_comb;
    p1_smul_90246 <= p1_smul_90246_comb;
    p1_smul_89731 <= p1_smul_89731_comb;
    p1_smul_89732 <= p1_smul_89732_comb;
    p1_smul_89733 <= p1_smul_89733_comb;
    p1_smul_89734 <= p1_smul_89734_comb;
    p1_smul_90247 <= p1_smul_90247_comb;
    p1_smul_90248 <= p1_smul_90248_comb;
    p1_smul_90249 <= p1_smul_90249_comb;
    p1_smul_90250 <= p1_smul_90250_comb;
    p1_smul_90251 <= p1_smul_90251_comb;
    p1_smul_90252 <= p1_smul_90252_comb;
    p1_smul_89735 <= p1_smul_89735_comb;
    p1_smul_89736 <= p1_smul_89736_comb;
    p1_smul_89737 <= p1_smul_89737_comb;
    p1_smul_89738 <= p1_smul_89738_comb;
    p1_smul_90253 <= p1_smul_90253_comb;
    p1_smul_90254 <= p1_smul_90254_comb;
    p1_smul_90255 <= p1_smul_90255_comb;
    p1_smul_90256 <= p1_smul_90256_comb;
    p1_smul_90257 <= p1_smul_90257_comb;
    p1_smul_90258 <= p1_smul_90258_comb;
    p1_smul_89739 <= p1_smul_89739_comb;
    p1_smul_89740 <= p1_smul_89740_comb;
    p1_smul_89741 <= p1_smul_89741_comb;
    p1_smul_89742 <= p1_smul_89742_comb;
    p1_smul_90259 <= p1_smul_90259_comb;
    p1_smul_90260 <= p1_smul_90260_comb;
    p1_smul_90261 <= p1_smul_90261_comb;
    p1_smul_90262 <= p1_smul_90262_comb;
    p1_smul_90263 <= p1_smul_90263_comb;
    p1_smul_90264 <= p1_smul_90264_comb;
    p1_smul_89743 <= p1_smul_89743_comb;
    p1_smul_89744 <= p1_smul_89744_comb;
    p1_smul_89745 <= p1_smul_89745_comb;
    p1_smul_89746 <= p1_smul_89746_comb;
    p1_smul_90265 <= p1_smul_90265_comb;
    p1_smul_90266 <= p1_smul_90266_comb;
    p1_smul_90267 <= p1_smul_90267_comb;
    p1_smul_90268 <= p1_smul_90268_comb;
    p1_smul_90269 <= p1_smul_90269_comb;
    p1_smul_90270 <= p1_smul_90270_comb;
    p1_smul_89747 <= p1_smul_89747_comb;
    p1_smul_89748 <= p1_smul_89748_comb;
    p1_smul_89749 <= p1_smul_89749_comb;
    p1_smul_89750 <= p1_smul_89750_comb;
    p1_smul_90271 <= p1_smul_90271_comb;
    p1_smul_90272 <= p1_smul_90272_comb;
    p1_smul_90273 <= p1_smul_90273_comb;
    p1_smul_90274 <= p1_smul_90274_comb;
    p1_smul_90275 <= p1_smul_90275_comb;
    p1_smul_90276 <= p1_smul_90276_comb;
    p1_smul_89751 <= p1_smul_89751_comb;
    p1_smul_89752 <= p1_smul_89752_comb;
    p1_smul_89753 <= p1_smul_89753_comb;
    p1_smul_89754 <= p1_smul_89754_comb;
    p1_smul_90277 <= p1_smul_90277_comb;
    p1_smul_90278 <= p1_smul_90278_comb;
    p1_smul_90279 <= p1_smul_90279_comb;
    p1_smul_90280 <= p1_smul_90280_comb;
    p1_smul_90281 <= p1_smul_90281_comb;
    p1_smul_90282 <= p1_smul_90282_comb;
    p1_smul_89755 <= p1_smul_89755_comb;
    p1_smul_89756 <= p1_smul_89756_comb;
    p1_smul_89757 <= p1_smul_89757_comb;
    p1_smul_89758 <= p1_smul_89758_comb;
    p1_smul_90283 <= p1_smul_90283_comb;
    p1_smul_90284 <= p1_smul_90284_comb;
    p1_smul_90285 <= p1_smul_90285_comb;
    p1_smul_90286 <= p1_smul_90286_comb;
    p1_smul_90287 <= p1_smul_90287_comb;
    p1_smul_90288 <= p1_smul_90288_comb;
    p1_smul_89759 <= p1_smul_89759_comb;
    p1_smul_89760 <= p1_smul_89760_comb;
    p1_smul_89761 <= p1_smul_89761_comb;
    p1_smul_89762 <= p1_smul_89762_comb;
    p1_smul_90289 <= p1_smul_90289_comb;
    p1_smul_90290 <= p1_smul_90290_comb;
    p1_smul_90291 <= p1_smul_90291_comb;
    p1_smul_90292 <= p1_smul_90292_comb;
    p1_smul_90293 <= p1_smul_90293_comb;
    p1_smul_90294 <= p1_smul_90294_comb;
    p1_smul_89763 <= p1_smul_89763_comb;
    p1_smul_89764 <= p1_smul_89764_comb;
    p1_smul_89765 <= p1_smul_89765_comb;
    p1_smul_89766 <= p1_smul_89766_comb;
    p1_smul_90295 <= p1_smul_90295_comb;
    p1_smul_90296 <= p1_smul_90296_comb;
    p1_smul_90297 <= p1_smul_90297_comb;
    p1_smul_90298 <= p1_smul_90298_comb;
    p1_smul_90299 <= p1_smul_90299_comb;
    p1_smul_90300 <= p1_smul_90300_comb;
    p1_smul_89767 <= p1_smul_89767_comb;
    p1_smul_89768 <= p1_smul_89768_comb;
    p1_smul_89769 <= p1_smul_89769_comb;
    p1_smul_89770 <= p1_smul_89770_comb;
    p1_smul_90301 <= p1_smul_90301_comb;
    p1_smul_90302 <= p1_smul_90302_comb;
    p1_smul_90303 <= p1_smul_90303_comb;
    p1_smul_90304 <= p1_smul_90304_comb;
    p1_smul_90305 <= p1_smul_90305_comb;
    p1_smul_90306 <= p1_smul_90306_comb;
    p1_smul_89771 <= p1_smul_89771_comb;
    p1_smul_89772 <= p1_smul_89772_comb;
    p1_smul_89773 <= p1_smul_89773_comb;
    p1_smul_89774 <= p1_smul_89774_comb;
    p1_smul_90307 <= p1_smul_90307_comb;
    p1_smul_90308 <= p1_smul_90308_comb;
    p1_smul_90309 <= p1_smul_90309_comb;
    p1_smul_90310 <= p1_smul_90310_comb;
    p1_smul_90311 <= p1_smul_90311_comb;
    p1_smul_90312 <= p1_smul_90312_comb;
    p1_smul_89775 <= p1_smul_89775_comb;
    p1_smul_89776 <= p1_smul_89776_comb;
    p1_smul_89777 <= p1_smul_89777_comb;
    p1_smul_89778 <= p1_smul_89778_comb;
    p1_smul_90313 <= p1_smul_90313_comb;
    p1_smul_90314 <= p1_smul_90314_comb;
    p1_smul_90315 <= p1_smul_90315_comb;
    p1_smul_90316 <= p1_smul_90316_comb;
    p1_smul_90317 <= p1_smul_90317_comb;
    p1_smul_90318 <= p1_smul_90318_comb;
    p1_smul_89779 <= p1_smul_89779_comb;
    p1_smul_89780 <= p1_smul_89780_comb;
    p1_smul_89781 <= p1_smul_89781_comb;
    p1_smul_89782 <= p1_smul_89782_comb;
    p1_smul_90319 <= p1_smul_90319_comb;
    p1_smul_90320 <= p1_smul_90320_comb;
    p1_smul_90321 <= p1_smul_90321_comb;
    p1_smul_90322 <= p1_smul_90322_comb;
    p1_smul_90323 <= p1_smul_90323_comb;
    p1_smul_90324 <= p1_smul_90324_comb;
    p1_smul_89783 <= p1_smul_89783_comb;
    p1_smul_89784 <= p1_smul_89784_comb;
    p1_smul_89785 <= p1_smul_89785_comb;
    p1_smul_89786 <= p1_smul_89786_comb;
    p1_smul_90325 <= p1_smul_90325_comb;
    p1_smul_90326 <= p1_smul_90326_comb;
    p1_smul_90327 <= p1_smul_90327_comb;
    p1_smul_90328 <= p1_smul_90328_comb;
    p1_smul_90329 <= p1_smul_90329_comb;
    p1_smul_90330 <= p1_smul_90330_comb;
    p1_smul_89787 <= p1_smul_89787_comb;
    p1_smul_89788 <= p1_smul_89788_comb;
    p1_smul_89789 <= p1_smul_89789_comb;
    p1_smul_89790 <= p1_smul_89790_comb;
    p1_smul_90331 <= p1_smul_90331_comb;
    p1_smul_90332 <= p1_smul_90332_comb;
    p1_smul_90333 <= p1_smul_90333_comb;
    p1_smul_90334 <= p1_smul_90334_comb;
    p1_smul_90335 <= p1_smul_90335_comb;
    p1_smul_90336 <= p1_smul_90336_comb;
    p1_smul_89791 <= p1_smul_89791_comb;
    p1_smul_89792 <= p1_smul_89792_comb;
    p1_smul_89793 <= p1_smul_89793_comb;
    p1_smul_89794 <= p1_smul_89794_comb;
    p1_smul_90337 <= p1_smul_90337_comb;
    p1_smul_90338 <= p1_smul_90338_comb;
    p1_smul_90339 <= p1_smul_90339_comb;
    p1_smul_90340 <= p1_smul_90340_comb;
    p1_smul_90341 <= p1_smul_90341_comb;
    p1_smul_90342 <= p1_smul_90342_comb;
    p1_smul_89795 <= p1_smul_89795_comb;
    p1_smul_89796 <= p1_smul_89796_comb;
    p1_smul_89797 <= p1_smul_89797_comb;
    p1_smul_89798 <= p1_smul_89798_comb;
    p1_smul_90343 <= p1_smul_90343_comb;
    p1_smul_90344 <= p1_smul_90344_comb;
    p1_smul_90345 <= p1_smul_90345_comb;
    p1_smul_90346 <= p1_smul_90346_comb;
    p1_smul_90347 <= p1_smul_90347_comb;
    p1_smul_90348 <= p1_smul_90348_comb;
    p1_smul_89799 <= p1_smul_89799_comb;
    p1_smul_89800 <= p1_smul_89800_comb;
    p1_smul_89801 <= p1_smul_89801_comb;
    p1_smul_89802 <= p1_smul_89802_comb;
    p1_smul_90349 <= p1_smul_90349_comb;
    p1_smul_90350 <= p1_smul_90350_comb;
    p1_smul_90351 <= p1_smul_90351_comb;
    p1_smul_90352 <= p1_smul_90352_comb;
    p1_smul_90353 <= p1_smul_90353_comb;
    p1_smul_90354 <= p1_smul_90354_comb;
    p1_smul_89803 <= p1_smul_89803_comb;
    p1_smul_89804 <= p1_smul_89804_comb;
    p1_smul_89805 <= p1_smul_89805_comb;
    p1_smul_89806 <= p1_smul_89806_comb;
    p1_smul_90355 <= p1_smul_90355_comb;
    p1_smul_90356 <= p1_smul_90356_comb;
    p1_smul_90357 <= p1_smul_90357_comb;
    p1_smul_90358 <= p1_smul_90358_comb;
    p1_smul_90359 <= p1_smul_90359_comb;
    p1_smul_90360 <= p1_smul_90360_comb;
    p1_smul_89807 <= p1_smul_89807_comb;
    p1_smul_89808 <= p1_smul_89808_comb;
    p1_smul_89809 <= p1_smul_89809_comb;
    p1_smul_89810 <= p1_smul_89810_comb;
    p1_smul_90361 <= p1_smul_90361_comb;
    p1_smul_90362 <= p1_smul_90362_comb;
    p1_smul_90363 <= p1_smul_90363_comb;
    p1_smul_90364 <= p1_smul_90364_comb;
    p1_smul_90365 <= p1_smul_90365_comb;
    p1_smul_90366 <= p1_smul_90366_comb;
    p1_smul_89811 <= p1_smul_89811_comb;
    p1_smul_89812 <= p1_smul_89812_comb;
    p1_smul_89813 <= p1_smul_89813_comb;
    p1_smul_89814 <= p1_smul_89814_comb;
    p1_smul_90367 <= p1_smul_90367_comb;
    p1_smul_90368 <= p1_smul_90368_comb;
    p1_smul_90369 <= p1_smul_90369_comb;
    p1_smul_90370 <= p1_smul_90370_comb;
    p1_smul_90371 <= p1_smul_90371_comb;
    p1_smul_90372 <= p1_smul_90372_comb;
    p1_smul_89815 <= p1_smul_89815_comb;
    p1_smul_89816 <= p1_smul_89816_comb;
    p1_smul_89817 <= p1_smul_89817_comb;
    p1_smul_89818 <= p1_smul_89818_comb;
    p1_smul_90373 <= p1_smul_90373_comb;
    p1_smul_90374 <= p1_smul_90374_comb;
    p1_smul_90375 <= p1_smul_90375_comb;
    p1_smul_90376 <= p1_smul_90376_comb;
    p1_smul_90377 <= p1_smul_90377_comb;
    p1_smul_90378 <= p1_smul_90378_comb;
    p1_smul_89819 <= p1_smul_89819_comb;
    p1_smul_89820 <= p1_smul_89820_comb;
    p1_smul_89821 <= p1_smul_89821_comb;
    p1_smul_89822 <= p1_smul_89822_comb;
    p1_smul_90379 <= p1_smul_90379_comb;
    p1_smul_90380 <= p1_smul_90380_comb;
    p1_smul_90381 <= p1_smul_90381_comb;
    p1_smul_90382 <= p1_smul_90382_comb;
    p1_smul_90383 <= p1_smul_90383_comb;
    p1_smul_90384 <= p1_smul_90384_comb;
    p1_smul_89823 <= p1_smul_89823_comb;
    p1_smul_89824 <= p1_smul_89824_comb;
    p1_smul_89825 <= p1_smul_89825_comb;
    p1_smul_89826 <= p1_smul_89826_comb;
    p1_smul_90385 <= p1_smul_90385_comb;
    p1_smul_90386 <= p1_smul_90386_comb;
    p1_smul_90387 <= p1_smul_90387_comb;
    p1_smul_90388 <= p1_smul_90388_comb;
    p1_smul_90389 <= p1_smul_90389_comb;
    p1_smul_90390 <= p1_smul_90390_comb;
    p1_smul_89827 <= p1_smul_89827_comb;
    p1_smul_89828 <= p1_smul_89828_comb;
    p1_smul_89829 <= p1_smul_89829_comb;
    p1_smul_89830 <= p1_smul_89830_comb;
    p1_smul_90391 <= p1_smul_90391_comb;
    p1_smul_90392 <= p1_smul_90392_comb;
    p1_smul_90393 <= p1_smul_90393_comb;
    p1_smul_90394 <= p1_smul_90394_comb;
    p1_smul_90395 <= p1_smul_90395_comb;
    p1_smul_90396 <= p1_smul_90396_comb;
    p1_smul_89831 <= p1_smul_89831_comb;
    p1_smul_89832 <= p1_smul_89832_comb;
    p1_smul_89833 <= p1_smul_89833_comb;
    p1_smul_89834 <= p1_smul_89834_comb;
    p1_smul_90397 <= p1_smul_90397_comb;
    p1_smul_90398 <= p1_smul_90398_comb;
    p1_smul_90399 <= p1_smul_90399_comb;
    p1_smul_90400 <= p1_smul_90400_comb;
    p1_smul_90401 <= p1_smul_90401_comb;
    p1_smul_90402 <= p1_smul_90402_comb;
    p1_smul_89835 <= p1_smul_89835_comb;
    p1_smul_89836 <= p1_smul_89836_comb;
    p1_smul_89837 <= p1_smul_89837_comb;
    p1_smul_89838 <= p1_smul_89838_comb;
    p1_smul_90403 <= p1_smul_90403_comb;
    p1_smul_90404 <= p1_smul_90404_comb;
    p1_smul_90405 <= p1_smul_90405_comb;
    p1_smul_90406 <= p1_smul_90406_comb;
    p1_smul_90407 <= p1_smul_90407_comb;
    p1_smul_90408 <= p1_smul_90408_comb;
    p1_smul_89839 <= p1_smul_89839_comb;
    p1_smul_89840 <= p1_smul_89840_comb;
    p1_smul_89841 <= p1_smul_89841_comb;
    p1_smul_89842 <= p1_smul_89842_comb;
    p1_smul_90409 <= p1_smul_90409_comb;
    p1_smul_90410 <= p1_smul_90410_comb;
    p1_smul_90411 <= p1_smul_90411_comb;
    p1_smul_90412 <= p1_smul_90412_comb;
    p1_smul_90413 <= p1_smul_90413_comb;
    p1_smul_90414 <= p1_smul_90414_comb;
    p1_smul_89843 <= p1_smul_89843_comb;
    p1_smul_89844 <= p1_smul_89844_comb;
    p1_smul_89845 <= p1_smul_89845_comb;
    p1_smul_89846 <= p1_smul_89846_comb;
    p1_smul_90415 <= p1_smul_90415_comb;
    p1_smul_90416 <= p1_smul_90416_comb;
    p1_smul_90417 <= p1_smul_90417_comb;
    p1_smul_90418 <= p1_smul_90418_comb;
    p1_smul_90419 <= p1_smul_90419_comb;
    p1_smul_90420 <= p1_smul_90420_comb;
    p1_smul_89847 <= p1_smul_89847_comb;
    p1_smul_89848 <= p1_smul_89848_comb;
    p1_smul_89849 <= p1_smul_89849_comb;
    p1_smul_89850 <= p1_smul_89850_comb;
    p1_smul_90421 <= p1_smul_90421_comb;
    p1_smul_90422 <= p1_smul_90422_comb;
    p1_smul_90423 <= p1_smul_90423_comb;
    p1_smul_90424 <= p1_smul_90424_comb;
    p1_smul_90425 <= p1_smul_90425_comb;
    p1_smul_90426 <= p1_smul_90426_comb;
    p1_smul_89851 <= p1_smul_89851_comb;
    p1_smul_89852 <= p1_smul_89852_comb;
    p1_smul_89853 <= p1_smul_89853_comb;
    p1_smul_89854 <= p1_smul_89854_comb;
    p1_smul_90427 <= p1_smul_90427_comb;
    p1_smul_90428 <= p1_smul_90428_comb;
    p1_smul_90429 <= p1_smul_90429_comb;
    p1_smul_90430 <= p1_smul_90430_comb;
    p1_smul_90431 <= p1_smul_90431_comb;
    p1_smul_90432 <= p1_smul_90432_comb;
    p1_smul_89855 <= p1_smul_89855_comb;
    p1_smul_89856 <= p1_smul_89856_comb;
    p1_smul_89857 <= p1_smul_89857_comb;
    p1_smul_89858 <= p1_smul_89858_comb;
    p1_smul_90433 <= p1_smul_90433_comb;
    p1_smul_90434 <= p1_smul_90434_comb;
    p1_smul_90435 <= p1_smul_90435_comb;
    p1_smul_90436 <= p1_smul_90436_comb;
    p1_smul_90437 <= p1_smul_90437_comb;
    p1_smul_90438 <= p1_smul_90438_comb;
    p1_smul_89859 <= p1_smul_89859_comb;
    p1_smul_89860 <= p1_smul_89860_comb;
    p1_smul_89861 <= p1_smul_89861_comb;
    p1_smul_89862 <= p1_smul_89862_comb;
    p1_smul_90439 <= p1_smul_90439_comb;
    p1_smul_90440 <= p1_smul_90440_comb;
    p1_smul_90441 <= p1_smul_90441_comb;
    p1_smul_90442 <= p1_smul_90442_comb;
    p1_smul_90443 <= p1_smul_90443_comb;
    p1_smul_90444 <= p1_smul_90444_comb;
    p1_smul_89863 <= p1_smul_89863_comb;
    p1_smul_89864 <= p1_smul_89864_comb;
    p1_smul_89865 <= p1_smul_89865_comb;
    p1_smul_89866 <= p1_smul_89866_comb;
    p1_smul_90445 <= p1_smul_90445_comb;
    p1_smul_90446 <= p1_smul_90446_comb;
    p1_smul_90447 <= p1_smul_90447_comb;
    p1_smul_90448 <= p1_smul_90448_comb;
    p1_smul_90449 <= p1_smul_90449_comb;
    p1_smul_90450 <= p1_smul_90450_comb;
    p1_smul_89867 <= p1_smul_89867_comb;
    p1_smul_89868 <= p1_smul_89868_comb;
    p1_smul_89869 <= p1_smul_89869_comb;
    p1_smul_89870 <= p1_smul_89870_comb;
    p1_smul_90451 <= p1_smul_90451_comb;
    p1_smul_90452 <= p1_smul_90452_comb;
    p1_smul_90453 <= p1_smul_90453_comb;
    p1_smul_90454 <= p1_smul_90454_comb;
    p1_smul_90455 <= p1_smul_90455_comb;
    p1_smul_90456 <= p1_smul_90456_comb;
    p1_smul_89871 <= p1_smul_89871_comb;
    p1_smul_89872 <= p1_smul_89872_comb;
    p1_smul_89873 <= p1_smul_89873_comb;
    p1_smul_89874 <= p1_smul_89874_comb;
    p1_smul_90457 <= p1_smul_90457_comb;
    p1_smul_90458 <= p1_smul_90458_comb;
    p1_smul_90459 <= p1_smul_90459_comb;
    p1_smul_90460 <= p1_smul_90460_comb;
    p1_smul_90461 <= p1_smul_90461_comb;
    p1_smul_90462 <= p1_smul_90462_comb;
    p1_smul_89875 <= p1_smul_89875_comb;
    p1_smul_89876 <= p1_smul_89876_comb;
    p1_smul_89877 <= p1_smul_89877_comb;
    p1_smul_89878 <= p1_smul_89878_comb;
    p1_smul_90463 <= p1_smul_90463_comb;
    p1_smul_90464 <= p1_smul_90464_comb;
    p1_smul_90465 <= p1_smul_90465_comb;
    p1_smul_90466 <= p1_smul_90466_comb;
    p1_smul_90467 <= p1_smul_90467_comb;
    p1_smul_90468 <= p1_smul_90468_comb;
    p1_smul_89879 <= p1_smul_89879_comb;
    p1_smul_89880 <= p1_smul_89880_comb;
    p1_smul_89881 <= p1_smul_89881_comb;
    p1_smul_89882 <= p1_smul_89882_comb;
    p1_smul_90469 <= p1_smul_90469_comb;
    p1_smul_90470 <= p1_smul_90470_comb;
    p1_smul_90471 <= p1_smul_90471_comb;
    p1_smul_90472 <= p1_smul_90472_comb;
    p1_smul_90473 <= p1_smul_90473_comb;
    p1_smul_90474 <= p1_smul_90474_comb;
    p1_smul_89883 <= p1_smul_89883_comb;
    p1_smul_89884 <= p1_smul_89884_comb;
    p1_smul_89885 <= p1_smul_89885_comb;
    p1_smul_89886 <= p1_smul_89886_comb;
    p1_smul_90475 <= p1_smul_90475_comb;
    p1_smul_90476 <= p1_smul_90476_comb;
    p1_smul_90477 <= p1_smul_90477_comb;
    p1_smul_90478 <= p1_smul_90478_comb;
    p1_smul_90479 <= p1_smul_90479_comb;
    p1_smul_90480 <= p1_smul_90480_comb;
    p1_smul_89887 <= p1_smul_89887_comb;
    p1_smul_89888 <= p1_smul_89888_comb;
    p1_smul_89889 <= p1_smul_89889_comb;
    p1_smul_89890 <= p1_smul_89890_comb;
    p1_smul_90481 <= p1_smul_90481_comb;
    p1_smul_90482 <= p1_smul_90482_comb;
    p1_smul_90483 <= p1_smul_90483_comb;
    p1_smul_90484 <= p1_smul_90484_comb;
    p1_smul_90485 <= p1_smul_90485_comb;
    p1_smul_90486 <= p1_smul_90486_comb;
    p1_smul_89891 <= p1_smul_89891_comb;
    p1_smul_89892 <= p1_smul_89892_comb;
    p1_smul_89893 <= p1_smul_89893_comb;
    p1_smul_89894 <= p1_smul_89894_comb;
    p1_smul_90487 <= p1_smul_90487_comb;
    p1_smul_90488 <= p1_smul_90488_comb;
    p1_smul_90489 <= p1_smul_90489_comb;
    p1_smul_90490 <= p1_smul_90490_comb;
    p1_smul_90491 <= p1_smul_90491_comb;
    p1_smul_90492 <= p1_smul_90492_comb;
    p1_smul_89895 <= p1_smul_89895_comb;
    p1_smul_89896 <= p1_smul_89896_comb;
    p1_smul_89897 <= p1_smul_89897_comb;
    p1_smul_89898 <= p1_smul_89898_comb;
    p1_smul_90493 <= p1_smul_90493_comb;
    p1_smul_90494 <= p1_smul_90494_comb;
    p1_smul_90495 <= p1_smul_90495_comb;
    p1_smul_90496 <= p1_smul_90496_comb;
    p1_smul_90497 <= p1_smul_90497_comb;
    p1_smul_90498 <= p1_smul_90498_comb;
  end

  // ===== Pipe stage 2:
  wire [31:0] p2_add_92711_comb;
  wire [31:0] p2_add_92712_comb;
  wire [31:0] p2_add_93111_comb;
  wire [31:0] p2_add_93112_comb;
  wire [31:0] p2_add_92709_comb;
  wire [31:0] p2_add_92710_comb;
  wire [31:0] p2_add_93107_comb;
  wire [31:0] p2_add_93108_comb;
  wire [31:0] p2_add_92707_comb;
  wire [31:0] p2_add_92708_comb;
  wire [31:0] p2_add_93103_comb;
  wire [31:0] p2_add_93104_comb;
  wire [31:0] p2_add_92705_comb;
  wire [31:0] p2_add_92706_comb;
  wire [31:0] p2_add_93099_comb;
  wire [31:0] p2_add_93100_comb;
  wire [31:0] p2_add_92703_comb;
  wire [31:0] p2_add_92704_comb;
  wire [31:0] p2_add_93095_comb;
  wire [31:0] p2_add_93096_comb;
  wire [31:0] p2_add_92701_comb;
  wire [31:0] p2_add_92702_comb;
  wire [31:0] p2_add_93091_comb;
  wire [31:0] p2_add_93092_comb;
  wire [31:0] p2_add_92699_comb;
  wire [31:0] p2_add_92700_comb;
  wire [31:0] p2_add_93087_comb;
  wire [31:0] p2_add_93088_comb;
  wire [31:0] p2_add_92697_comb;
  wire [31:0] p2_add_92698_comb;
  wire [31:0] p2_add_93083_comb;
  wire [31:0] p2_add_93084_comb;
  wire [31:0] p2_add_92695_comb;
  wire [31:0] p2_add_92696_comb;
  wire [31:0] p2_add_93079_comb;
  wire [31:0] p2_add_93080_comb;
  wire [31:0] p2_add_92693_comb;
  wire [31:0] p2_add_92694_comb;
  wire [31:0] p2_add_93075_comb;
  wire [31:0] p2_add_93076_comb;
  wire [31:0] p2_add_92691_comb;
  wire [31:0] p2_add_92692_comb;
  wire [31:0] p2_add_93071_comb;
  wire [31:0] p2_add_93072_comb;
  wire [31:0] p2_add_92689_comb;
  wire [31:0] p2_add_92690_comb;
  wire [31:0] p2_add_93067_comb;
  wire [31:0] p2_add_93068_comb;
  wire [31:0] p2_add_92687_comb;
  wire [31:0] p2_add_92688_comb;
  wire [31:0] p2_add_93063_comb;
  wire [31:0] p2_add_93064_comb;
  wire [31:0] p2_add_92685_comb;
  wire [31:0] p2_add_92686_comb;
  wire [31:0] p2_add_93059_comb;
  wire [31:0] p2_add_93060_comb;
  wire [31:0] p2_add_92683_comb;
  wire [31:0] p2_add_92684_comb;
  wire [31:0] p2_add_93055_comb;
  wire [31:0] p2_add_93056_comb;
  wire [31:0] p2_add_92681_comb;
  wire [31:0] p2_add_92682_comb;
  wire [31:0] p2_add_93051_comb;
  wire [31:0] p2_add_93052_comb;
  wire [31:0] p2_add_92679_comb;
  wire [31:0] p2_add_92680_comb;
  wire [31:0] p2_add_93047_comb;
  wire [31:0] p2_add_93048_comb;
  wire [31:0] p2_add_92677_comb;
  wire [31:0] p2_add_92678_comb;
  wire [31:0] p2_add_93043_comb;
  wire [31:0] p2_add_93044_comb;
  wire [31:0] p2_add_92675_comb;
  wire [31:0] p2_add_92676_comb;
  wire [31:0] p2_add_93039_comb;
  wire [31:0] p2_add_93040_comb;
  wire [31:0] p2_add_92673_comb;
  wire [31:0] p2_add_92674_comb;
  wire [31:0] p2_add_93035_comb;
  wire [31:0] p2_add_93036_comb;
  wire [31:0] p2_add_92671_comb;
  wire [31:0] p2_add_92672_comb;
  wire [31:0] p2_add_93031_comb;
  wire [31:0] p2_add_93032_comb;
  wire [31:0] p2_add_92669_comb;
  wire [31:0] p2_add_92670_comb;
  wire [31:0] p2_add_93027_comb;
  wire [31:0] p2_add_93028_comb;
  wire [31:0] p2_add_92667_comb;
  wire [31:0] p2_add_92668_comb;
  wire [31:0] p2_add_93023_comb;
  wire [31:0] p2_add_93024_comb;
  wire [31:0] p2_add_92665_comb;
  wire [31:0] p2_add_92666_comb;
  wire [31:0] p2_add_93019_comb;
  wire [31:0] p2_add_93020_comb;
  wire [31:0] p2_add_92663_comb;
  wire [31:0] p2_add_92664_comb;
  wire [31:0] p2_add_93015_comb;
  wire [31:0] p2_add_93016_comb;
  wire [31:0] p2_add_92661_comb;
  wire [31:0] p2_add_92662_comb;
  wire [31:0] p2_add_93011_comb;
  wire [31:0] p2_add_93012_comb;
  wire [31:0] p2_add_92659_comb;
  wire [31:0] p2_add_92660_comb;
  wire [31:0] p2_add_93007_comb;
  wire [31:0] p2_add_93008_comb;
  wire [31:0] p2_add_92657_comb;
  wire [31:0] p2_add_92658_comb;
  wire [31:0] p2_add_93003_comb;
  wire [31:0] p2_add_93004_comb;
  wire [31:0] p2_add_92655_comb;
  wire [31:0] p2_add_92656_comb;
  wire [31:0] p2_add_92999_comb;
  wire [31:0] p2_add_93000_comb;
  wire [31:0] p2_add_92653_comb;
  wire [31:0] p2_add_92654_comb;
  wire [31:0] p2_add_92995_comb;
  wire [31:0] p2_add_92996_comb;
  wire [31:0] p2_add_92651_comb;
  wire [31:0] p2_add_92652_comb;
  wire [31:0] p2_add_92991_comb;
  wire [31:0] p2_add_92992_comb;
  wire [31:0] p2_add_92649_comb;
  wire [31:0] p2_add_92650_comb;
  wire [31:0] p2_add_92987_comb;
  wire [31:0] p2_add_92988_comb;
  wire [31:0] p2_add_92647_comb;
  wire [31:0] p2_add_92648_comb;
  wire [31:0] p2_add_92983_comb;
  wire [31:0] p2_add_92984_comb;
  wire [31:0] p2_add_92645_comb;
  wire [31:0] p2_add_92646_comb;
  wire [31:0] p2_add_92979_comb;
  wire [31:0] p2_add_92980_comb;
  wire [31:0] p2_add_92643_comb;
  wire [31:0] p2_add_92644_comb;
  wire [31:0] p2_add_92975_comb;
  wire [31:0] p2_add_92976_comb;
  wire [31:0] p2_add_92641_comb;
  wire [31:0] p2_add_92642_comb;
  wire [31:0] p2_add_92971_comb;
  wire [31:0] p2_add_92972_comb;
  wire [31:0] p2_add_92639_comb;
  wire [31:0] p2_add_92640_comb;
  wire [31:0] p2_add_92967_comb;
  wire [31:0] p2_add_92968_comb;
  wire [31:0] p2_add_92637_comb;
  wire [31:0] p2_add_92638_comb;
  wire [31:0] p2_add_92963_comb;
  wire [31:0] p2_add_92964_comb;
  wire [31:0] p2_add_92635_comb;
  wire [31:0] p2_add_92636_comb;
  wire [31:0] p2_add_92959_comb;
  wire [31:0] p2_add_92960_comb;
  wire [31:0] p2_add_92633_comb;
  wire [31:0] p2_add_92634_comb;
  wire [31:0] p2_add_92955_comb;
  wire [31:0] p2_add_92956_comb;
  wire [31:0] p2_add_92631_comb;
  wire [31:0] p2_add_92632_comb;
  wire [31:0] p2_add_92951_comb;
  wire [31:0] p2_add_92952_comb;
  wire [31:0] p2_add_92629_comb;
  wire [31:0] p2_add_92630_comb;
  wire [31:0] p2_add_92947_comb;
  wire [31:0] p2_add_92948_comb;
  wire [31:0] p2_add_92627_comb;
  wire [31:0] p2_add_92628_comb;
  wire [31:0] p2_add_92943_comb;
  wire [31:0] p2_add_92944_comb;
  wire [31:0] p2_add_92625_comb;
  wire [31:0] p2_add_92626_comb;
  wire [31:0] p2_add_92939_comb;
  wire [31:0] p2_add_92940_comb;
  wire [31:0] p2_add_92623_comb;
  wire [31:0] p2_add_92624_comb;
  wire [31:0] p2_add_92935_comb;
  wire [31:0] p2_add_92936_comb;
  wire [31:0] p2_add_92621_comb;
  wire [31:0] p2_add_92622_comb;
  wire [31:0] p2_add_92931_comb;
  wire [31:0] p2_add_92932_comb;
  wire [31:0] p2_add_92619_comb;
  wire [31:0] p2_add_92620_comb;
  wire [31:0] p2_add_92927_comb;
  wire [31:0] p2_add_92928_comb;
  wire [31:0] p2_add_92617_comb;
  wire [31:0] p2_add_92618_comb;
  wire [31:0] p2_add_92923_comb;
  wire [31:0] p2_add_92924_comb;
  wire [31:0] p2_add_92615_comb;
  wire [31:0] p2_add_92616_comb;
  wire [31:0] p2_add_92919_comb;
  wire [31:0] p2_add_92920_comb;
  wire [31:0] p2_add_92613_comb;
  wire [31:0] p2_add_92614_comb;
  wire [31:0] p2_add_92915_comb;
  wire [31:0] p2_add_92916_comb;
  wire [31:0] p2_add_92611_comb;
  wire [31:0] p2_add_92612_comb;
  wire [31:0] p2_add_92911_comb;
  wire [31:0] p2_add_92912_comb;
  wire [31:0] p2_add_92609_comb;
  wire [31:0] p2_add_92610_comb;
  wire [31:0] p2_add_92907_comb;
  wire [31:0] p2_add_92908_comb;
  wire [31:0] p2_add_92607_comb;
  wire [31:0] p2_add_92608_comb;
  wire [31:0] p2_add_92903_comb;
  wire [31:0] p2_add_92904_comb;
  wire [31:0] p2_add_92605_comb;
  wire [31:0] p2_add_92606_comb;
  wire [31:0] p2_add_92899_comb;
  wire [31:0] p2_add_92900_comb;
  wire [31:0] p2_add_92603_comb;
  wire [31:0] p2_add_92604_comb;
  wire [31:0] p2_add_92895_comb;
  wire [31:0] p2_add_92896_comb;
  wire [31:0] p2_add_92601_comb;
  wire [31:0] p2_add_92602_comb;
  wire [31:0] p2_add_92891_comb;
  wire [31:0] p2_add_92892_comb;
  wire [31:0] p2_add_92599_comb;
  wire [31:0] p2_add_92600_comb;
  wire [31:0] p2_add_92887_comb;
  wire [31:0] p2_add_92888_comb;
  wire [31:0] p2_add_92597_comb;
  wire [31:0] p2_add_92598_comb;
  wire [31:0] p2_add_92883_comb;
  wire [31:0] p2_add_92884_comb;
  wire [31:0] p2_add_92595_comb;
  wire [31:0] p2_add_92596_comb;
  wire [31:0] p2_add_92879_comb;
  wire [31:0] p2_add_92880_comb;
  wire [31:0] p2_add_92593_comb;
  wire [31:0] p2_add_92594_comb;
  wire [31:0] p2_add_92875_comb;
  wire [31:0] p2_add_92876_comb;
  wire [31:0] p2_add_92591_comb;
  wire [31:0] p2_add_92592_comb;
  wire [31:0] p2_add_92871_comb;
  wire [31:0] p2_add_92872_comb;
  wire [31:0] p2_add_92589_comb;
  wire [31:0] p2_add_92590_comb;
  wire [31:0] p2_add_92867_comb;
  wire [31:0] p2_add_92868_comb;
  wire [31:0] p2_add_92587_comb;
  wire [31:0] p2_add_92588_comb;
  wire [31:0] p2_add_92863_comb;
  wire [31:0] p2_add_92864_comb;
  wire [31:0] p2_add_92585_comb;
  wire [31:0] p2_add_92586_comb;
  wire [31:0] p2_add_92859_comb;
  wire [31:0] p2_add_92860_comb;
  wire [31:0] p2_add_92583_comb;
  wire [31:0] p2_add_92584_comb;
  wire [31:0] p2_add_92855_comb;
  wire [31:0] p2_add_92856_comb;
  wire [31:0] p2_add_92581_comb;
  wire [31:0] p2_add_92582_comb;
  wire [31:0] p2_add_92851_comb;
  wire [31:0] p2_add_92852_comb;
  wire [31:0] p2_add_92579_comb;
  wire [31:0] p2_add_92580_comb;
  wire [31:0] p2_add_92847_comb;
  wire [31:0] p2_add_92848_comb;
  wire [31:0] p2_add_92577_comb;
  wire [31:0] p2_add_92578_comb;
  wire [31:0] p2_add_92843_comb;
  wire [31:0] p2_add_92844_comb;
  wire [31:0] p2_add_92575_comb;
  wire [31:0] p2_add_92576_comb;
  wire [31:0] p2_add_92839_comb;
  wire [31:0] p2_add_92840_comb;
  wire [31:0] p2_add_92573_comb;
  wire [31:0] p2_add_92574_comb;
  wire [31:0] p2_add_92835_comb;
  wire [31:0] p2_add_92836_comb;
  wire [31:0] p2_add_92571_comb;
  wire [31:0] p2_add_92572_comb;
  wire [31:0] p2_add_92831_comb;
  wire [31:0] p2_add_92832_comb;
  wire [31:0] p2_add_92569_comb;
  wire [31:0] p2_add_92570_comb;
  wire [31:0] p2_add_92827_comb;
  wire [31:0] p2_add_92828_comb;
  wire [31:0] p2_add_92567_comb;
  wire [31:0] p2_add_92568_comb;
  wire [31:0] p2_add_92823_comb;
  wire [31:0] p2_add_92824_comb;
  wire [31:0] p2_add_92565_comb;
  wire [31:0] p2_add_92566_comb;
  wire [31:0] p2_add_92819_comb;
  wire [31:0] p2_add_92820_comb;
  wire [31:0] p2_add_92563_comb;
  wire [31:0] p2_add_92564_comb;
  wire [31:0] p2_add_92815_comb;
  wire [31:0] p2_add_92816_comb;
  wire [31:0] p2_add_92561_comb;
  wire [31:0] p2_add_92562_comb;
  wire [31:0] p2_add_92811_comb;
  wire [31:0] p2_add_92812_comb;
  wire [31:0] p2_add_92559_comb;
  wire [31:0] p2_add_92560_comb;
  wire [31:0] p2_add_92807_comb;
  wire [31:0] p2_add_92808_comb;
  wire [31:0] p2_add_92557_comb;
  wire [31:0] p2_add_92558_comb;
  wire [31:0] p2_add_92803_comb;
  wire [31:0] p2_add_92804_comb;
  wire [31:0] p2_add_92555_comb;
  wire [31:0] p2_add_92556_comb;
  wire [31:0] p2_add_92799_comb;
  wire [31:0] p2_add_92800_comb;
  wire [31:0] p2_add_92553_comb;
  wire [31:0] p2_add_92554_comb;
  wire [31:0] p2_add_92795_comb;
  wire [31:0] p2_add_92796_comb;
  wire [31:0] p2_add_92551_comb;
  wire [31:0] p2_add_92552_comb;
  wire [31:0] p2_add_92791_comb;
  wire [31:0] p2_add_92792_comb;
  wire [31:0] p2_add_92549_comb;
  wire [31:0] p2_add_92550_comb;
  wire [31:0] p2_add_92787_comb;
  wire [31:0] p2_add_92788_comb;
  wire [31:0] p2_add_92547_comb;
  wire [31:0] p2_add_92548_comb;
  wire [31:0] p2_add_92783_comb;
  wire [31:0] p2_add_92784_comb;
  wire [31:0] p2_add_92545_comb;
  wire [31:0] p2_add_92546_comb;
  wire [31:0] p2_add_92779_comb;
  wire [31:0] p2_add_92780_comb;
  wire [31:0] p2_add_92543_comb;
  wire [31:0] p2_add_92544_comb;
  wire [31:0] p2_add_92775_comb;
  wire [31:0] p2_add_92776_comb;
  wire [31:0] p2_add_92541_comb;
  wire [31:0] p2_add_92542_comb;
  wire [31:0] p2_add_92771_comb;
  wire [31:0] p2_add_92772_comb;
  wire [31:0] p2_add_92539_comb;
  wire [31:0] p2_add_92540_comb;
  wire [31:0] p2_add_92767_comb;
  wire [31:0] p2_add_92768_comb;
  wire [31:0] p2_add_92537_comb;
  wire [31:0] p2_add_92538_comb;
  wire [31:0] p2_add_92763_comb;
  wire [31:0] p2_add_92764_comb;
  wire [31:0] p2_add_92535_comb;
  wire [31:0] p2_add_92536_comb;
  wire [31:0] p2_add_92759_comb;
  wire [31:0] p2_add_92760_comb;
  wire [31:0] p2_add_92533_comb;
  wire [31:0] p2_add_92534_comb;
  wire [31:0] p2_add_92755_comb;
  wire [31:0] p2_add_92756_comb;
  wire [31:0] p2_add_92531_comb;
  wire [31:0] p2_add_92532_comb;
  wire [31:0] p2_add_92751_comb;
  wire [31:0] p2_add_92752_comb;
  wire [31:0] p2_add_92529_comb;
  wire [31:0] p2_add_92530_comb;
  wire [31:0] p2_add_92747_comb;
  wire [31:0] p2_add_92748_comb;
  wire [31:0] p2_add_92527_comb;
  wire [31:0] p2_add_92528_comb;
  wire [31:0] p2_add_92743_comb;
  wire [31:0] p2_add_92744_comb;
  wire [31:0] p2_add_92525_comb;
  wire [31:0] p2_add_92526_comb;
  wire [31:0] p2_add_92739_comb;
  wire [31:0] p2_add_92740_comb;
  wire [31:0] p2_add_92523_comb;
  wire [31:0] p2_add_92524_comb;
  wire [31:0] p2_add_92735_comb;
  wire [31:0] p2_add_92736_comb;
  wire [31:0] p2_add_92521_comb;
  wire [31:0] p2_add_92522_comb;
  wire [31:0] p2_add_92731_comb;
  wire [31:0] p2_add_92732_comb;
  wire [31:0] p2_add_92519_comb;
  wire [31:0] p2_add_92520_comb;
  wire [31:0] p2_add_92727_comb;
  wire [31:0] p2_add_92728_comb;
  wire [31:0] p2_add_92517_comb;
  wire [31:0] p2_add_92518_comb;
  wire [31:0] p2_add_92723_comb;
  wire [31:0] p2_add_92724_comb;
  wire [31:0] p2_add_92515_comb;
  wire [31:0] p2_add_92516_comb;
  wire [31:0] p2_add_92719_comb;
  wire [31:0] p2_add_92720_comb;
  wire [31:0] p2_add_92513_comb;
  wire [31:0] p2_add_92514_comb;
  wire [31:0] p2_add_92715_comb;
  wire [31:0] p2_add_92716_comb;
  wire [31:0] p2_add_93109_comb;
  wire [31:0] p2_add_93110_comb;
  wire [31:0] p2_add_93212_comb;
  wire [31:0] p2_add_93105_comb;
  wire [31:0] p2_add_93106_comb;
  wire [31:0] p2_add_93211_comb;
  wire [31:0] p2_add_93101_comb;
  wire [31:0] p2_add_93102_comb;
  wire [31:0] p2_add_93210_comb;
  wire [31:0] p2_add_93097_comb;
  wire [31:0] p2_add_93098_comb;
  wire [31:0] p2_add_93209_comb;
  wire [31:0] p2_add_93093_comb;
  wire [31:0] p2_add_93094_comb;
  wire [31:0] p2_add_93208_comb;
  wire [31:0] p2_add_93089_comb;
  wire [31:0] p2_add_93090_comb;
  wire [31:0] p2_add_93207_comb;
  wire [31:0] p2_add_93085_comb;
  wire [31:0] p2_add_93086_comb;
  wire [31:0] p2_add_93206_comb;
  wire [31:0] p2_add_93081_comb;
  wire [31:0] p2_add_93082_comb;
  wire [31:0] p2_add_93205_comb;
  wire [31:0] p2_add_93077_comb;
  wire [31:0] p2_add_93078_comb;
  wire [31:0] p2_add_93204_comb;
  wire [31:0] p2_add_93073_comb;
  wire [31:0] p2_add_93074_comb;
  wire [31:0] p2_add_93203_comb;
  wire [31:0] p2_add_93069_comb;
  wire [31:0] p2_add_93070_comb;
  wire [31:0] p2_add_93202_comb;
  wire [31:0] p2_add_93065_comb;
  wire [31:0] p2_add_93066_comb;
  wire [31:0] p2_add_93201_comb;
  wire [31:0] p2_add_93061_comb;
  wire [31:0] p2_add_93062_comb;
  wire [31:0] p2_add_93200_comb;
  wire [31:0] p2_add_93057_comb;
  wire [31:0] p2_add_93058_comb;
  wire [31:0] p2_add_93199_comb;
  wire [31:0] p2_add_93053_comb;
  wire [31:0] p2_add_93054_comb;
  wire [31:0] p2_add_93198_comb;
  wire [31:0] p2_add_93049_comb;
  wire [31:0] p2_add_93050_comb;
  wire [31:0] p2_add_93197_comb;
  wire [31:0] p2_add_93045_comb;
  wire [31:0] p2_add_93046_comb;
  wire [31:0] p2_add_93196_comb;
  wire [31:0] p2_add_93041_comb;
  wire [31:0] p2_add_93042_comb;
  wire [31:0] p2_add_93195_comb;
  wire [31:0] p2_add_93037_comb;
  wire [31:0] p2_add_93038_comb;
  wire [31:0] p2_add_93194_comb;
  wire [31:0] p2_add_93033_comb;
  wire [31:0] p2_add_93034_comb;
  wire [31:0] p2_add_93193_comb;
  wire [31:0] p2_add_93029_comb;
  wire [31:0] p2_add_93030_comb;
  wire [31:0] p2_add_93192_comb;
  wire [31:0] p2_add_93025_comb;
  wire [31:0] p2_add_93026_comb;
  wire [31:0] p2_add_93191_comb;
  wire [31:0] p2_add_93021_comb;
  wire [31:0] p2_add_93022_comb;
  wire [31:0] p2_add_93190_comb;
  wire [31:0] p2_add_93017_comb;
  wire [31:0] p2_add_93018_comb;
  wire [31:0] p2_add_93189_comb;
  wire [31:0] p2_add_93013_comb;
  wire [31:0] p2_add_93014_comb;
  wire [31:0] p2_add_93188_comb;
  wire [31:0] p2_add_93009_comb;
  wire [31:0] p2_add_93010_comb;
  wire [31:0] p2_add_93187_comb;
  wire [31:0] p2_add_93005_comb;
  wire [31:0] p2_add_93006_comb;
  wire [31:0] p2_add_93186_comb;
  wire [31:0] p2_add_93001_comb;
  wire [31:0] p2_add_93002_comb;
  wire [31:0] p2_add_93185_comb;
  wire [31:0] p2_add_92997_comb;
  wire [31:0] p2_add_92998_comb;
  wire [31:0] p2_add_93184_comb;
  wire [31:0] p2_add_92993_comb;
  wire [31:0] p2_add_92994_comb;
  wire [31:0] p2_add_93183_comb;
  wire [31:0] p2_add_92989_comb;
  wire [31:0] p2_add_92990_comb;
  wire [31:0] p2_add_93182_comb;
  wire [31:0] p2_add_92985_comb;
  wire [31:0] p2_add_92986_comb;
  wire [31:0] p2_add_93181_comb;
  wire [31:0] p2_add_92981_comb;
  wire [31:0] p2_add_92982_comb;
  wire [31:0] p2_add_93180_comb;
  wire [31:0] p2_add_92977_comb;
  wire [31:0] p2_add_92978_comb;
  wire [31:0] p2_add_93179_comb;
  wire [31:0] p2_add_92973_comb;
  wire [31:0] p2_add_92974_comb;
  wire [31:0] p2_add_93178_comb;
  wire [31:0] p2_add_92969_comb;
  wire [31:0] p2_add_92970_comb;
  wire [31:0] p2_add_93177_comb;
  wire [31:0] p2_add_92965_comb;
  wire [31:0] p2_add_92966_comb;
  wire [31:0] p2_add_93176_comb;
  wire [31:0] p2_add_92961_comb;
  wire [31:0] p2_add_92962_comb;
  wire [31:0] p2_add_93175_comb;
  wire [31:0] p2_add_92957_comb;
  wire [31:0] p2_add_92958_comb;
  wire [31:0] p2_add_93174_comb;
  wire [31:0] p2_add_92953_comb;
  wire [31:0] p2_add_92954_comb;
  wire [31:0] p2_add_93173_comb;
  wire [31:0] p2_add_92949_comb;
  wire [31:0] p2_add_92950_comb;
  wire [31:0] p2_add_93172_comb;
  wire [31:0] p2_add_92945_comb;
  wire [31:0] p2_add_92946_comb;
  wire [31:0] p2_add_93171_comb;
  wire [31:0] p2_add_92941_comb;
  wire [31:0] p2_add_92942_comb;
  wire [31:0] p2_add_93170_comb;
  wire [31:0] p2_add_92937_comb;
  wire [31:0] p2_add_92938_comb;
  wire [31:0] p2_add_93169_comb;
  wire [31:0] p2_add_92933_comb;
  wire [31:0] p2_add_92934_comb;
  wire [31:0] p2_add_93168_comb;
  wire [31:0] p2_add_92929_comb;
  wire [31:0] p2_add_92930_comb;
  wire [31:0] p2_add_93167_comb;
  wire [31:0] p2_add_92925_comb;
  wire [31:0] p2_add_92926_comb;
  wire [31:0] p2_add_93166_comb;
  wire [31:0] p2_add_92921_comb;
  wire [31:0] p2_add_92922_comb;
  wire [31:0] p2_add_93165_comb;
  wire [31:0] p2_add_92917_comb;
  wire [31:0] p2_add_92918_comb;
  wire [31:0] p2_add_93164_comb;
  wire [31:0] p2_add_92913_comb;
  wire [31:0] p2_add_92914_comb;
  wire [31:0] p2_add_93163_comb;
  wire [31:0] p2_add_92909_comb;
  wire [31:0] p2_add_92910_comb;
  wire [31:0] p2_add_93162_comb;
  wire [31:0] p2_add_92905_comb;
  wire [31:0] p2_add_92906_comb;
  wire [31:0] p2_add_93161_comb;
  wire [31:0] p2_add_92901_comb;
  wire [31:0] p2_add_92902_comb;
  wire [31:0] p2_add_93160_comb;
  wire [31:0] p2_add_92897_comb;
  wire [31:0] p2_add_92898_comb;
  wire [31:0] p2_add_93159_comb;
  wire [31:0] p2_add_92893_comb;
  wire [31:0] p2_add_92894_comb;
  wire [31:0] p2_add_93158_comb;
  wire [31:0] p2_add_92889_comb;
  wire [31:0] p2_add_92890_comb;
  wire [31:0] p2_add_93157_comb;
  wire [31:0] p2_add_92885_comb;
  wire [31:0] p2_add_92886_comb;
  wire [31:0] p2_add_93156_comb;
  wire [31:0] p2_add_92881_comb;
  wire [31:0] p2_add_92882_comb;
  wire [31:0] p2_add_93155_comb;
  wire [31:0] p2_add_92877_comb;
  wire [31:0] p2_add_92878_comb;
  wire [31:0] p2_add_93154_comb;
  wire [31:0] p2_add_92873_comb;
  wire [31:0] p2_add_92874_comb;
  wire [31:0] p2_add_93153_comb;
  wire [31:0] p2_add_92869_comb;
  wire [31:0] p2_add_92870_comb;
  wire [31:0] p2_add_93152_comb;
  wire [31:0] p2_add_92865_comb;
  wire [31:0] p2_add_92866_comb;
  wire [31:0] p2_add_93151_comb;
  wire [31:0] p2_add_92861_comb;
  wire [31:0] p2_add_92862_comb;
  wire [31:0] p2_add_93150_comb;
  wire [31:0] p2_add_92857_comb;
  wire [31:0] p2_add_92858_comb;
  wire [31:0] p2_add_93149_comb;
  wire [31:0] p2_add_92853_comb;
  wire [31:0] p2_add_92854_comb;
  wire [31:0] p2_add_93148_comb;
  wire [31:0] p2_add_92849_comb;
  wire [31:0] p2_add_92850_comb;
  wire [31:0] p2_add_93147_comb;
  wire [31:0] p2_add_92845_comb;
  wire [31:0] p2_add_92846_comb;
  wire [31:0] p2_add_93146_comb;
  wire [31:0] p2_add_92841_comb;
  wire [31:0] p2_add_92842_comb;
  wire [31:0] p2_add_93145_comb;
  wire [31:0] p2_add_92837_comb;
  wire [31:0] p2_add_92838_comb;
  wire [31:0] p2_add_93144_comb;
  wire [31:0] p2_add_92833_comb;
  wire [31:0] p2_add_92834_comb;
  wire [31:0] p2_add_93143_comb;
  wire [31:0] p2_add_92829_comb;
  wire [31:0] p2_add_92830_comb;
  wire [31:0] p2_add_93142_comb;
  wire [31:0] p2_add_92825_comb;
  wire [31:0] p2_add_92826_comb;
  wire [31:0] p2_add_93141_comb;
  wire [31:0] p2_add_92821_comb;
  wire [31:0] p2_add_92822_comb;
  wire [31:0] p2_add_93140_comb;
  wire [31:0] p2_add_92817_comb;
  wire [31:0] p2_add_92818_comb;
  wire [31:0] p2_add_93139_comb;
  wire [31:0] p2_add_92813_comb;
  wire [31:0] p2_add_92814_comb;
  wire [31:0] p2_add_93138_comb;
  wire [31:0] p2_add_92809_comb;
  wire [31:0] p2_add_92810_comb;
  wire [31:0] p2_add_93137_comb;
  wire [31:0] p2_add_92805_comb;
  wire [31:0] p2_add_92806_comb;
  wire [31:0] p2_add_93136_comb;
  wire [31:0] p2_add_92801_comb;
  wire [31:0] p2_add_92802_comb;
  wire [31:0] p2_add_93135_comb;
  wire [31:0] p2_add_92797_comb;
  wire [31:0] p2_add_92798_comb;
  wire [31:0] p2_add_93134_comb;
  wire [31:0] p2_add_92793_comb;
  wire [31:0] p2_add_92794_comb;
  wire [31:0] p2_add_93133_comb;
  wire [31:0] p2_add_92789_comb;
  wire [31:0] p2_add_92790_comb;
  wire [31:0] p2_add_93132_comb;
  wire [31:0] p2_add_92785_comb;
  wire [31:0] p2_add_92786_comb;
  wire [31:0] p2_add_93131_comb;
  wire [31:0] p2_add_92781_comb;
  wire [31:0] p2_add_92782_comb;
  wire [31:0] p2_add_93130_comb;
  wire [31:0] p2_add_92777_comb;
  wire [31:0] p2_add_92778_comb;
  wire [31:0] p2_add_93129_comb;
  wire [31:0] p2_add_92773_comb;
  wire [31:0] p2_add_92774_comb;
  wire [31:0] p2_add_93128_comb;
  wire [31:0] p2_add_92769_comb;
  wire [31:0] p2_add_92770_comb;
  wire [31:0] p2_add_93127_comb;
  wire [31:0] p2_add_92765_comb;
  wire [31:0] p2_add_92766_comb;
  wire [31:0] p2_add_93126_comb;
  wire [31:0] p2_add_92761_comb;
  wire [31:0] p2_add_92762_comb;
  wire [31:0] p2_add_93125_comb;
  wire [31:0] p2_add_92757_comb;
  wire [31:0] p2_add_92758_comb;
  wire [31:0] p2_add_93124_comb;
  wire [31:0] p2_add_92753_comb;
  wire [31:0] p2_add_92754_comb;
  wire [31:0] p2_add_93123_comb;
  wire [31:0] p2_add_92749_comb;
  wire [31:0] p2_add_92750_comb;
  wire [31:0] p2_add_93122_comb;
  wire [31:0] p2_add_92745_comb;
  wire [31:0] p2_add_92746_comb;
  wire [31:0] p2_add_93121_comb;
  wire [31:0] p2_add_92741_comb;
  wire [31:0] p2_add_92742_comb;
  wire [31:0] p2_add_93120_comb;
  wire [31:0] p2_add_92737_comb;
  wire [31:0] p2_add_92738_comb;
  wire [31:0] p2_add_93119_comb;
  wire [31:0] p2_add_92733_comb;
  wire [31:0] p2_add_92734_comb;
  wire [31:0] p2_add_93118_comb;
  wire [31:0] p2_add_92729_comb;
  wire [31:0] p2_add_92730_comb;
  wire [31:0] p2_add_93117_comb;
  wire [31:0] p2_add_92725_comb;
  wire [31:0] p2_add_92726_comb;
  wire [31:0] p2_add_93116_comb;
  wire [31:0] p2_add_92721_comb;
  wire [31:0] p2_add_92722_comb;
  wire [31:0] p2_add_93115_comb;
  wire [31:0] p2_add_92717_comb;
  wire [31:0] p2_add_92718_comb;
  wire [31:0] p2_add_93114_comb;
  wire [31:0] p2_add_92713_comb;
  wire [31:0] p2_add_92714_comb;
  wire [31:0] p2_add_93113_comb;
  assign p2_add_92711_comb = p1_smul_89895 + p1_smul_89896;
  assign p2_add_92712_comb = p1_smul_89897 + p1_smul_89898;
  assign p2_add_93111_comb = p1_smul_90495 + p1_smul_90496;
  assign p2_add_93112_comb = p1_smul_90497 + p1_smul_90498;
  assign p2_add_92709_comb = p1_smul_89891 + p1_smul_89892;
  assign p2_add_92710_comb = p1_smul_89893 + p1_smul_89894;
  assign p2_add_93107_comb = p1_smul_90489 + p1_smul_90490;
  assign p2_add_93108_comb = p1_smul_90491 + p1_smul_90492;
  assign p2_add_92707_comb = p1_smul_89887 + p1_smul_89888;
  assign p2_add_92708_comb = p1_smul_89889 + p1_smul_89890;
  assign p2_add_93103_comb = p1_smul_90483 + p1_smul_90484;
  assign p2_add_93104_comb = p1_smul_90485 + p1_smul_90486;
  assign p2_add_92705_comb = p1_smul_89883 + p1_smul_89884;
  assign p2_add_92706_comb = p1_smul_89885 + p1_smul_89886;
  assign p2_add_93099_comb = p1_smul_90477 + p1_smul_90478;
  assign p2_add_93100_comb = p1_smul_90479 + p1_smul_90480;
  assign p2_add_92703_comb = p1_smul_89879 + p1_smul_89880;
  assign p2_add_92704_comb = p1_smul_89881 + p1_smul_89882;
  assign p2_add_93095_comb = p1_smul_90471 + p1_smul_90472;
  assign p2_add_93096_comb = p1_smul_90473 + p1_smul_90474;
  assign p2_add_92701_comb = p1_smul_89875 + p1_smul_89876;
  assign p2_add_92702_comb = p1_smul_89877 + p1_smul_89878;
  assign p2_add_93091_comb = p1_smul_90465 + p1_smul_90466;
  assign p2_add_93092_comb = p1_smul_90467 + p1_smul_90468;
  assign p2_add_92699_comb = p1_smul_89871 + p1_smul_89872;
  assign p2_add_92700_comb = p1_smul_89873 + p1_smul_89874;
  assign p2_add_93087_comb = p1_smul_90459 + p1_smul_90460;
  assign p2_add_93088_comb = p1_smul_90461 + p1_smul_90462;
  assign p2_add_92697_comb = p1_smul_89867 + p1_smul_89868;
  assign p2_add_92698_comb = p1_smul_89869 + p1_smul_89870;
  assign p2_add_93083_comb = p1_smul_90453 + p1_smul_90454;
  assign p2_add_93084_comb = p1_smul_90455 + p1_smul_90456;
  assign p2_add_92695_comb = p1_smul_89863 + p1_smul_89864;
  assign p2_add_92696_comb = p1_smul_89865 + p1_smul_89866;
  assign p2_add_93079_comb = p1_smul_90447 + p1_smul_90448;
  assign p2_add_93080_comb = p1_smul_90449 + p1_smul_90450;
  assign p2_add_92693_comb = p1_smul_89859 + p1_smul_89860;
  assign p2_add_92694_comb = p1_smul_89861 + p1_smul_89862;
  assign p2_add_93075_comb = p1_smul_90441 + p1_smul_90442;
  assign p2_add_93076_comb = p1_smul_90443 + p1_smul_90444;
  assign p2_add_92691_comb = p1_smul_89855 + p1_smul_89856;
  assign p2_add_92692_comb = p1_smul_89857 + p1_smul_89858;
  assign p2_add_93071_comb = p1_smul_90435 + p1_smul_90436;
  assign p2_add_93072_comb = p1_smul_90437 + p1_smul_90438;
  assign p2_add_92689_comb = p1_smul_89851 + p1_smul_89852;
  assign p2_add_92690_comb = p1_smul_89853 + p1_smul_89854;
  assign p2_add_93067_comb = p1_smul_90429 + p1_smul_90430;
  assign p2_add_93068_comb = p1_smul_90431 + p1_smul_90432;
  assign p2_add_92687_comb = p1_smul_89847 + p1_smul_89848;
  assign p2_add_92688_comb = p1_smul_89849 + p1_smul_89850;
  assign p2_add_93063_comb = p1_smul_90423 + p1_smul_90424;
  assign p2_add_93064_comb = p1_smul_90425 + p1_smul_90426;
  assign p2_add_92685_comb = p1_smul_89843 + p1_smul_89844;
  assign p2_add_92686_comb = p1_smul_89845 + p1_smul_89846;
  assign p2_add_93059_comb = p1_smul_90417 + p1_smul_90418;
  assign p2_add_93060_comb = p1_smul_90419 + p1_smul_90420;
  assign p2_add_92683_comb = p1_smul_89839 + p1_smul_89840;
  assign p2_add_92684_comb = p1_smul_89841 + p1_smul_89842;
  assign p2_add_93055_comb = p1_smul_90411 + p1_smul_90412;
  assign p2_add_93056_comb = p1_smul_90413 + p1_smul_90414;
  assign p2_add_92681_comb = p1_smul_89835 + p1_smul_89836;
  assign p2_add_92682_comb = p1_smul_89837 + p1_smul_89838;
  assign p2_add_93051_comb = p1_smul_90405 + p1_smul_90406;
  assign p2_add_93052_comb = p1_smul_90407 + p1_smul_90408;
  assign p2_add_92679_comb = p1_smul_89831 + p1_smul_89832;
  assign p2_add_92680_comb = p1_smul_89833 + p1_smul_89834;
  assign p2_add_93047_comb = p1_smul_90399 + p1_smul_90400;
  assign p2_add_93048_comb = p1_smul_90401 + p1_smul_90402;
  assign p2_add_92677_comb = p1_smul_89827 + p1_smul_89828;
  assign p2_add_92678_comb = p1_smul_89829 + p1_smul_89830;
  assign p2_add_93043_comb = p1_smul_90393 + p1_smul_90394;
  assign p2_add_93044_comb = p1_smul_90395 + p1_smul_90396;
  assign p2_add_92675_comb = p1_smul_89823 + p1_smul_89824;
  assign p2_add_92676_comb = p1_smul_89825 + p1_smul_89826;
  assign p2_add_93039_comb = p1_smul_90387 + p1_smul_90388;
  assign p2_add_93040_comb = p1_smul_90389 + p1_smul_90390;
  assign p2_add_92673_comb = p1_smul_89819 + p1_smul_89820;
  assign p2_add_92674_comb = p1_smul_89821 + p1_smul_89822;
  assign p2_add_93035_comb = p1_smul_90381 + p1_smul_90382;
  assign p2_add_93036_comb = p1_smul_90383 + p1_smul_90384;
  assign p2_add_92671_comb = p1_smul_89815 + p1_smul_89816;
  assign p2_add_92672_comb = p1_smul_89817 + p1_smul_89818;
  assign p2_add_93031_comb = p1_smul_90375 + p1_smul_90376;
  assign p2_add_93032_comb = p1_smul_90377 + p1_smul_90378;
  assign p2_add_92669_comb = p1_smul_89811 + p1_smul_89812;
  assign p2_add_92670_comb = p1_smul_89813 + p1_smul_89814;
  assign p2_add_93027_comb = p1_smul_90369 + p1_smul_90370;
  assign p2_add_93028_comb = p1_smul_90371 + p1_smul_90372;
  assign p2_add_92667_comb = p1_smul_89807 + p1_smul_89808;
  assign p2_add_92668_comb = p1_smul_89809 + p1_smul_89810;
  assign p2_add_93023_comb = p1_smul_90363 + p1_smul_90364;
  assign p2_add_93024_comb = p1_smul_90365 + p1_smul_90366;
  assign p2_add_92665_comb = p1_smul_89803 + p1_smul_89804;
  assign p2_add_92666_comb = p1_smul_89805 + p1_smul_89806;
  assign p2_add_93019_comb = p1_smul_90357 + p1_smul_90358;
  assign p2_add_93020_comb = p1_smul_90359 + p1_smul_90360;
  assign p2_add_92663_comb = p1_smul_89799 + p1_smul_89800;
  assign p2_add_92664_comb = p1_smul_89801 + p1_smul_89802;
  assign p2_add_93015_comb = p1_smul_90351 + p1_smul_90352;
  assign p2_add_93016_comb = p1_smul_90353 + p1_smul_90354;
  assign p2_add_92661_comb = p1_smul_89795 + p1_smul_89796;
  assign p2_add_92662_comb = p1_smul_89797 + p1_smul_89798;
  assign p2_add_93011_comb = p1_smul_90345 + p1_smul_90346;
  assign p2_add_93012_comb = p1_smul_90347 + p1_smul_90348;
  assign p2_add_92659_comb = p1_smul_89791 + p1_smul_89792;
  assign p2_add_92660_comb = p1_smul_89793 + p1_smul_89794;
  assign p2_add_93007_comb = p1_smul_90339 + p1_smul_90340;
  assign p2_add_93008_comb = p1_smul_90341 + p1_smul_90342;
  assign p2_add_92657_comb = p1_smul_89787 + p1_smul_89788;
  assign p2_add_92658_comb = p1_smul_89789 + p1_smul_89790;
  assign p2_add_93003_comb = p1_smul_90333 + p1_smul_90334;
  assign p2_add_93004_comb = p1_smul_90335 + p1_smul_90336;
  assign p2_add_92655_comb = p1_smul_89783 + p1_smul_89784;
  assign p2_add_92656_comb = p1_smul_89785 + p1_smul_89786;
  assign p2_add_92999_comb = p1_smul_90327 + p1_smul_90328;
  assign p2_add_93000_comb = p1_smul_90329 + p1_smul_90330;
  assign p2_add_92653_comb = p1_smul_89779 + p1_smul_89780;
  assign p2_add_92654_comb = p1_smul_89781 + p1_smul_89782;
  assign p2_add_92995_comb = p1_smul_90321 + p1_smul_90322;
  assign p2_add_92996_comb = p1_smul_90323 + p1_smul_90324;
  assign p2_add_92651_comb = p1_smul_89775 + p1_smul_89776;
  assign p2_add_92652_comb = p1_smul_89777 + p1_smul_89778;
  assign p2_add_92991_comb = p1_smul_90315 + p1_smul_90316;
  assign p2_add_92992_comb = p1_smul_90317 + p1_smul_90318;
  assign p2_add_92649_comb = p1_smul_89771 + p1_smul_89772;
  assign p2_add_92650_comb = p1_smul_89773 + p1_smul_89774;
  assign p2_add_92987_comb = p1_smul_90309 + p1_smul_90310;
  assign p2_add_92988_comb = p1_smul_90311 + p1_smul_90312;
  assign p2_add_92647_comb = p1_smul_89767 + p1_smul_89768;
  assign p2_add_92648_comb = p1_smul_89769 + p1_smul_89770;
  assign p2_add_92983_comb = p1_smul_90303 + p1_smul_90304;
  assign p2_add_92984_comb = p1_smul_90305 + p1_smul_90306;
  assign p2_add_92645_comb = p1_smul_89763 + p1_smul_89764;
  assign p2_add_92646_comb = p1_smul_89765 + p1_smul_89766;
  assign p2_add_92979_comb = p1_smul_90297 + p1_smul_90298;
  assign p2_add_92980_comb = p1_smul_90299 + p1_smul_90300;
  assign p2_add_92643_comb = p1_smul_89759 + p1_smul_89760;
  assign p2_add_92644_comb = p1_smul_89761 + p1_smul_89762;
  assign p2_add_92975_comb = p1_smul_90291 + p1_smul_90292;
  assign p2_add_92976_comb = p1_smul_90293 + p1_smul_90294;
  assign p2_add_92641_comb = p1_smul_89755 + p1_smul_89756;
  assign p2_add_92642_comb = p1_smul_89757 + p1_smul_89758;
  assign p2_add_92971_comb = p1_smul_90285 + p1_smul_90286;
  assign p2_add_92972_comb = p1_smul_90287 + p1_smul_90288;
  assign p2_add_92639_comb = p1_smul_89751 + p1_smul_89752;
  assign p2_add_92640_comb = p1_smul_89753 + p1_smul_89754;
  assign p2_add_92967_comb = p1_smul_90279 + p1_smul_90280;
  assign p2_add_92968_comb = p1_smul_90281 + p1_smul_90282;
  assign p2_add_92637_comb = p1_smul_89747 + p1_smul_89748;
  assign p2_add_92638_comb = p1_smul_89749 + p1_smul_89750;
  assign p2_add_92963_comb = p1_smul_90273 + p1_smul_90274;
  assign p2_add_92964_comb = p1_smul_90275 + p1_smul_90276;
  assign p2_add_92635_comb = p1_smul_89743 + p1_smul_89744;
  assign p2_add_92636_comb = p1_smul_89745 + p1_smul_89746;
  assign p2_add_92959_comb = p1_smul_90267 + p1_smul_90268;
  assign p2_add_92960_comb = p1_smul_90269 + p1_smul_90270;
  assign p2_add_92633_comb = p1_smul_89739 + p1_smul_89740;
  assign p2_add_92634_comb = p1_smul_89741 + p1_smul_89742;
  assign p2_add_92955_comb = p1_smul_90261 + p1_smul_90262;
  assign p2_add_92956_comb = p1_smul_90263 + p1_smul_90264;
  assign p2_add_92631_comb = p1_smul_89735 + p1_smul_89736;
  assign p2_add_92632_comb = p1_smul_89737 + p1_smul_89738;
  assign p2_add_92951_comb = p1_smul_90255 + p1_smul_90256;
  assign p2_add_92952_comb = p1_smul_90257 + p1_smul_90258;
  assign p2_add_92629_comb = p1_smul_89731 + p1_smul_89732;
  assign p2_add_92630_comb = p1_smul_89733 + p1_smul_89734;
  assign p2_add_92947_comb = p1_smul_90249 + p1_smul_90250;
  assign p2_add_92948_comb = p1_smul_90251 + p1_smul_90252;
  assign p2_add_92627_comb = p1_smul_89727 + p1_smul_89728;
  assign p2_add_92628_comb = p1_smul_89729 + p1_smul_89730;
  assign p2_add_92943_comb = p1_smul_90243 + p1_smul_90244;
  assign p2_add_92944_comb = p1_smul_90245 + p1_smul_90246;
  assign p2_add_92625_comb = p1_smul_89723 + p1_smul_89724;
  assign p2_add_92626_comb = p1_smul_89725 + p1_smul_89726;
  assign p2_add_92939_comb = p1_smul_90237 + p1_smul_90238;
  assign p2_add_92940_comb = p1_smul_90239 + p1_smul_90240;
  assign p2_add_92623_comb = p1_smul_89719 + p1_smul_89720;
  assign p2_add_92624_comb = p1_smul_89721 + p1_smul_89722;
  assign p2_add_92935_comb = p1_smul_90231 + p1_smul_90232;
  assign p2_add_92936_comb = p1_smul_90233 + p1_smul_90234;
  assign p2_add_92621_comb = p1_smul_89715 + p1_smul_89716;
  assign p2_add_92622_comb = p1_smul_89717 + p1_smul_89718;
  assign p2_add_92931_comb = p1_smul_90225 + p1_smul_90226;
  assign p2_add_92932_comb = p1_smul_90227 + p1_smul_90228;
  assign p2_add_92619_comb = p1_smul_89711 + p1_smul_89712;
  assign p2_add_92620_comb = p1_smul_89713 + p1_smul_89714;
  assign p2_add_92927_comb = p1_smul_90219 + p1_smul_90220;
  assign p2_add_92928_comb = p1_smul_90221 + p1_smul_90222;
  assign p2_add_92617_comb = p1_smul_89707 + p1_smul_89708;
  assign p2_add_92618_comb = p1_smul_89709 + p1_smul_89710;
  assign p2_add_92923_comb = p1_smul_90213 + p1_smul_90214;
  assign p2_add_92924_comb = p1_smul_90215 + p1_smul_90216;
  assign p2_add_92615_comb = p1_smul_89703 + p1_smul_89704;
  assign p2_add_92616_comb = p1_smul_89705 + p1_smul_89706;
  assign p2_add_92919_comb = p1_smul_90207 + p1_smul_90208;
  assign p2_add_92920_comb = p1_smul_90209 + p1_smul_90210;
  assign p2_add_92613_comb = p1_smul_89699 + p1_smul_89700;
  assign p2_add_92614_comb = p1_smul_89701 + p1_smul_89702;
  assign p2_add_92915_comb = p1_smul_90201 + p1_smul_90202;
  assign p2_add_92916_comb = p1_smul_90203 + p1_smul_90204;
  assign p2_add_92611_comb = p1_smul_89695 + p1_smul_89696;
  assign p2_add_92612_comb = p1_smul_89697 + p1_smul_89698;
  assign p2_add_92911_comb = p1_smul_90195 + p1_smul_90196;
  assign p2_add_92912_comb = p1_smul_90197 + p1_smul_90198;
  assign p2_add_92609_comb = p1_smul_89691 + p1_smul_89692;
  assign p2_add_92610_comb = p1_smul_89693 + p1_smul_89694;
  assign p2_add_92907_comb = p1_smul_90189 + p1_smul_90190;
  assign p2_add_92908_comb = p1_smul_90191 + p1_smul_90192;
  assign p2_add_92607_comb = p1_smul_89687 + p1_smul_89688;
  assign p2_add_92608_comb = p1_smul_89689 + p1_smul_89690;
  assign p2_add_92903_comb = p1_smul_90183 + p1_smul_90184;
  assign p2_add_92904_comb = p1_smul_90185 + p1_smul_90186;
  assign p2_add_92605_comb = p1_smul_89683 + p1_smul_89684;
  assign p2_add_92606_comb = p1_smul_89685 + p1_smul_89686;
  assign p2_add_92899_comb = p1_smul_90177 + p1_smul_90178;
  assign p2_add_92900_comb = p1_smul_90179 + p1_smul_90180;
  assign p2_add_92603_comb = p1_smul_89679 + p1_smul_89680;
  assign p2_add_92604_comb = p1_smul_89681 + p1_smul_89682;
  assign p2_add_92895_comb = p1_smul_90171 + p1_smul_90172;
  assign p2_add_92896_comb = p1_smul_90173 + p1_smul_90174;
  assign p2_add_92601_comb = p1_smul_89675 + p1_smul_89676;
  assign p2_add_92602_comb = p1_smul_89677 + p1_smul_89678;
  assign p2_add_92891_comb = p1_smul_90165 + p1_smul_90166;
  assign p2_add_92892_comb = p1_smul_90167 + p1_smul_90168;
  assign p2_add_92599_comb = p1_smul_89671 + p1_smul_89672;
  assign p2_add_92600_comb = p1_smul_89673 + p1_smul_89674;
  assign p2_add_92887_comb = p1_smul_90159 + p1_smul_90160;
  assign p2_add_92888_comb = p1_smul_90161 + p1_smul_90162;
  assign p2_add_92597_comb = p1_smul_89667 + p1_smul_89668;
  assign p2_add_92598_comb = p1_smul_89669 + p1_smul_89670;
  assign p2_add_92883_comb = p1_smul_90153 + p1_smul_90154;
  assign p2_add_92884_comb = p1_smul_90155 + p1_smul_90156;
  assign p2_add_92595_comb = p1_smul_89663 + p1_smul_89664;
  assign p2_add_92596_comb = p1_smul_89665 + p1_smul_89666;
  assign p2_add_92879_comb = p1_smul_90147 + p1_smul_90148;
  assign p2_add_92880_comb = p1_smul_90149 + p1_smul_90150;
  assign p2_add_92593_comb = p1_smul_89659 + p1_smul_89660;
  assign p2_add_92594_comb = p1_smul_89661 + p1_smul_89662;
  assign p2_add_92875_comb = p1_smul_90141 + p1_smul_90142;
  assign p2_add_92876_comb = p1_smul_90143 + p1_smul_90144;
  assign p2_add_92591_comb = p1_smul_89655 + p1_smul_89656;
  assign p2_add_92592_comb = p1_smul_89657 + p1_smul_89658;
  assign p2_add_92871_comb = p1_smul_90135 + p1_smul_90136;
  assign p2_add_92872_comb = p1_smul_90137 + p1_smul_90138;
  assign p2_add_92589_comb = p1_smul_89651 + p1_smul_89652;
  assign p2_add_92590_comb = p1_smul_89653 + p1_smul_89654;
  assign p2_add_92867_comb = p1_smul_90129 + p1_smul_90130;
  assign p2_add_92868_comb = p1_smul_90131 + p1_smul_90132;
  assign p2_add_92587_comb = p1_smul_89647 + p1_smul_89648;
  assign p2_add_92588_comb = p1_smul_89649 + p1_smul_89650;
  assign p2_add_92863_comb = p1_smul_90123 + p1_smul_90124;
  assign p2_add_92864_comb = p1_smul_90125 + p1_smul_90126;
  assign p2_add_92585_comb = p1_smul_89643 + p1_smul_89644;
  assign p2_add_92586_comb = p1_smul_89645 + p1_smul_89646;
  assign p2_add_92859_comb = p1_smul_90117 + p1_smul_90118;
  assign p2_add_92860_comb = p1_smul_90119 + p1_smul_90120;
  assign p2_add_92583_comb = p1_smul_89639 + p1_smul_89640;
  assign p2_add_92584_comb = p1_smul_89641 + p1_smul_89642;
  assign p2_add_92855_comb = p1_smul_90111 + p1_smul_90112;
  assign p2_add_92856_comb = p1_smul_90113 + p1_smul_90114;
  assign p2_add_92581_comb = p1_smul_89635 + p1_smul_89636;
  assign p2_add_92582_comb = p1_smul_89637 + p1_smul_89638;
  assign p2_add_92851_comb = p1_smul_90105 + p1_smul_90106;
  assign p2_add_92852_comb = p1_smul_90107 + p1_smul_90108;
  assign p2_add_92579_comb = p1_smul_89631 + p1_smul_89632;
  assign p2_add_92580_comb = p1_smul_89633 + p1_smul_89634;
  assign p2_add_92847_comb = p1_smul_90099 + p1_smul_90100;
  assign p2_add_92848_comb = p1_smul_90101 + p1_smul_90102;
  assign p2_add_92577_comb = p1_smul_89627 + p1_smul_89628;
  assign p2_add_92578_comb = p1_smul_89629 + p1_smul_89630;
  assign p2_add_92843_comb = p1_smul_90093 + p1_smul_90094;
  assign p2_add_92844_comb = p1_smul_90095 + p1_smul_90096;
  assign p2_add_92575_comb = p1_smul_89623 + p1_smul_89624;
  assign p2_add_92576_comb = p1_smul_89625 + p1_smul_89626;
  assign p2_add_92839_comb = p1_smul_90087 + p1_smul_90088;
  assign p2_add_92840_comb = p1_smul_90089 + p1_smul_90090;
  assign p2_add_92573_comb = p1_smul_89619 + p1_smul_89620;
  assign p2_add_92574_comb = p1_smul_89621 + p1_smul_89622;
  assign p2_add_92835_comb = p1_smul_90081 + p1_smul_90082;
  assign p2_add_92836_comb = p1_smul_90083 + p1_smul_90084;
  assign p2_add_92571_comb = p1_smul_89615 + p1_smul_89616;
  assign p2_add_92572_comb = p1_smul_89617 + p1_smul_89618;
  assign p2_add_92831_comb = p1_smul_90075 + p1_smul_90076;
  assign p2_add_92832_comb = p1_smul_90077 + p1_smul_90078;
  assign p2_add_92569_comb = p1_smul_89611 + p1_smul_89612;
  assign p2_add_92570_comb = p1_smul_89613 + p1_smul_89614;
  assign p2_add_92827_comb = p1_smul_90069 + p1_smul_90070;
  assign p2_add_92828_comb = p1_smul_90071 + p1_smul_90072;
  assign p2_add_92567_comb = p1_smul_89607 + p1_smul_89608;
  assign p2_add_92568_comb = p1_smul_89609 + p1_smul_89610;
  assign p2_add_92823_comb = p1_smul_90063 + p1_smul_90064;
  assign p2_add_92824_comb = p1_smul_90065 + p1_smul_90066;
  assign p2_add_92565_comb = p1_smul_89603 + p1_smul_89604;
  assign p2_add_92566_comb = p1_smul_89605 + p1_smul_89606;
  assign p2_add_92819_comb = p1_smul_90057 + p1_smul_90058;
  assign p2_add_92820_comb = p1_smul_90059 + p1_smul_90060;
  assign p2_add_92563_comb = p1_smul_89599 + p1_smul_89600;
  assign p2_add_92564_comb = p1_smul_89601 + p1_smul_89602;
  assign p2_add_92815_comb = p1_smul_90051 + p1_smul_90052;
  assign p2_add_92816_comb = p1_smul_90053 + p1_smul_90054;
  assign p2_add_92561_comb = p1_smul_89595 + p1_smul_89596;
  assign p2_add_92562_comb = p1_smul_89597 + p1_smul_89598;
  assign p2_add_92811_comb = p1_smul_90045 + p1_smul_90046;
  assign p2_add_92812_comb = p1_smul_90047 + p1_smul_90048;
  assign p2_add_92559_comb = p1_smul_89591 + p1_smul_89592;
  assign p2_add_92560_comb = p1_smul_89593 + p1_smul_89594;
  assign p2_add_92807_comb = p1_smul_90039 + p1_smul_90040;
  assign p2_add_92808_comb = p1_smul_90041 + p1_smul_90042;
  assign p2_add_92557_comb = p1_smul_89587 + p1_smul_89588;
  assign p2_add_92558_comb = p1_smul_89589 + p1_smul_89590;
  assign p2_add_92803_comb = p1_smul_90033 + p1_smul_90034;
  assign p2_add_92804_comb = p1_smul_90035 + p1_smul_90036;
  assign p2_add_92555_comb = p1_smul_89583 + p1_smul_89584;
  assign p2_add_92556_comb = p1_smul_89585 + p1_smul_89586;
  assign p2_add_92799_comb = p1_smul_90027 + p1_smul_90028;
  assign p2_add_92800_comb = p1_smul_90029 + p1_smul_90030;
  assign p2_add_92553_comb = p1_smul_89579 + p1_smul_89580;
  assign p2_add_92554_comb = p1_smul_89581 + p1_smul_89582;
  assign p2_add_92795_comb = p1_smul_90021 + p1_smul_90022;
  assign p2_add_92796_comb = p1_smul_90023 + p1_smul_90024;
  assign p2_add_92551_comb = p1_smul_89575 + p1_smul_89576;
  assign p2_add_92552_comb = p1_smul_89577 + p1_smul_89578;
  assign p2_add_92791_comb = p1_smul_90015 + p1_smul_90016;
  assign p2_add_92792_comb = p1_smul_90017 + p1_smul_90018;
  assign p2_add_92549_comb = p1_smul_89571 + p1_smul_89572;
  assign p2_add_92550_comb = p1_smul_89573 + p1_smul_89574;
  assign p2_add_92787_comb = p1_smul_90009 + p1_smul_90010;
  assign p2_add_92788_comb = p1_smul_90011 + p1_smul_90012;
  assign p2_add_92547_comb = p1_smul_89567 + p1_smul_89568;
  assign p2_add_92548_comb = p1_smul_89569 + p1_smul_89570;
  assign p2_add_92783_comb = p1_smul_90003 + p1_smul_90004;
  assign p2_add_92784_comb = p1_smul_90005 + p1_smul_90006;
  assign p2_add_92545_comb = p1_smul_89563 + p1_smul_89564;
  assign p2_add_92546_comb = p1_smul_89565 + p1_smul_89566;
  assign p2_add_92779_comb = p1_smul_89997 + p1_smul_89998;
  assign p2_add_92780_comb = p1_smul_89999 + p1_smul_90000;
  assign p2_add_92543_comb = p1_smul_89559 + p1_smul_89560;
  assign p2_add_92544_comb = p1_smul_89561 + p1_smul_89562;
  assign p2_add_92775_comb = p1_smul_89991 + p1_smul_89992;
  assign p2_add_92776_comb = p1_smul_89993 + p1_smul_89994;
  assign p2_add_92541_comb = p1_smul_89555 + p1_smul_89556;
  assign p2_add_92542_comb = p1_smul_89557 + p1_smul_89558;
  assign p2_add_92771_comb = p1_smul_89985 + p1_smul_89986;
  assign p2_add_92772_comb = p1_smul_89987 + p1_smul_89988;
  assign p2_add_92539_comb = p1_smul_89551 + p1_smul_89552;
  assign p2_add_92540_comb = p1_smul_89553 + p1_smul_89554;
  assign p2_add_92767_comb = p1_smul_89979 + p1_smul_89980;
  assign p2_add_92768_comb = p1_smul_89981 + p1_smul_89982;
  assign p2_add_92537_comb = p1_smul_89547 + p1_smul_89548;
  assign p2_add_92538_comb = p1_smul_89549 + p1_smul_89550;
  assign p2_add_92763_comb = p1_smul_89973 + p1_smul_89974;
  assign p2_add_92764_comb = p1_smul_89975 + p1_smul_89976;
  assign p2_add_92535_comb = p1_smul_89543 + p1_smul_89544;
  assign p2_add_92536_comb = p1_smul_89545 + p1_smul_89546;
  assign p2_add_92759_comb = p1_smul_89967 + p1_smul_89968;
  assign p2_add_92760_comb = p1_smul_89969 + p1_smul_89970;
  assign p2_add_92533_comb = p1_smul_89539 + p1_smul_89540;
  assign p2_add_92534_comb = p1_smul_89541 + p1_smul_89542;
  assign p2_add_92755_comb = p1_smul_89961 + p1_smul_89962;
  assign p2_add_92756_comb = p1_smul_89963 + p1_smul_89964;
  assign p2_add_92531_comb = p1_smul_89535 + p1_smul_89536;
  assign p2_add_92532_comb = p1_smul_89537 + p1_smul_89538;
  assign p2_add_92751_comb = p1_smul_89955 + p1_smul_89956;
  assign p2_add_92752_comb = p1_smul_89957 + p1_smul_89958;
  assign p2_add_92529_comb = p1_smul_89531 + p1_smul_89532;
  assign p2_add_92530_comb = p1_smul_89533 + p1_smul_89534;
  assign p2_add_92747_comb = p1_smul_89949 + p1_smul_89950;
  assign p2_add_92748_comb = p1_smul_89951 + p1_smul_89952;
  assign p2_add_92527_comb = p1_smul_89527 + p1_smul_89528;
  assign p2_add_92528_comb = p1_smul_89529 + p1_smul_89530;
  assign p2_add_92743_comb = p1_smul_89943 + p1_smul_89944;
  assign p2_add_92744_comb = p1_smul_89945 + p1_smul_89946;
  assign p2_add_92525_comb = p1_smul_89523 + p1_smul_89524;
  assign p2_add_92526_comb = p1_smul_89525 + p1_smul_89526;
  assign p2_add_92739_comb = p1_smul_89937 + p1_smul_89938;
  assign p2_add_92740_comb = p1_smul_89939 + p1_smul_89940;
  assign p2_add_92523_comb = p1_smul_89519 + p1_smul_89520;
  assign p2_add_92524_comb = p1_smul_89521 + p1_smul_89522;
  assign p2_add_92735_comb = p1_smul_89931 + p1_smul_89932;
  assign p2_add_92736_comb = p1_smul_89933 + p1_smul_89934;
  assign p2_add_92521_comb = p1_smul_89515 + p1_smul_89516;
  assign p2_add_92522_comb = p1_smul_89517 + p1_smul_89518;
  assign p2_add_92731_comb = p1_smul_89925 + p1_smul_89926;
  assign p2_add_92732_comb = p1_smul_89927 + p1_smul_89928;
  assign p2_add_92519_comb = p1_smul_89511 + p1_smul_89512;
  assign p2_add_92520_comb = p1_smul_89513 + p1_smul_89514;
  assign p2_add_92727_comb = p1_smul_89919 + p1_smul_89920;
  assign p2_add_92728_comb = p1_smul_89921 + p1_smul_89922;
  assign p2_add_92517_comb = p1_smul_89507 + p1_smul_89508;
  assign p2_add_92518_comb = p1_smul_89509 + p1_smul_89510;
  assign p2_add_92723_comb = p1_smul_89913 + p1_smul_89914;
  assign p2_add_92724_comb = p1_smul_89915 + p1_smul_89916;
  assign p2_add_92515_comb = p1_smul_89503 + p1_smul_89504;
  assign p2_add_92516_comb = p1_smul_89505 + p1_smul_89506;
  assign p2_add_92719_comb = p1_smul_89907 + p1_smul_89908;
  assign p2_add_92720_comb = p1_smul_89909 + p1_smul_89910;
  assign p2_add_92513_comb = p1_smul_89499 + p1_smul_89500;
  assign p2_add_92514_comb = p1_smul_89501 + p1_smul_89502;
  assign p2_add_92715_comb = p1_smul_89901 + p1_smul_89902;
  assign p2_add_92716_comb = p1_smul_89903 + p1_smul_89904;
  assign p2_add_93109_comb = p2_add_92711_comb + p2_add_92712_comb;
  assign p2_add_93110_comb = p1_smul_90493 + p1_smul_90494;
  assign p2_add_93212_comb = p2_add_93111_comb + p2_add_93112_comb;
  assign p2_add_93105_comb = p2_add_92709_comb + p2_add_92710_comb;
  assign p2_add_93106_comb = p1_smul_90487 + p1_smul_90488;
  assign p2_add_93211_comb = p2_add_93107_comb + p2_add_93108_comb;
  assign p2_add_93101_comb = p2_add_92707_comb + p2_add_92708_comb;
  assign p2_add_93102_comb = p1_smul_90481 + p1_smul_90482;
  assign p2_add_93210_comb = p2_add_93103_comb + p2_add_93104_comb;
  assign p2_add_93097_comb = p2_add_92705_comb + p2_add_92706_comb;
  assign p2_add_93098_comb = p1_smul_90475 + p1_smul_90476;
  assign p2_add_93209_comb = p2_add_93099_comb + p2_add_93100_comb;
  assign p2_add_93093_comb = p2_add_92703_comb + p2_add_92704_comb;
  assign p2_add_93094_comb = p1_smul_90469 + p1_smul_90470;
  assign p2_add_93208_comb = p2_add_93095_comb + p2_add_93096_comb;
  assign p2_add_93089_comb = p2_add_92701_comb + p2_add_92702_comb;
  assign p2_add_93090_comb = p1_smul_90463 + p1_smul_90464;
  assign p2_add_93207_comb = p2_add_93091_comb + p2_add_93092_comb;
  assign p2_add_93085_comb = p2_add_92699_comb + p2_add_92700_comb;
  assign p2_add_93086_comb = p1_smul_90457 + p1_smul_90458;
  assign p2_add_93206_comb = p2_add_93087_comb + p2_add_93088_comb;
  assign p2_add_93081_comb = p2_add_92697_comb + p2_add_92698_comb;
  assign p2_add_93082_comb = p1_smul_90451 + p1_smul_90452;
  assign p2_add_93205_comb = p2_add_93083_comb + p2_add_93084_comb;
  assign p2_add_93077_comb = p2_add_92695_comb + p2_add_92696_comb;
  assign p2_add_93078_comb = p1_smul_90445 + p1_smul_90446;
  assign p2_add_93204_comb = p2_add_93079_comb + p2_add_93080_comb;
  assign p2_add_93073_comb = p2_add_92693_comb + p2_add_92694_comb;
  assign p2_add_93074_comb = p1_smul_90439 + p1_smul_90440;
  assign p2_add_93203_comb = p2_add_93075_comb + p2_add_93076_comb;
  assign p2_add_93069_comb = p2_add_92691_comb + p2_add_92692_comb;
  assign p2_add_93070_comb = p1_smul_90433 + p1_smul_90434;
  assign p2_add_93202_comb = p2_add_93071_comb + p2_add_93072_comb;
  assign p2_add_93065_comb = p2_add_92689_comb + p2_add_92690_comb;
  assign p2_add_93066_comb = p1_smul_90427 + p1_smul_90428;
  assign p2_add_93201_comb = p2_add_93067_comb + p2_add_93068_comb;
  assign p2_add_93061_comb = p2_add_92687_comb + p2_add_92688_comb;
  assign p2_add_93062_comb = p1_smul_90421 + p1_smul_90422;
  assign p2_add_93200_comb = p2_add_93063_comb + p2_add_93064_comb;
  assign p2_add_93057_comb = p2_add_92685_comb + p2_add_92686_comb;
  assign p2_add_93058_comb = p1_smul_90415 + p1_smul_90416;
  assign p2_add_93199_comb = p2_add_93059_comb + p2_add_93060_comb;
  assign p2_add_93053_comb = p2_add_92683_comb + p2_add_92684_comb;
  assign p2_add_93054_comb = p1_smul_90409 + p1_smul_90410;
  assign p2_add_93198_comb = p2_add_93055_comb + p2_add_93056_comb;
  assign p2_add_93049_comb = p2_add_92681_comb + p2_add_92682_comb;
  assign p2_add_93050_comb = p1_smul_90403 + p1_smul_90404;
  assign p2_add_93197_comb = p2_add_93051_comb + p2_add_93052_comb;
  assign p2_add_93045_comb = p2_add_92679_comb + p2_add_92680_comb;
  assign p2_add_93046_comb = p1_smul_90397 + p1_smul_90398;
  assign p2_add_93196_comb = p2_add_93047_comb + p2_add_93048_comb;
  assign p2_add_93041_comb = p2_add_92677_comb + p2_add_92678_comb;
  assign p2_add_93042_comb = p1_smul_90391 + p1_smul_90392;
  assign p2_add_93195_comb = p2_add_93043_comb + p2_add_93044_comb;
  assign p2_add_93037_comb = p2_add_92675_comb + p2_add_92676_comb;
  assign p2_add_93038_comb = p1_smul_90385 + p1_smul_90386;
  assign p2_add_93194_comb = p2_add_93039_comb + p2_add_93040_comb;
  assign p2_add_93033_comb = p2_add_92673_comb + p2_add_92674_comb;
  assign p2_add_93034_comb = p1_smul_90379 + p1_smul_90380;
  assign p2_add_93193_comb = p2_add_93035_comb + p2_add_93036_comb;
  assign p2_add_93029_comb = p2_add_92671_comb + p2_add_92672_comb;
  assign p2_add_93030_comb = p1_smul_90373 + p1_smul_90374;
  assign p2_add_93192_comb = p2_add_93031_comb + p2_add_93032_comb;
  assign p2_add_93025_comb = p2_add_92669_comb + p2_add_92670_comb;
  assign p2_add_93026_comb = p1_smul_90367 + p1_smul_90368;
  assign p2_add_93191_comb = p2_add_93027_comb + p2_add_93028_comb;
  assign p2_add_93021_comb = p2_add_92667_comb + p2_add_92668_comb;
  assign p2_add_93022_comb = p1_smul_90361 + p1_smul_90362;
  assign p2_add_93190_comb = p2_add_93023_comb + p2_add_93024_comb;
  assign p2_add_93017_comb = p2_add_92665_comb + p2_add_92666_comb;
  assign p2_add_93018_comb = p1_smul_90355 + p1_smul_90356;
  assign p2_add_93189_comb = p2_add_93019_comb + p2_add_93020_comb;
  assign p2_add_93013_comb = p2_add_92663_comb + p2_add_92664_comb;
  assign p2_add_93014_comb = p1_smul_90349 + p1_smul_90350;
  assign p2_add_93188_comb = p2_add_93015_comb + p2_add_93016_comb;
  assign p2_add_93009_comb = p2_add_92661_comb + p2_add_92662_comb;
  assign p2_add_93010_comb = p1_smul_90343 + p1_smul_90344;
  assign p2_add_93187_comb = p2_add_93011_comb + p2_add_93012_comb;
  assign p2_add_93005_comb = p2_add_92659_comb + p2_add_92660_comb;
  assign p2_add_93006_comb = p1_smul_90337 + p1_smul_90338;
  assign p2_add_93186_comb = p2_add_93007_comb + p2_add_93008_comb;
  assign p2_add_93001_comb = p2_add_92657_comb + p2_add_92658_comb;
  assign p2_add_93002_comb = p1_smul_90331 + p1_smul_90332;
  assign p2_add_93185_comb = p2_add_93003_comb + p2_add_93004_comb;
  assign p2_add_92997_comb = p2_add_92655_comb + p2_add_92656_comb;
  assign p2_add_92998_comb = p1_smul_90325 + p1_smul_90326;
  assign p2_add_93184_comb = p2_add_92999_comb + p2_add_93000_comb;
  assign p2_add_92993_comb = p2_add_92653_comb + p2_add_92654_comb;
  assign p2_add_92994_comb = p1_smul_90319 + p1_smul_90320;
  assign p2_add_93183_comb = p2_add_92995_comb + p2_add_92996_comb;
  assign p2_add_92989_comb = p2_add_92651_comb + p2_add_92652_comb;
  assign p2_add_92990_comb = p1_smul_90313 + p1_smul_90314;
  assign p2_add_93182_comb = p2_add_92991_comb + p2_add_92992_comb;
  assign p2_add_92985_comb = p2_add_92649_comb + p2_add_92650_comb;
  assign p2_add_92986_comb = p1_smul_90307 + p1_smul_90308;
  assign p2_add_93181_comb = p2_add_92987_comb + p2_add_92988_comb;
  assign p2_add_92981_comb = p2_add_92647_comb + p2_add_92648_comb;
  assign p2_add_92982_comb = p1_smul_90301 + p1_smul_90302;
  assign p2_add_93180_comb = p2_add_92983_comb + p2_add_92984_comb;
  assign p2_add_92977_comb = p2_add_92645_comb + p2_add_92646_comb;
  assign p2_add_92978_comb = p1_smul_90295 + p1_smul_90296;
  assign p2_add_93179_comb = p2_add_92979_comb + p2_add_92980_comb;
  assign p2_add_92973_comb = p2_add_92643_comb + p2_add_92644_comb;
  assign p2_add_92974_comb = p1_smul_90289 + p1_smul_90290;
  assign p2_add_93178_comb = p2_add_92975_comb + p2_add_92976_comb;
  assign p2_add_92969_comb = p2_add_92641_comb + p2_add_92642_comb;
  assign p2_add_92970_comb = p1_smul_90283 + p1_smul_90284;
  assign p2_add_93177_comb = p2_add_92971_comb + p2_add_92972_comb;
  assign p2_add_92965_comb = p2_add_92639_comb + p2_add_92640_comb;
  assign p2_add_92966_comb = p1_smul_90277 + p1_smul_90278;
  assign p2_add_93176_comb = p2_add_92967_comb + p2_add_92968_comb;
  assign p2_add_92961_comb = p2_add_92637_comb + p2_add_92638_comb;
  assign p2_add_92962_comb = p1_smul_90271 + p1_smul_90272;
  assign p2_add_93175_comb = p2_add_92963_comb + p2_add_92964_comb;
  assign p2_add_92957_comb = p2_add_92635_comb + p2_add_92636_comb;
  assign p2_add_92958_comb = p1_smul_90265 + p1_smul_90266;
  assign p2_add_93174_comb = p2_add_92959_comb + p2_add_92960_comb;
  assign p2_add_92953_comb = p2_add_92633_comb + p2_add_92634_comb;
  assign p2_add_92954_comb = p1_smul_90259 + p1_smul_90260;
  assign p2_add_93173_comb = p2_add_92955_comb + p2_add_92956_comb;
  assign p2_add_92949_comb = p2_add_92631_comb + p2_add_92632_comb;
  assign p2_add_92950_comb = p1_smul_90253 + p1_smul_90254;
  assign p2_add_93172_comb = p2_add_92951_comb + p2_add_92952_comb;
  assign p2_add_92945_comb = p2_add_92629_comb + p2_add_92630_comb;
  assign p2_add_92946_comb = p1_smul_90247 + p1_smul_90248;
  assign p2_add_93171_comb = p2_add_92947_comb + p2_add_92948_comb;
  assign p2_add_92941_comb = p2_add_92627_comb + p2_add_92628_comb;
  assign p2_add_92942_comb = p1_smul_90241 + p1_smul_90242;
  assign p2_add_93170_comb = p2_add_92943_comb + p2_add_92944_comb;
  assign p2_add_92937_comb = p2_add_92625_comb + p2_add_92626_comb;
  assign p2_add_92938_comb = p1_smul_90235 + p1_smul_90236;
  assign p2_add_93169_comb = p2_add_92939_comb + p2_add_92940_comb;
  assign p2_add_92933_comb = p2_add_92623_comb + p2_add_92624_comb;
  assign p2_add_92934_comb = p1_smul_90229 + p1_smul_90230;
  assign p2_add_93168_comb = p2_add_92935_comb + p2_add_92936_comb;
  assign p2_add_92929_comb = p2_add_92621_comb + p2_add_92622_comb;
  assign p2_add_92930_comb = p1_smul_90223 + p1_smul_90224;
  assign p2_add_93167_comb = p2_add_92931_comb + p2_add_92932_comb;
  assign p2_add_92925_comb = p2_add_92619_comb + p2_add_92620_comb;
  assign p2_add_92926_comb = p1_smul_90217 + p1_smul_90218;
  assign p2_add_93166_comb = p2_add_92927_comb + p2_add_92928_comb;
  assign p2_add_92921_comb = p2_add_92617_comb + p2_add_92618_comb;
  assign p2_add_92922_comb = p1_smul_90211 + p1_smul_90212;
  assign p2_add_93165_comb = p2_add_92923_comb + p2_add_92924_comb;
  assign p2_add_92917_comb = p2_add_92615_comb + p2_add_92616_comb;
  assign p2_add_92918_comb = p1_smul_90205 + p1_smul_90206;
  assign p2_add_93164_comb = p2_add_92919_comb + p2_add_92920_comb;
  assign p2_add_92913_comb = p2_add_92613_comb + p2_add_92614_comb;
  assign p2_add_92914_comb = p1_smul_90199 + p1_smul_90200;
  assign p2_add_93163_comb = p2_add_92915_comb + p2_add_92916_comb;
  assign p2_add_92909_comb = p2_add_92611_comb + p2_add_92612_comb;
  assign p2_add_92910_comb = p1_smul_90193 + p1_smul_90194;
  assign p2_add_93162_comb = p2_add_92911_comb + p2_add_92912_comb;
  assign p2_add_92905_comb = p2_add_92609_comb + p2_add_92610_comb;
  assign p2_add_92906_comb = p1_smul_90187 + p1_smul_90188;
  assign p2_add_93161_comb = p2_add_92907_comb + p2_add_92908_comb;
  assign p2_add_92901_comb = p2_add_92607_comb + p2_add_92608_comb;
  assign p2_add_92902_comb = p1_smul_90181 + p1_smul_90182;
  assign p2_add_93160_comb = p2_add_92903_comb + p2_add_92904_comb;
  assign p2_add_92897_comb = p2_add_92605_comb + p2_add_92606_comb;
  assign p2_add_92898_comb = p1_smul_90175 + p1_smul_90176;
  assign p2_add_93159_comb = p2_add_92899_comb + p2_add_92900_comb;
  assign p2_add_92893_comb = p2_add_92603_comb + p2_add_92604_comb;
  assign p2_add_92894_comb = p1_smul_90169 + p1_smul_90170;
  assign p2_add_93158_comb = p2_add_92895_comb + p2_add_92896_comb;
  assign p2_add_92889_comb = p2_add_92601_comb + p2_add_92602_comb;
  assign p2_add_92890_comb = p1_smul_90163 + p1_smul_90164;
  assign p2_add_93157_comb = p2_add_92891_comb + p2_add_92892_comb;
  assign p2_add_92885_comb = p2_add_92599_comb + p2_add_92600_comb;
  assign p2_add_92886_comb = p1_smul_90157 + p1_smul_90158;
  assign p2_add_93156_comb = p2_add_92887_comb + p2_add_92888_comb;
  assign p2_add_92881_comb = p2_add_92597_comb + p2_add_92598_comb;
  assign p2_add_92882_comb = p1_smul_90151 + p1_smul_90152;
  assign p2_add_93155_comb = p2_add_92883_comb + p2_add_92884_comb;
  assign p2_add_92877_comb = p2_add_92595_comb + p2_add_92596_comb;
  assign p2_add_92878_comb = p1_smul_90145 + p1_smul_90146;
  assign p2_add_93154_comb = p2_add_92879_comb + p2_add_92880_comb;
  assign p2_add_92873_comb = p2_add_92593_comb + p2_add_92594_comb;
  assign p2_add_92874_comb = p1_smul_90139 + p1_smul_90140;
  assign p2_add_93153_comb = p2_add_92875_comb + p2_add_92876_comb;
  assign p2_add_92869_comb = p2_add_92591_comb + p2_add_92592_comb;
  assign p2_add_92870_comb = p1_smul_90133 + p1_smul_90134;
  assign p2_add_93152_comb = p2_add_92871_comb + p2_add_92872_comb;
  assign p2_add_92865_comb = p2_add_92589_comb + p2_add_92590_comb;
  assign p2_add_92866_comb = p1_smul_90127 + p1_smul_90128;
  assign p2_add_93151_comb = p2_add_92867_comb + p2_add_92868_comb;
  assign p2_add_92861_comb = p2_add_92587_comb + p2_add_92588_comb;
  assign p2_add_92862_comb = p1_smul_90121 + p1_smul_90122;
  assign p2_add_93150_comb = p2_add_92863_comb + p2_add_92864_comb;
  assign p2_add_92857_comb = p2_add_92585_comb + p2_add_92586_comb;
  assign p2_add_92858_comb = p1_smul_90115 + p1_smul_90116;
  assign p2_add_93149_comb = p2_add_92859_comb + p2_add_92860_comb;
  assign p2_add_92853_comb = p2_add_92583_comb + p2_add_92584_comb;
  assign p2_add_92854_comb = p1_smul_90109 + p1_smul_90110;
  assign p2_add_93148_comb = p2_add_92855_comb + p2_add_92856_comb;
  assign p2_add_92849_comb = p2_add_92581_comb + p2_add_92582_comb;
  assign p2_add_92850_comb = p1_smul_90103 + p1_smul_90104;
  assign p2_add_93147_comb = p2_add_92851_comb + p2_add_92852_comb;
  assign p2_add_92845_comb = p2_add_92579_comb + p2_add_92580_comb;
  assign p2_add_92846_comb = p1_smul_90097 + p1_smul_90098;
  assign p2_add_93146_comb = p2_add_92847_comb + p2_add_92848_comb;
  assign p2_add_92841_comb = p2_add_92577_comb + p2_add_92578_comb;
  assign p2_add_92842_comb = p1_smul_90091 + p1_smul_90092;
  assign p2_add_93145_comb = p2_add_92843_comb + p2_add_92844_comb;
  assign p2_add_92837_comb = p2_add_92575_comb + p2_add_92576_comb;
  assign p2_add_92838_comb = p1_smul_90085 + p1_smul_90086;
  assign p2_add_93144_comb = p2_add_92839_comb + p2_add_92840_comb;
  assign p2_add_92833_comb = p2_add_92573_comb + p2_add_92574_comb;
  assign p2_add_92834_comb = p1_smul_90079 + p1_smul_90080;
  assign p2_add_93143_comb = p2_add_92835_comb + p2_add_92836_comb;
  assign p2_add_92829_comb = p2_add_92571_comb + p2_add_92572_comb;
  assign p2_add_92830_comb = p1_smul_90073 + p1_smul_90074;
  assign p2_add_93142_comb = p2_add_92831_comb + p2_add_92832_comb;
  assign p2_add_92825_comb = p2_add_92569_comb + p2_add_92570_comb;
  assign p2_add_92826_comb = p1_smul_90067 + p1_smul_90068;
  assign p2_add_93141_comb = p2_add_92827_comb + p2_add_92828_comb;
  assign p2_add_92821_comb = p2_add_92567_comb + p2_add_92568_comb;
  assign p2_add_92822_comb = p1_smul_90061 + p1_smul_90062;
  assign p2_add_93140_comb = p2_add_92823_comb + p2_add_92824_comb;
  assign p2_add_92817_comb = p2_add_92565_comb + p2_add_92566_comb;
  assign p2_add_92818_comb = p1_smul_90055 + p1_smul_90056;
  assign p2_add_93139_comb = p2_add_92819_comb + p2_add_92820_comb;
  assign p2_add_92813_comb = p2_add_92563_comb + p2_add_92564_comb;
  assign p2_add_92814_comb = p1_smul_90049 + p1_smul_90050;
  assign p2_add_93138_comb = p2_add_92815_comb + p2_add_92816_comb;
  assign p2_add_92809_comb = p2_add_92561_comb + p2_add_92562_comb;
  assign p2_add_92810_comb = p1_smul_90043 + p1_smul_90044;
  assign p2_add_93137_comb = p2_add_92811_comb + p2_add_92812_comb;
  assign p2_add_92805_comb = p2_add_92559_comb + p2_add_92560_comb;
  assign p2_add_92806_comb = p1_smul_90037 + p1_smul_90038;
  assign p2_add_93136_comb = p2_add_92807_comb + p2_add_92808_comb;
  assign p2_add_92801_comb = p2_add_92557_comb + p2_add_92558_comb;
  assign p2_add_92802_comb = p1_smul_90031 + p1_smul_90032;
  assign p2_add_93135_comb = p2_add_92803_comb + p2_add_92804_comb;
  assign p2_add_92797_comb = p2_add_92555_comb + p2_add_92556_comb;
  assign p2_add_92798_comb = p1_smul_90025 + p1_smul_90026;
  assign p2_add_93134_comb = p2_add_92799_comb + p2_add_92800_comb;
  assign p2_add_92793_comb = p2_add_92553_comb + p2_add_92554_comb;
  assign p2_add_92794_comb = p1_smul_90019 + p1_smul_90020;
  assign p2_add_93133_comb = p2_add_92795_comb + p2_add_92796_comb;
  assign p2_add_92789_comb = p2_add_92551_comb + p2_add_92552_comb;
  assign p2_add_92790_comb = p1_smul_90013 + p1_smul_90014;
  assign p2_add_93132_comb = p2_add_92791_comb + p2_add_92792_comb;
  assign p2_add_92785_comb = p2_add_92549_comb + p2_add_92550_comb;
  assign p2_add_92786_comb = p1_smul_90007 + p1_smul_90008;
  assign p2_add_93131_comb = p2_add_92787_comb + p2_add_92788_comb;
  assign p2_add_92781_comb = p2_add_92547_comb + p2_add_92548_comb;
  assign p2_add_92782_comb = p1_smul_90001 + p1_smul_90002;
  assign p2_add_93130_comb = p2_add_92783_comb + p2_add_92784_comb;
  assign p2_add_92777_comb = p2_add_92545_comb + p2_add_92546_comb;
  assign p2_add_92778_comb = p1_smul_89995 + p1_smul_89996;
  assign p2_add_93129_comb = p2_add_92779_comb + p2_add_92780_comb;
  assign p2_add_92773_comb = p2_add_92543_comb + p2_add_92544_comb;
  assign p2_add_92774_comb = p1_smul_89989 + p1_smul_89990;
  assign p2_add_93128_comb = p2_add_92775_comb + p2_add_92776_comb;
  assign p2_add_92769_comb = p2_add_92541_comb + p2_add_92542_comb;
  assign p2_add_92770_comb = p1_smul_89983 + p1_smul_89984;
  assign p2_add_93127_comb = p2_add_92771_comb + p2_add_92772_comb;
  assign p2_add_92765_comb = p2_add_92539_comb + p2_add_92540_comb;
  assign p2_add_92766_comb = p1_smul_89977 + p1_smul_89978;
  assign p2_add_93126_comb = p2_add_92767_comb + p2_add_92768_comb;
  assign p2_add_92761_comb = p2_add_92537_comb + p2_add_92538_comb;
  assign p2_add_92762_comb = p1_smul_89971 + p1_smul_89972;
  assign p2_add_93125_comb = p2_add_92763_comb + p2_add_92764_comb;
  assign p2_add_92757_comb = p2_add_92535_comb + p2_add_92536_comb;
  assign p2_add_92758_comb = p1_smul_89965 + p1_smul_89966;
  assign p2_add_93124_comb = p2_add_92759_comb + p2_add_92760_comb;
  assign p2_add_92753_comb = p2_add_92533_comb + p2_add_92534_comb;
  assign p2_add_92754_comb = p1_smul_89959 + p1_smul_89960;
  assign p2_add_93123_comb = p2_add_92755_comb + p2_add_92756_comb;
  assign p2_add_92749_comb = p2_add_92531_comb + p2_add_92532_comb;
  assign p2_add_92750_comb = p1_smul_89953 + p1_smul_89954;
  assign p2_add_93122_comb = p2_add_92751_comb + p2_add_92752_comb;
  assign p2_add_92745_comb = p2_add_92529_comb + p2_add_92530_comb;
  assign p2_add_92746_comb = p1_smul_89947 + p1_smul_89948;
  assign p2_add_93121_comb = p2_add_92747_comb + p2_add_92748_comb;
  assign p2_add_92741_comb = p2_add_92527_comb + p2_add_92528_comb;
  assign p2_add_92742_comb = p1_smul_89941 + p1_smul_89942;
  assign p2_add_93120_comb = p2_add_92743_comb + p2_add_92744_comb;
  assign p2_add_92737_comb = p2_add_92525_comb + p2_add_92526_comb;
  assign p2_add_92738_comb = p1_smul_89935 + p1_smul_89936;
  assign p2_add_93119_comb = p2_add_92739_comb + p2_add_92740_comb;
  assign p2_add_92733_comb = p2_add_92523_comb + p2_add_92524_comb;
  assign p2_add_92734_comb = p1_smul_89929 + p1_smul_89930;
  assign p2_add_93118_comb = p2_add_92735_comb + p2_add_92736_comb;
  assign p2_add_92729_comb = p2_add_92521_comb + p2_add_92522_comb;
  assign p2_add_92730_comb = p1_smul_89923 + p1_smul_89924;
  assign p2_add_93117_comb = p2_add_92731_comb + p2_add_92732_comb;
  assign p2_add_92725_comb = p2_add_92519_comb + p2_add_92520_comb;
  assign p2_add_92726_comb = p1_smul_89917 + p1_smul_89918;
  assign p2_add_93116_comb = p2_add_92727_comb + p2_add_92728_comb;
  assign p2_add_92721_comb = p2_add_92517_comb + p2_add_92518_comb;
  assign p2_add_92722_comb = p1_smul_89911 + p1_smul_89912;
  assign p2_add_93115_comb = p2_add_92723_comb + p2_add_92724_comb;
  assign p2_add_92717_comb = p2_add_92515_comb + p2_add_92516_comb;
  assign p2_add_92718_comb = p1_smul_89905 + p1_smul_89906;
  assign p2_add_93114_comb = p2_add_92719_comb + p2_add_92720_comb;
  assign p2_add_92713_comb = p2_add_92513_comb + p2_add_92514_comb;
  assign p2_add_92714_comb = p1_smul_89899 + p1_smul_89900;
  assign p2_add_93113_comb = p2_add_92715_comb + p2_add_92716_comb;

  // Registers for pipe stage 2:
  reg [31:0] p2_add_93109;
  reg [31:0] p2_add_93110;
  reg [31:0] p2_add_93212;
  reg [31:0] p2_add_93105;
  reg [31:0] p2_add_93106;
  reg [31:0] p2_add_93211;
  reg [31:0] p2_add_93101;
  reg [31:0] p2_add_93102;
  reg [31:0] p2_add_93210;
  reg [31:0] p2_add_93097;
  reg [31:0] p2_add_93098;
  reg [31:0] p2_add_93209;
  reg [31:0] p2_add_93093;
  reg [31:0] p2_add_93094;
  reg [31:0] p2_add_93208;
  reg [31:0] p2_add_93089;
  reg [31:0] p2_add_93090;
  reg [31:0] p2_add_93207;
  reg [31:0] p2_add_93085;
  reg [31:0] p2_add_93086;
  reg [31:0] p2_add_93206;
  reg [31:0] p2_add_93081;
  reg [31:0] p2_add_93082;
  reg [31:0] p2_add_93205;
  reg [31:0] p2_add_93077;
  reg [31:0] p2_add_93078;
  reg [31:0] p2_add_93204;
  reg [31:0] p2_add_93073;
  reg [31:0] p2_add_93074;
  reg [31:0] p2_add_93203;
  reg [31:0] p2_add_93069;
  reg [31:0] p2_add_93070;
  reg [31:0] p2_add_93202;
  reg [31:0] p2_add_93065;
  reg [31:0] p2_add_93066;
  reg [31:0] p2_add_93201;
  reg [31:0] p2_add_93061;
  reg [31:0] p2_add_93062;
  reg [31:0] p2_add_93200;
  reg [31:0] p2_add_93057;
  reg [31:0] p2_add_93058;
  reg [31:0] p2_add_93199;
  reg [31:0] p2_add_93053;
  reg [31:0] p2_add_93054;
  reg [31:0] p2_add_93198;
  reg [31:0] p2_add_93049;
  reg [31:0] p2_add_93050;
  reg [31:0] p2_add_93197;
  reg [31:0] p2_add_93045;
  reg [31:0] p2_add_93046;
  reg [31:0] p2_add_93196;
  reg [31:0] p2_add_93041;
  reg [31:0] p2_add_93042;
  reg [31:0] p2_add_93195;
  reg [31:0] p2_add_93037;
  reg [31:0] p2_add_93038;
  reg [31:0] p2_add_93194;
  reg [31:0] p2_add_93033;
  reg [31:0] p2_add_93034;
  reg [31:0] p2_add_93193;
  reg [31:0] p2_add_93029;
  reg [31:0] p2_add_93030;
  reg [31:0] p2_add_93192;
  reg [31:0] p2_add_93025;
  reg [31:0] p2_add_93026;
  reg [31:0] p2_add_93191;
  reg [31:0] p2_add_93021;
  reg [31:0] p2_add_93022;
  reg [31:0] p2_add_93190;
  reg [31:0] p2_add_93017;
  reg [31:0] p2_add_93018;
  reg [31:0] p2_add_93189;
  reg [31:0] p2_add_93013;
  reg [31:0] p2_add_93014;
  reg [31:0] p2_add_93188;
  reg [31:0] p2_add_93009;
  reg [31:0] p2_add_93010;
  reg [31:0] p2_add_93187;
  reg [31:0] p2_add_93005;
  reg [31:0] p2_add_93006;
  reg [31:0] p2_add_93186;
  reg [31:0] p2_add_93001;
  reg [31:0] p2_add_93002;
  reg [31:0] p2_add_93185;
  reg [31:0] p2_add_92997;
  reg [31:0] p2_add_92998;
  reg [31:0] p2_add_93184;
  reg [31:0] p2_add_92993;
  reg [31:0] p2_add_92994;
  reg [31:0] p2_add_93183;
  reg [31:0] p2_add_92989;
  reg [31:0] p2_add_92990;
  reg [31:0] p2_add_93182;
  reg [31:0] p2_add_92985;
  reg [31:0] p2_add_92986;
  reg [31:0] p2_add_93181;
  reg [31:0] p2_add_92981;
  reg [31:0] p2_add_92982;
  reg [31:0] p2_add_93180;
  reg [31:0] p2_add_92977;
  reg [31:0] p2_add_92978;
  reg [31:0] p2_add_93179;
  reg [31:0] p2_add_92973;
  reg [31:0] p2_add_92974;
  reg [31:0] p2_add_93178;
  reg [31:0] p2_add_92969;
  reg [31:0] p2_add_92970;
  reg [31:0] p2_add_93177;
  reg [31:0] p2_add_92965;
  reg [31:0] p2_add_92966;
  reg [31:0] p2_add_93176;
  reg [31:0] p2_add_92961;
  reg [31:0] p2_add_92962;
  reg [31:0] p2_add_93175;
  reg [31:0] p2_add_92957;
  reg [31:0] p2_add_92958;
  reg [31:0] p2_add_93174;
  reg [31:0] p2_add_92953;
  reg [31:0] p2_add_92954;
  reg [31:0] p2_add_93173;
  reg [31:0] p2_add_92949;
  reg [31:0] p2_add_92950;
  reg [31:0] p2_add_93172;
  reg [31:0] p2_add_92945;
  reg [31:0] p2_add_92946;
  reg [31:0] p2_add_93171;
  reg [31:0] p2_add_92941;
  reg [31:0] p2_add_92942;
  reg [31:0] p2_add_93170;
  reg [31:0] p2_add_92937;
  reg [31:0] p2_add_92938;
  reg [31:0] p2_add_93169;
  reg [31:0] p2_add_92933;
  reg [31:0] p2_add_92934;
  reg [31:0] p2_add_93168;
  reg [31:0] p2_add_92929;
  reg [31:0] p2_add_92930;
  reg [31:0] p2_add_93167;
  reg [31:0] p2_add_92925;
  reg [31:0] p2_add_92926;
  reg [31:0] p2_add_93166;
  reg [31:0] p2_add_92921;
  reg [31:0] p2_add_92922;
  reg [31:0] p2_add_93165;
  reg [31:0] p2_add_92917;
  reg [31:0] p2_add_92918;
  reg [31:0] p2_add_93164;
  reg [31:0] p2_add_92913;
  reg [31:0] p2_add_92914;
  reg [31:0] p2_add_93163;
  reg [31:0] p2_add_92909;
  reg [31:0] p2_add_92910;
  reg [31:0] p2_add_93162;
  reg [31:0] p2_add_92905;
  reg [31:0] p2_add_92906;
  reg [31:0] p2_add_93161;
  reg [31:0] p2_add_92901;
  reg [31:0] p2_add_92902;
  reg [31:0] p2_add_93160;
  reg [31:0] p2_add_92897;
  reg [31:0] p2_add_92898;
  reg [31:0] p2_add_93159;
  reg [31:0] p2_add_92893;
  reg [31:0] p2_add_92894;
  reg [31:0] p2_add_93158;
  reg [31:0] p2_add_92889;
  reg [31:0] p2_add_92890;
  reg [31:0] p2_add_93157;
  reg [31:0] p2_add_92885;
  reg [31:0] p2_add_92886;
  reg [31:0] p2_add_93156;
  reg [31:0] p2_add_92881;
  reg [31:0] p2_add_92882;
  reg [31:0] p2_add_93155;
  reg [31:0] p2_add_92877;
  reg [31:0] p2_add_92878;
  reg [31:0] p2_add_93154;
  reg [31:0] p2_add_92873;
  reg [31:0] p2_add_92874;
  reg [31:0] p2_add_93153;
  reg [31:0] p2_add_92869;
  reg [31:0] p2_add_92870;
  reg [31:0] p2_add_93152;
  reg [31:0] p2_add_92865;
  reg [31:0] p2_add_92866;
  reg [31:0] p2_add_93151;
  reg [31:0] p2_add_92861;
  reg [31:0] p2_add_92862;
  reg [31:0] p2_add_93150;
  reg [31:0] p2_add_92857;
  reg [31:0] p2_add_92858;
  reg [31:0] p2_add_93149;
  reg [31:0] p2_add_92853;
  reg [31:0] p2_add_92854;
  reg [31:0] p2_add_93148;
  reg [31:0] p2_add_92849;
  reg [31:0] p2_add_92850;
  reg [31:0] p2_add_93147;
  reg [31:0] p2_add_92845;
  reg [31:0] p2_add_92846;
  reg [31:0] p2_add_93146;
  reg [31:0] p2_add_92841;
  reg [31:0] p2_add_92842;
  reg [31:0] p2_add_93145;
  reg [31:0] p2_add_92837;
  reg [31:0] p2_add_92838;
  reg [31:0] p2_add_93144;
  reg [31:0] p2_add_92833;
  reg [31:0] p2_add_92834;
  reg [31:0] p2_add_93143;
  reg [31:0] p2_add_92829;
  reg [31:0] p2_add_92830;
  reg [31:0] p2_add_93142;
  reg [31:0] p2_add_92825;
  reg [31:0] p2_add_92826;
  reg [31:0] p2_add_93141;
  reg [31:0] p2_add_92821;
  reg [31:0] p2_add_92822;
  reg [31:0] p2_add_93140;
  reg [31:0] p2_add_92817;
  reg [31:0] p2_add_92818;
  reg [31:0] p2_add_93139;
  reg [31:0] p2_add_92813;
  reg [31:0] p2_add_92814;
  reg [31:0] p2_add_93138;
  reg [31:0] p2_add_92809;
  reg [31:0] p2_add_92810;
  reg [31:0] p2_add_93137;
  reg [31:0] p2_add_92805;
  reg [31:0] p2_add_92806;
  reg [31:0] p2_add_93136;
  reg [31:0] p2_add_92801;
  reg [31:0] p2_add_92802;
  reg [31:0] p2_add_93135;
  reg [31:0] p2_add_92797;
  reg [31:0] p2_add_92798;
  reg [31:0] p2_add_93134;
  reg [31:0] p2_add_92793;
  reg [31:0] p2_add_92794;
  reg [31:0] p2_add_93133;
  reg [31:0] p2_add_92789;
  reg [31:0] p2_add_92790;
  reg [31:0] p2_add_93132;
  reg [31:0] p2_add_92785;
  reg [31:0] p2_add_92786;
  reg [31:0] p2_add_93131;
  reg [31:0] p2_add_92781;
  reg [31:0] p2_add_92782;
  reg [31:0] p2_add_93130;
  reg [31:0] p2_add_92777;
  reg [31:0] p2_add_92778;
  reg [31:0] p2_add_93129;
  reg [31:0] p2_add_92773;
  reg [31:0] p2_add_92774;
  reg [31:0] p2_add_93128;
  reg [31:0] p2_add_92769;
  reg [31:0] p2_add_92770;
  reg [31:0] p2_add_93127;
  reg [31:0] p2_add_92765;
  reg [31:0] p2_add_92766;
  reg [31:0] p2_add_93126;
  reg [31:0] p2_add_92761;
  reg [31:0] p2_add_92762;
  reg [31:0] p2_add_93125;
  reg [31:0] p2_add_92757;
  reg [31:0] p2_add_92758;
  reg [31:0] p2_add_93124;
  reg [31:0] p2_add_92753;
  reg [31:0] p2_add_92754;
  reg [31:0] p2_add_93123;
  reg [31:0] p2_add_92749;
  reg [31:0] p2_add_92750;
  reg [31:0] p2_add_93122;
  reg [31:0] p2_add_92745;
  reg [31:0] p2_add_92746;
  reg [31:0] p2_add_93121;
  reg [31:0] p2_add_92741;
  reg [31:0] p2_add_92742;
  reg [31:0] p2_add_93120;
  reg [31:0] p2_add_92737;
  reg [31:0] p2_add_92738;
  reg [31:0] p2_add_93119;
  reg [31:0] p2_add_92733;
  reg [31:0] p2_add_92734;
  reg [31:0] p2_add_93118;
  reg [31:0] p2_add_92729;
  reg [31:0] p2_add_92730;
  reg [31:0] p2_add_93117;
  reg [31:0] p2_add_92725;
  reg [31:0] p2_add_92726;
  reg [31:0] p2_add_93116;
  reg [31:0] p2_add_92721;
  reg [31:0] p2_add_92722;
  reg [31:0] p2_add_93115;
  reg [31:0] p2_add_92717;
  reg [31:0] p2_add_92718;
  reg [31:0] p2_add_93114;
  reg [31:0] p2_add_92713;
  reg [31:0] p2_add_92714;
  reg [31:0] p2_add_93113;
  always_ff @ (posedge clk) begin
    p2_add_93109 <= p2_add_93109_comb;
    p2_add_93110 <= p2_add_93110_comb;
    p2_add_93212 <= p2_add_93212_comb;
    p2_add_93105 <= p2_add_93105_comb;
    p2_add_93106 <= p2_add_93106_comb;
    p2_add_93211 <= p2_add_93211_comb;
    p2_add_93101 <= p2_add_93101_comb;
    p2_add_93102 <= p2_add_93102_comb;
    p2_add_93210 <= p2_add_93210_comb;
    p2_add_93097 <= p2_add_93097_comb;
    p2_add_93098 <= p2_add_93098_comb;
    p2_add_93209 <= p2_add_93209_comb;
    p2_add_93093 <= p2_add_93093_comb;
    p2_add_93094 <= p2_add_93094_comb;
    p2_add_93208 <= p2_add_93208_comb;
    p2_add_93089 <= p2_add_93089_comb;
    p2_add_93090 <= p2_add_93090_comb;
    p2_add_93207 <= p2_add_93207_comb;
    p2_add_93085 <= p2_add_93085_comb;
    p2_add_93086 <= p2_add_93086_comb;
    p2_add_93206 <= p2_add_93206_comb;
    p2_add_93081 <= p2_add_93081_comb;
    p2_add_93082 <= p2_add_93082_comb;
    p2_add_93205 <= p2_add_93205_comb;
    p2_add_93077 <= p2_add_93077_comb;
    p2_add_93078 <= p2_add_93078_comb;
    p2_add_93204 <= p2_add_93204_comb;
    p2_add_93073 <= p2_add_93073_comb;
    p2_add_93074 <= p2_add_93074_comb;
    p2_add_93203 <= p2_add_93203_comb;
    p2_add_93069 <= p2_add_93069_comb;
    p2_add_93070 <= p2_add_93070_comb;
    p2_add_93202 <= p2_add_93202_comb;
    p2_add_93065 <= p2_add_93065_comb;
    p2_add_93066 <= p2_add_93066_comb;
    p2_add_93201 <= p2_add_93201_comb;
    p2_add_93061 <= p2_add_93061_comb;
    p2_add_93062 <= p2_add_93062_comb;
    p2_add_93200 <= p2_add_93200_comb;
    p2_add_93057 <= p2_add_93057_comb;
    p2_add_93058 <= p2_add_93058_comb;
    p2_add_93199 <= p2_add_93199_comb;
    p2_add_93053 <= p2_add_93053_comb;
    p2_add_93054 <= p2_add_93054_comb;
    p2_add_93198 <= p2_add_93198_comb;
    p2_add_93049 <= p2_add_93049_comb;
    p2_add_93050 <= p2_add_93050_comb;
    p2_add_93197 <= p2_add_93197_comb;
    p2_add_93045 <= p2_add_93045_comb;
    p2_add_93046 <= p2_add_93046_comb;
    p2_add_93196 <= p2_add_93196_comb;
    p2_add_93041 <= p2_add_93041_comb;
    p2_add_93042 <= p2_add_93042_comb;
    p2_add_93195 <= p2_add_93195_comb;
    p2_add_93037 <= p2_add_93037_comb;
    p2_add_93038 <= p2_add_93038_comb;
    p2_add_93194 <= p2_add_93194_comb;
    p2_add_93033 <= p2_add_93033_comb;
    p2_add_93034 <= p2_add_93034_comb;
    p2_add_93193 <= p2_add_93193_comb;
    p2_add_93029 <= p2_add_93029_comb;
    p2_add_93030 <= p2_add_93030_comb;
    p2_add_93192 <= p2_add_93192_comb;
    p2_add_93025 <= p2_add_93025_comb;
    p2_add_93026 <= p2_add_93026_comb;
    p2_add_93191 <= p2_add_93191_comb;
    p2_add_93021 <= p2_add_93021_comb;
    p2_add_93022 <= p2_add_93022_comb;
    p2_add_93190 <= p2_add_93190_comb;
    p2_add_93017 <= p2_add_93017_comb;
    p2_add_93018 <= p2_add_93018_comb;
    p2_add_93189 <= p2_add_93189_comb;
    p2_add_93013 <= p2_add_93013_comb;
    p2_add_93014 <= p2_add_93014_comb;
    p2_add_93188 <= p2_add_93188_comb;
    p2_add_93009 <= p2_add_93009_comb;
    p2_add_93010 <= p2_add_93010_comb;
    p2_add_93187 <= p2_add_93187_comb;
    p2_add_93005 <= p2_add_93005_comb;
    p2_add_93006 <= p2_add_93006_comb;
    p2_add_93186 <= p2_add_93186_comb;
    p2_add_93001 <= p2_add_93001_comb;
    p2_add_93002 <= p2_add_93002_comb;
    p2_add_93185 <= p2_add_93185_comb;
    p2_add_92997 <= p2_add_92997_comb;
    p2_add_92998 <= p2_add_92998_comb;
    p2_add_93184 <= p2_add_93184_comb;
    p2_add_92993 <= p2_add_92993_comb;
    p2_add_92994 <= p2_add_92994_comb;
    p2_add_93183 <= p2_add_93183_comb;
    p2_add_92989 <= p2_add_92989_comb;
    p2_add_92990 <= p2_add_92990_comb;
    p2_add_93182 <= p2_add_93182_comb;
    p2_add_92985 <= p2_add_92985_comb;
    p2_add_92986 <= p2_add_92986_comb;
    p2_add_93181 <= p2_add_93181_comb;
    p2_add_92981 <= p2_add_92981_comb;
    p2_add_92982 <= p2_add_92982_comb;
    p2_add_93180 <= p2_add_93180_comb;
    p2_add_92977 <= p2_add_92977_comb;
    p2_add_92978 <= p2_add_92978_comb;
    p2_add_93179 <= p2_add_93179_comb;
    p2_add_92973 <= p2_add_92973_comb;
    p2_add_92974 <= p2_add_92974_comb;
    p2_add_93178 <= p2_add_93178_comb;
    p2_add_92969 <= p2_add_92969_comb;
    p2_add_92970 <= p2_add_92970_comb;
    p2_add_93177 <= p2_add_93177_comb;
    p2_add_92965 <= p2_add_92965_comb;
    p2_add_92966 <= p2_add_92966_comb;
    p2_add_93176 <= p2_add_93176_comb;
    p2_add_92961 <= p2_add_92961_comb;
    p2_add_92962 <= p2_add_92962_comb;
    p2_add_93175 <= p2_add_93175_comb;
    p2_add_92957 <= p2_add_92957_comb;
    p2_add_92958 <= p2_add_92958_comb;
    p2_add_93174 <= p2_add_93174_comb;
    p2_add_92953 <= p2_add_92953_comb;
    p2_add_92954 <= p2_add_92954_comb;
    p2_add_93173 <= p2_add_93173_comb;
    p2_add_92949 <= p2_add_92949_comb;
    p2_add_92950 <= p2_add_92950_comb;
    p2_add_93172 <= p2_add_93172_comb;
    p2_add_92945 <= p2_add_92945_comb;
    p2_add_92946 <= p2_add_92946_comb;
    p2_add_93171 <= p2_add_93171_comb;
    p2_add_92941 <= p2_add_92941_comb;
    p2_add_92942 <= p2_add_92942_comb;
    p2_add_93170 <= p2_add_93170_comb;
    p2_add_92937 <= p2_add_92937_comb;
    p2_add_92938 <= p2_add_92938_comb;
    p2_add_93169 <= p2_add_93169_comb;
    p2_add_92933 <= p2_add_92933_comb;
    p2_add_92934 <= p2_add_92934_comb;
    p2_add_93168 <= p2_add_93168_comb;
    p2_add_92929 <= p2_add_92929_comb;
    p2_add_92930 <= p2_add_92930_comb;
    p2_add_93167 <= p2_add_93167_comb;
    p2_add_92925 <= p2_add_92925_comb;
    p2_add_92926 <= p2_add_92926_comb;
    p2_add_93166 <= p2_add_93166_comb;
    p2_add_92921 <= p2_add_92921_comb;
    p2_add_92922 <= p2_add_92922_comb;
    p2_add_93165 <= p2_add_93165_comb;
    p2_add_92917 <= p2_add_92917_comb;
    p2_add_92918 <= p2_add_92918_comb;
    p2_add_93164 <= p2_add_93164_comb;
    p2_add_92913 <= p2_add_92913_comb;
    p2_add_92914 <= p2_add_92914_comb;
    p2_add_93163 <= p2_add_93163_comb;
    p2_add_92909 <= p2_add_92909_comb;
    p2_add_92910 <= p2_add_92910_comb;
    p2_add_93162 <= p2_add_93162_comb;
    p2_add_92905 <= p2_add_92905_comb;
    p2_add_92906 <= p2_add_92906_comb;
    p2_add_93161 <= p2_add_93161_comb;
    p2_add_92901 <= p2_add_92901_comb;
    p2_add_92902 <= p2_add_92902_comb;
    p2_add_93160 <= p2_add_93160_comb;
    p2_add_92897 <= p2_add_92897_comb;
    p2_add_92898 <= p2_add_92898_comb;
    p2_add_93159 <= p2_add_93159_comb;
    p2_add_92893 <= p2_add_92893_comb;
    p2_add_92894 <= p2_add_92894_comb;
    p2_add_93158 <= p2_add_93158_comb;
    p2_add_92889 <= p2_add_92889_comb;
    p2_add_92890 <= p2_add_92890_comb;
    p2_add_93157 <= p2_add_93157_comb;
    p2_add_92885 <= p2_add_92885_comb;
    p2_add_92886 <= p2_add_92886_comb;
    p2_add_93156 <= p2_add_93156_comb;
    p2_add_92881 <= p2_add_92881_comb;
    p2_add_92882 <= p2_add_92882_comb;
    p2_add_93155 <= p2_add_93155_comb;
    p2_add_92877 <= p2_add_92877_comb;
    p2_add_92878 <= p2_add_92878_comb;
    p2_add_93154 <= p2_add_93154_comb;
    p2_add_92873 <= p2_add_92873_comb;
    p2_add_92874 <= p2_add_92874_comb;
    p2_add_93153 <= p2_add_93153_comb;
    p2_add_92869 <= p2_add_92869_comb;
    p2_add_92870 <= p2_add_92870_comb;
    p2_add_93152 <= p2_add_93152_comb;
    p2_add_92865 <= p2_add_92865_comb;
    p2_add_92866 <= p2_add_92866_comb;
    p2_add_93151 <= p2_add_93151_comb;
    p2_add_92861 <= p2_add_92861_comb;
    p2_add_92862 <= p2_add_92862_comb;
    p2_add_93150 <= p2_add_93150_comb;
    p2_add_92857 <= p2_add_92857_comb;
    p2_add_92858 <= p2_add_92858_comb;
    p2_add_93149 <= p2_add_93149_comb;
    p2_add_92853 <= p2_add_92853_comb;
    p2_add_92854 <= p2_add_92854_comb;
    p2_add_93148 <= p2_add_93148_comb;
    p2_add_92849 <= p2_add_92849_comb;
    p2_add_92850 <= p2_add_92850_comb;
    p2_add_93147 <= p2_add_93147_comb;
    p2_add_92845 <= p2_add_92845_comb;
    p2_add_92846 <= p2_add_92846_comb;
    p2_add_93146 <= p2_add_93146_comb;
    p2_add_92841 <= p2_add_92841_comb;
    p2_add_92842 <= p2_add_92842_comb;
    p2_add_93145 <= p2_add_93145_comb;
    p2_add_92837 <= p2_add_92837_comb;
    p2_add_92838 <= p2_add_92838_comb;
    p2_add_93144 <= p2_add_93144_comb;
    p2_add_92833 <= p2_add_92833_comb;
    p2_add_92834 <= p2_add_92834_comb;
    p2_add_93143 <= p2_add_93143_comb;
    p2_add_92829 <= p2_add_92829_comb;
    p2_add_92830 <= p2_add_92830_comb;
    p2_add_93142 <= p2_add_93142_comb;
    p2_add_92825 <= p2_add_92825_comb;
    p2_add_92826 <= p2_add_92826_comb;
    p2_add_93141 <= p2_add_93141_comb;
    p2_add_92821 <= p2_add_92821_comb;
    p2_add_92822 <= p2_add_92822_comb;
    p2_add_93140 <= p2_add_93140_comb;
    p2_add_92817 <= p2_add_92817_comb;
    p2_add_92818 <= p2_add_92818_comb;
    p2_add_93139 <= p2_add_93139_comb;
    p2_add_92813 <= p2_add_92813_comb;
    p2_add_92814 <= p2_add_92814_comb;
    p2_add_93138 <= p2_add_93138_comb;
    p2_add_92809 <= p2_add_92809_comb;
    p2_add_92810 <= p2_add_92810_comb;
    p2_add_93137 <= p2_add_93137_comb;
    p2_add_92805 <= p2_add_92805_comb;
    p2_add_92806 <= p2_add_92806_comb;
    p2_add_93136 <= p2_add_93136_comb;
    p2_add_92801 <= p2_add_92801_comb;
    p2_add_92802 <= p2_add_92802_comb;
    p2_add_93135 <= p2_add_93135_comb;
    p2_add_92797 <= p2_add_92797_comb;
    p2_add_92798 <= p2_add_92798_comb;
    p2_add_93134 <= p2_add_93134_comb;
    p2_add_92793 <= p2_add_92793_comb;
    p2_add_92794 <= p2_add_92794_comb;
    p2_add_93133 <= p2_add_93133_comb;
    p2_add_92789 <= p2_add_92789_comb;
    p2_add_92790 <= p2_add_92790_comb;
    p2_add_93132 <= p2_add_93132_comb;
    p2_add_92785 <= p2_add_92785_comb;
    p2_add_92786 <= p2_add_92786_comb;
    p2_add_93131 <= p2_add_93131_comb;
    p2_add_92781 <= p2_add_92781_comb;
    p2_add_92782 <= p2_add_92782_comb;
    p2_add_93130 <= p2_add_93130_comb;
    p2_add_92777 <= p2_add_92777_comb;
    p2_add_92778 <= p2_add_92778_comb;
    p2_add_93129 <= p2_add_93129_comb;
    p2_add_92773 <= p2_add_92773_comb;
    p2_add_92774 <= p2_add_92774_comb;
    p2_add_93128 <= p2_add_93128_comb;
    p2_add_92769 <= p2_add_92769_comb;
    p2_add_92770 <= p2_add_92770_comb;
    p2_add_93127 <= p2_add_93127_comb;
    p2_add_92765 <= p2_add_92765_comb;
    p2_add_92766 <= p2_add_92766_comb;
    p2_add_93126 <= p2_add_93126_comb;
    p2_add_92761 <= p2_add_92761_comb;
    p2_add_92762 <= p2_add_92762_comb;
    p2_add_93125 <= p2_add_93125_comb;
    p2_add_92757 <= p2_add_92757_comb;
    p2_add_92758 <= p2_add_92758_comb;
    p2_add_93124 <= p2_add_93124_comb;
    p2_add_92753 <= p2_add_92753_comb;
    p2_add_92754 <= p2_add_92754_comb;
    p2_add_93123 <= p2_add_93123_comb;
    p2_add_92749 <= p2_add_92749_comb;
    p2_add_92750 <= p2_add_92750_comb;
    p2_add_93122 <= p2_add_93122_comb;
    p2_add_92745 <= p2_add_92745_comb;
    p2_add_92746 <= p2_add_92746_comb;
    p2_add_93121 <= p2_add_93121_comb;
    p2_add_92741 <= p2_add_92741_comb;
    p2_add_92742 <= p2_add_92742_comb;
    p2_add_93120 <= p2_add_93120_comb;
    p2_add_92737 <= p2_add_92737_comb;
    p2_add_92738 <= p2_add_92738_comb;
    p2_add_93119 <= p2_add_93119_comb;
    p2_add_92733 <= p2_add_92733_comb;
    p2_add_92734 <= p2_add_92734_comb;
    p2_add_93118 <= p2_add_93118_comb;
    p2_add_92729 <= p2_add_92729_comb;
    p2_add_92730 <= p2_add_92730_comb;
    p2_add_93117 <= p2_add_93117_comb;
    p2_add_92725 <= p2_add_92725_comb;
    p2_add_92726 <= p2_add_92726_comb;
    p2_add_93116 <= p2_add_93116_comb;
    p2_add_92721 <= p2_add_92721_comb;
    p2_add_92722 <= p2_add_92722_comb;
    p2_add_93115 <= p2_add_93115_comb;
    p2_add_92717 <= p2_add_92717_comb;
    p2_add_92718 <= p2_add_92718_comb;
    p2_add_93114 <= p2_add_93114_comb;
    p2_add_92713 <= p2_add_92713_comb;
    p2_add_92714 <= p2_add_92714_comb;
    p2_add_93113 <= p2_add_93113_comb;
  end

  // ===== Pipe stage 3:
  wire [31:0] p3_add_93925_comb;
  wire [31:0] p3_add_93924_comb;
  wire [31:0] p3_add_93923_comb;
  wire [31:0] p3_add_93922_comb;
  wire [31:0] p3_add_93921_comb;
  wire [31:0] p3_add_93920_comb;
  wire [31:0] p3_add_93919_comb;
  wire [31:0] p3_add_93918_comb;
  wire [31:0] p3_add_93917_comb;
  wire [31:0] p3_add_93916_comb;
  wire [31:0] p3_add_93915_comb;
  wire [31:0] p3_add_93914_comb;
  wire [31:0] p3_add_93913_comb;
  wire [31:0] p3_add_93912_comb;
  wire [31:0] p3_add_93911_comb;
  wire [31:0] p3_add_93910_comb;
  wire [31:0] p3_add_93909_comb;
  wire [31:0] p3_add_93908_comb;
  wire [31:0] p3_add_93907_comb;
  wire [31:0] p3_add_93906_comb;
  wire [31:0] p3_add_93905_comb;
  wire [31:0] p3_add_93904_comb;
  wire [31:0] p3_add_93903_comb;
  wire [31:0] p3_add_93902_comb;
  wire [31:0] p3_add_93901_comb;
  wire [31:0] p3_add_93900_comb;
  wire [31:0] p3_add_93899_comb;
  wire [31:0] p3_add_93898_comb;
  wire [31:0] p3_add_93897_comb;
  wire [31:0] p3_add_93896_comb;
  wire [31:0] p3_add_93895_comb;
  wire [31:0] p3_add_93894_comb;
  wire [31:0] p3_add_93893_comb;
  wire [31:0] p3_add_93892_comb;
  wire [31:0] p3_add_93891_comb;
  wire [31:0] p3_add_93890_comb;
  wire [31:0] p3_add_93889_comb;
  wire [31:0] p3_add_93888_comb;
  wire [31:0] p3_add_93887_comb;
  wire [31:0] p3_add_93886_comb;
  wire [31:0] p3_add_93885_comb;
  wire [31:0] p3_add_93884_comb;
  wire [31:0] p3_add_93883_comb;
  wire [31:0] p3_add_93882_comb;
  wire [31:0] p3_add_93881_comb;
  wire [31:0] p3_add_93880_comb;
  wire [31:0] p3_add_93879_comb;
  wire [31:0] p3_add_93878_comb;
  wire [31:0] p3_add_93877_comb;
  wire [31:0] p3_add_93876_comb;
  wire [31:0] p3_add_93875_comb;
  wire [31:0] p3_add_93874_comb;
  wire [31:0] p3_add_93873_comb;
  wire [31:0] p3_add_93872_comb;
  wire [31:0] p3_add_93871_comb;
  wire [31:0] p3_add_93870_comb;
  wire [31:0] p3_add_93869_comb;
  wire [31:0] p3_add_93868_comb;
  wire [31:0] p3_add_93867_comb;
  wire [31:0] p3_add_93866_comb;
  wire [31:0] p3_add_93865_comb;
  wire [31:0] p3_add_93864_comb;
  wire [31:0] p3_add_93863_comb;
  wire [31:0] p3_add_93862_comb;
  wire [31:0] p3_add_93861_comb;
  wire [31:0] p3_add_93860_comb;
  wire [31:0] p3_add_93859_comb;
  wire [31:0] p3_add_93858_comb;
  wire [31:0] p3_add_93857_comb;
  wire [31:0] p3_add_93856_comb;
  wire [31:0] p3_add_93855_comb;
  wire [31:0] p3_add_93854_comb;
  wire [31:0] p3_add_93853_comb;
  wire [31:0] p3_add_93852_comb;
  wire [31:0] p3_add_93851_comb;
  wire [31:0] p3_add_93850_comb;
  wire [31:0] p3_add_93849_comb;
  wire [31:0] p3_add_93848_comb;
  wire [31:0] p3_add_93847_comb;
  wire [31:0] p3_add_93846_comb;
  wire [31:0] p3_add_93845_comb;
  wire [31:0] p3_add_93844_comb;
  wire [31:0] p3_add_93843_comb;
  wire [31:0] p3_add_93842_comb;
  wire [31:0] p3_add_93841_comb;
  wire [31:0] p3_add_93840_comb;
  wire [31:0] p3_add_93839_comb;
  wire [31:0] p3_add_93838_comb;
  wire [31:0] p3_add_93837_comb;
  wire [31:0] p3_add_93836_comb;
  wire [31:0] p3_add_93835_comb;
  wire [31:0] p3_add_93834_comb;
  wire [31:0] p3_add_93833_comb;
  wire [31:0] p3_add_93832_comb;
  wire [31:0] p3_add_93831_comb;
  wire [31:0] p3_add_93830_comb;
  wire [31:0] p3_add_93829_comb;
  wire [31:0] p3_add_93828_comb;
  wire [31:0] p3_add_93827_comb;
  wire [31:0] p3_add_93826_comb;
  wire [31:0] p3_add_94025_comb;
  wire [31:0] p3_add_94024_comb;
  wire [31:0] p3_add_94023_comb;
  wire [31:0] p3_add_94022_comb;
  wire [31:0] p3_add_94021_comb;
  wire [31:0] p3_add_94020_comb;
  wire [31:0] p3_add_94019_comb;
  wire [31:0] p3_add_94018_comb;
  wire [31:0] p3_add_94017_comb;
  wire [31:0] p3_add_94016_comb;
  wire [31:0] p3_add_94015_comb;
  wire [31:0] p3_add_94014_comb;
  wire [31:0] p3_add_94013_comb;
  wire [31:0] p3_add_94012_comb;
  wire [31:0] p3_add_94011_comb;
  wire [31:0] p3_add_94010_comb;
  wire [31:0] p3_add_94009_comb;
  wire [31:0] p3_add_94008_comb;
  wire [31:0] p3_add_94007_comb;
  wire [31:0] p3_add_94006_comb;
  wire [31:0] p3_add_94005_comb;
  wire [31:0] p3_add_94004_comb;
  wire [31:0] p3_add_94003_comb;
  wire [31:0] p3_add_94002_comb;
  wire [31:0] p3_add_94001_comb;
  wire [31:0] p3_add_94000_comb;
  wire [31:0] p3_add_93999_comb;
  wire [31:0] p3_add_93998_comb;
  wire [31:0] p3_add_93997_comb;
  wire [31:0] p3_add_93996_comb;
  wire [31:0] p3_add_93995_comb;
  wire [31:0] p3_add_93994_comb;
  wire [31:0] p3_add_93993_comb;
  wire [31:0] p3_add_93992_comb;
  wire [31:0] p3_add_93991_comb;
  wire [31:0] p3_add_93990_comb;
  wire [31:0] p3_add_93989_comb;
  wire [31:0] p3_add_93988_comb;
  wire [31:0] p3_add_93987_comb;
  wire [31:0] p3_add_93986_comb;
  wire [31:0] p3_add_93985_comb;
  wire [31:0] p3_add_93984_comb;
  wire [31:0] p3_add_93983_comb;
  wire [31:0] p3_add_93982_comb;
  wire [31:0] p3_add_93981_comb;
  wire [31:0] p3_add_93980_comb;
  wire [31:0] p3_add_93979_comb;
  wire [31:0] p3_add_93978_comb;
  wire [31:0] p3_add_93977_comb;
  wire [31:0] p3_add_93976_comb;
  wire [31:0] p3_add_93975_comb;
  wire [31:0] p3_add_93974_comb;
  wire [31:0] p3_add_93973_comb;
  wire [31:0] p3_add_93972_comb;
  wire [31:0] p3_add_93971_comb;
  wire [31:0] p3_add_93970_comb;
  wire [31:0] p3_add_93969_comb;
  wire [31:0] p3_add_93968_comb;
  wire [31:0] p3_add_93967_comb;
  wire [31:0] p3_add_93966_comb;
  wire [31:0] p3_add_93965_comb;
  wire [31:0] p3_add_93964_comb;
  wire [31:0] p3_add_93963_comb;
  wire [31:0] p3_add_93962_comb;
  wire [31:0] p3_add_93961_comb;
  wire [31:0] p3_add_93960_comb;
  wire [31:0] p3_add_93959_comb;
  wire [31:0] p3_add_93958_comb;
  wire [31:0] p3_add_93957_comb;
  wire [31:0] p3_add_93956_comb;
  wire [31:0] p3_add_93955_comb;
  wire [31:0] p3_add_93954_comb;
  wire [31:0] p3_add_93953_comb;
  wire [31:0] p3_add_93952_comb;
  wire [31:0] p3_add_93951_comb;
  wire [31:0] p3_add_93950_comb;
  wire [31:0] p3_add_93949_comb;
  wire [31:0] p3_add_93948_comb;
  wire [31:0] p3_add_93947_comb;
  wire [31:0] p3_add_93946_comb;
  wire [31:0] p3_add_93945_comb;
  wire [31:0] p3_add_93944_comb;
  wire [31:0] p3_add_93943_comb;
  wire [31:0] p3_add_93942_comb;
  wire [31:0] p3_add_93941_comb;
  wire [31:0] p3_add_93940_comb;
  wire [31:0] p3_add_93939_comb;
  wire [31:0] p3_add_93938_comb;
  wire [31:0] p3_add_93937_comb;
  wire [31:0] p3_add_93936_comb;
  wire [31:0] p3_add_93935_comb;
  wire [31:0] p3_add_93934_comb;
  wire [31:0] p3_add_93933_comb;
  wire [31:0] p3_add_93932_comb;
  wire [31:0] p3_add_93931_comb;
  wire [31:0] p3_add_93930_comb;
  wire [31:0] p3_add_93929_comb;
  wire [31:0] p3_add_93928_comb;
  wire [31:0] p3_add_93927_comb;
  wire [31:0] p3_add_93926_comb;
  assign p3_add_93925_comb = p2_add_93109 + p2_add_93110;
  assign p3_add_93924_comb = p2_add_93105 + p2_add_93106;
  assign p3_add_93923_comb = p2_add_93101 + p2_add_93102;
  assign p3_add_93922_comb = p2_add_93097 + p2_add_93098;
  assign p3_add_93921_comb = p2_add_93093 + p2_add_93094;
  assign p3_add_93920_comb = p2_add_93089 + p2_add_93090;
  assign p3_add_93919_comb = p2_add_93085 + p2_add_93086;
  assign p3_add_93918_comb = p2_add_93081 + p2_add_93082;
  assign p3_add_93917_comb = p2_add_93077 + p2_add_93078;
  assign p3_add_93916_comb = p2_add_93073 + p2_add_93074;
  assign p3_add_93915_comb = p2_add_93069 + p2_add_93070;
  assign p3_add_93914_comb = p2_add_93065 + p2_add_93066;
  assign p3_add_93913_comb = p2_add_93061 + p2_add_93062;
  assign p3_add_93912_comb = p2_add_93057 + p2_add_93058;
  assign p3_add_93911_comb = p2_add_93053 + p2_add_93054;
  assign p3_add_93910_comb = p2_add_93049 + p2_add_93050;
  assign p3_add_93909_comb = p2_add_93045 + p2_add_93046;
  assign p3_add_93908_comb = p2_add_93041 + p2_add_93042;
  assign p3_add_93907_comb = p2_add_93037 + p2_add_93038;
  assign p3_add_93906_comb = p2_add_93033 + p2_add_93034;
  assign p3_add_93905_comb = p2_add_93029 + p2_add_93030;
  assign p3_add_93904_comb = p2_add_93025 + p2_add_93026;
  assign p3_add_93903_comb = p2_add_93021 + p2_add_93022;
  assign p3_add_93902_comb = p2_add_93017 + p2_add_93018;
  assign p3_add_93901_comb = p2_add_93013 + p2_add_93014;
  assign p3_add_93900_comb = p2_add_93009 + p2_add_93010;
  assign p3_add_93899_comb = p2_add_93005 + p2_add_93006;
  assign p3_add_93898_comb = p2_add_93001 + p2_add_93002;
  assign p3_add_93897_comb = p2_add_92997 + p2_add_92998;
  assign p3_add_93896_comb = p2_add_92993 + p2_add_92994;
  assign p3_add_93895_comb = p2_add_92989 + p2_add_92990;
  assign p3_add_93894_comb = p2_add_92985 + p2_add_92986;
  assign p3_add_93893_comb = p2_add_92981 + p2_add_92982;
  assign p3_add_93892_comb = p2_add_92977 + p2_add_92978;
  assign p3_add_93891_comb = p2_add_92973 + p2_add_92974;
  assign p3_add_93890_comb = p2_add_92969 + p2_add_92970;
  assign p3_add_93889_comb = p2_add_92965 + p2_add_92966;
  assign p3_add_93888_comb = p2_add_92961 + p2_add_92962;
  assign p3_add_93887_comb = p2_add_92957 + p2_add_92958;
  assign p3_add_93886_comb = p2_add_92953 + p2_add_92954;
  assign p3_add_93885_comb = p2_add_92949 + p2_add_92950;
  assign p3_add_93884_comb = p2_add_92945 + p2_add_92946;
  assign p3_add_93883_comb = p2_add_92941 + p2_add_92942;
  assign p3_add_93882_comb = p2_add_92937 + p2_add_92938;
  assign p3_add_93881_comb = p2_add_92933 + p2_add_92934;
  assign p3_add_93880_comb = p2_add_92929 + p2_add_92930;
  assign p3_add_93879_comb = p2_add_92925 + p2_add_92926;
  assign p3_add_93878_comb = p2_add_92921 + p2_add_92922;
  assign p3_add_93877_comb = p2_add_92917 + p2_add_92918;
  assign p3_add_93876_comb = p2_add_92913 + p2_add_92914;
  assign p3_add_93875_comb = p2_add_92909 + p2_add_92910;
  assign p3_add_93874_comb = p2_add_92905 + p2_add_92906;
  assign p3_add_93873_comb = p2_add_92901 + p2_add_92902;
  assign p3_add_93872_comb = p2_add_92897 + p2_add_92898;
  assign p3_add_93871_comb = p2_add_92893 + p2_add_92894;
  assign p3_add_93870_comb = p2_add_92889 + p2_add_92890;
  assign p3_add_93869_comb = p2_add_92885 + p2_add_92886;
  assign p3_add_93868_comb = p2_add_92881 + p2_add_92882;
  assign p3_add_93867_comb = p2_add_92877 + p2_add_92878;
  assign p3_add_93866_comb = p2_add_92873 + p2_add_92874;
  assign p3_add_93865_comb = p2_add_92869 + p2_add_92870;
  assign p3_add_93864_comb = p2_add_92865 + p2_add_92866;
  assign p3_add_93863_comb = p2_add_92861 + p2_add_92862;
  assign p3_add_93862_comb = p2_add_92857 + p2_add_92858;
  assign p3_add_93861_comb = p2_add_92853 + p2_add_92854;
  assign p3_add_93860_comb = p2_add_92849 + p2_add_92850;
  assign p3_add_93859_comb = p2_add_92845 + p2_add_92846;
  assign p3_add_93858_comb = p2_add_92841 + p2_add_92842;
  assign p3_add_93857_comb = p2_add_92837 + p2_add_92838;
  assign p3_add_93856_comb = p2_add_92833 + p2_add_92834;
  assign p3_add_93855_comb = p2_add_92829 + p2_add_92830;
  assign p3_add_93854_comb = p2_add_92825 + p2_add_92826;
  assign p3_add_93853_comb = p2_add_92821 + p2_add_92822;
  assign p3_add_93852_comb = p2_add_92817 + p2_add_92818;
  assign p3_add_93851_comb = p2_add_92813 + p2_add_92814;
  assign p3_add_93850_comb = p2_add_92809 + p2_add_92810;
  assign p3_add_93849_comb = p2_add_92805 + p2_add_92806;
  assign p3_add_93848_comb = p2_add_92801 + p2_add_92802;
  assign p3_add_93847_comb = p2_add_92797 + p2_add_92798;
  assign p3_add_93846_comb = p2_add_92793 + p2_add_92794;
  assign p3_add_93845_comb = p2_add_92789 + p2_add_92790;
  assign p3_add_93844_comb = p2_add_92785 + p2_add_92786;
  assign p3_add_93843_comb = p2_add_92781 + p2_add_92782;
  assign p3_add_93842_comb = p2_add_92777 + p2_add_92778;
  assign p3_add_93841_comb = p2_add_92773 + p2_add_92774;
  assign p3_add_93840_comb = p2_add_92769 + p2_add_92770;
  assign p3_add_93839_comb = p2_add_92765 + p2_add_92766;
  assign p3_add_93838_comb = p2_add_92761 + p2_add_92762;
  assign p3_add_93837_comb = p2_add_92757 + p2_add_92758;
  assign p3_add_93836_comb = p2_add_92753 + p2_add_92754;
  assign p3_add_93835_comb = p2_add_92749 + p2_add_92750;
  assign p3_add_93834_comb = p2_add_92745 + p2_add_92746;
  assign p3_add_93833_comb = p2_add_92741 + p2_add_92742;
  assign p3_add_93832_comb = p2_add_92737 + p2_add_92738;
  assign p3_add_93831_comb = p2_add_92733 + p2_add_92734;
  assign p3_add_93830_comb = p2_add_92729 + p2_add_92730;
  assign p3_add_93829_comb = p2_add_92725 + p2_add_92726;
  assign p3_add_93828_comb = p2_add_92721 + p2_add_92722;
  assign p3_add_93827_comb = p2_add_92717 + p2_add_92718;
  assign p3_add_93826_comb = p2_add_92713 + p2_add_92714;
  assign p3_add_94025_comb = p3_add_93925_comb + p2_add_93212;
  assign p3_add_94024_comb = p3_add_93924_comb + p2_add_93211;
  assign p3_add_94023_comb = p3_add_93923_comb + p2_add_93210;
  assign p3_add_94022_comb = p3_add_93922_comb + p2_add_93209;
  assign p3_add_94021_comb = p3_add_93921_comb + p2_add_93208;
  assign p3_add_94020_comb = p3_add_93920_comb + p2_add_93207;
  assign p3_add_94019_comb = p3_add_93919_comb + p2_add_93206;
  assign p3_add_94018_comb = p3_add_93918_comb + p2_add_93205;
  assign p3_add_94017_comb = p3_add_93917_comb + p2_add_93204;
  assign p3_add_94016_comb = p3_add_93916_comb + p2_add_93203;
  assign p3_add_94015_comb = p3_add_93915_comb + p2_add_93202;
  assign p3_add_94014_comb = p3_add_93914_comb + p2_add_93201;
  assign p3_add_94013_comb = p3_add_93913_comb + p2_add_93200;
  assign p3_add_94012_comb = p3_add_93912_comb + p2_add_93199;
  assign p3_add_94011_comb = p3_add_93911_comb + p2_add_93198;
  assign p3_add_94010_comb = p3_add_93910_comb + p2_add_93197;
  assign p3_add_94009_comb = p3_add_93909_comb + p2_add_93196;
  assign p3_add_94008_comb = p3_add_93908_comb + p2_add_93195;
  assign p3_add_94007_comb = p3_add_93907_comb + p2_add_93194;
  assign p3_add_94006_comb = p3_add_93906_comb + p2_add_93193;
  assign p3_add_94005_comb = p3_add_93905_comb + p2_add_93192;
  assign p3_add_94004_comb = p3_add_93904_comb + p2_add_93191;
  assign p3_add_94003_comb = p3_add_93903_comb + p2_add_93190;
  assign p3_add_94002_comb = p3_add_93902_comb + p2_add_93189;
  assign p3_add_94001_comb = p3_add_93901_comb + p2_add_93188;
  assign p3_add_94000_comb = p3_add_93900_comb + p2_add_93187;
  assign p3_add_93999_comb = p3_add_93899_comb + p2_add_93186;
  assign p3_add_93998_comb = p3_add_93898_comb + p2_add_93185;
  assign p3_add_93997_comb = p3_add_93897_comb + p2_add_93184;
  assign p3_add_93996_comb = p3_add_93896_comb + p2_add_93183;
  assign p3_add_93995_comb = p3_add_93895_comb + p2_add_93182;
  assign p3_add_93994_comb = p3_add_93894_comb + p2_add_93181;
  assign p3_add_93993_comb = p3_add_93893_comb + p2_add_93180;
  assign p3_add_93992_comb = p3_add_93892_comb + p2_add_93179;
  assign p3_add_93991_comb = p3_add_93891_comb + p2_add_93178;
  assign p3_add_93990_comb = p3_add_93890_comb + p2_add_93177;
  assign p3_add_93989_comb = p3_add_93889_comb + p2_add_93176;
  assign p3_add_93988_comb = p3_add_93888_comb + p2_add_93175;
  assign p3_add_93987_comb = p3_add_93887_comb + p2_add_93174;
  assign p3_add_93986_comb = p3_add_93886_comb + p2_add_93173;
  assign p3_add_93985_comb = p3_add_93885_comb + p2_add_93172;
  assign p3_add_93984_comb = p3_add_93884_comb + p2_add_93171;
  assign p3_add_93983_comb = p3_add_93883_comb + p2_add_93170;
  assign p3_add_93982_comb = p3_add_93882_comb + p2_add_93169;
  assign p3_add_93981_comb = p3_add_93881_comb + p2_add_93168;
  assign p3_add_93980_comb = p3_add_93880_comb + p2_add_93167;
  assign p3_add_93979_comb = p3_add_93879_comb + p2_add_93166;
  assign p3_add_93978_comb = p3_add_93878_comb + p2_add_93165;
  assign p3_add_93977_comb = p3_add_93877_comb + p2_add_93164;
  assign p3_add_93976_comb = p3_add_93876_comb + p2_add_93163;
  assign p3_add_93975_comb = p3_add_93875_comb + p2_add_93162;
  assign p3_add_93974_comb = p3_add_93874_comb + p2_add_93161;
  assign p3_add_93973_comb = p3_add_93873_comb + p2_add_93160;
  assign p3_add_93972_comb = p3_add_93872_comb + p2_add_93159;
  assign p3_add_93971_comb = p3_add_93871_comb + p2_add_93158;
  assign p3_add_93970_comb = p3_add_93870_comb + p2_add_93157;
  assign p3_add_93969_comb = p3_add_93869_comb + p2_add_93156;
  assign p3_add_93968_comb = p3_add_93868_comb + p2_add_93155;
  assign p3_add_93967_comb = p3_add_93867_comb + p2_add_93154;
  assign p3_add_93966_comb = p3_add_93866_comb + p2_add_93153;
  assign p3_add_93965_comb = p3_add_93865_comb + p2_add_93152;
  assign p3_add_93964_comb = p3_add_93864_comb + p2_add_93151;
  assign p3_add_93963_comb = p3_add_93863_comb + p2_add_93150;
  assign p3_add_93962_comb = p3_add_93862_comb + p2_add_93149;
  assign p3_add_93961_comb = p3_add_93861_comb + p2_add_93148;
  assign p3_add_93960_comb = p3_add_93860_comb + p2_add_93147;
  assign p3_add_93959_comb = p3_add_93859_comb + p2_add_93146;
  assign p3_add_93958_comb = p3_add_93858_comb + p2_add_93145;
  assign p3_add_93957_comb = p3_add_93857_comb + p2_add_93144;
  assign p3_add_93956_comb = p3_add_93856_comb + p2_add_93143;
  assign p3_add_93955_comb = p3_add_93855_comb + p2_add_93142;
  assign p3_add_93954_comb = p3_add_93854_comb + p2_add_93141;
  assign p3_add_93953_comb = p3_add_93853_comb + p2_add_93140;
  assign p3_add_93952_comb = p3_add_93852_comb + p2_add_93139;
  assign p3_add_93951_comb = p3_add_93851_comb + p2_add_93138;
  assign p3_add_93950_comb = p3_add_93850_comb + p2_add_93137;
  assign p3_add_93949_comb = p3_add_93849_comb + p2_add_93136;
  assign p3_add_93948_comb = p3_add_93848_comb + p2_add_93135;
  assign p3_add_93947_comb = p3_add_93847_comb + p2_add_93134;
  assign p3_add_93946_comb = p3_add_93846_comb + p2_add_93133;
  assign p3_add_93945_comb = p3_add_93845_comb + p2_add_93132;
  assign p3_add_93944_comb = p3_add_93844_comb + p2_add_93131;
  assign p3_add_93943_comb = p3_add_93843_comb + p2_add_93130;
  assign p3_add_93942_comb = p3_add_93842_comb + p2_add_93129;
  assign p3_add_93941_comb = p3_add_93841_comb + p2_add_93128;
  assign p3_add_93940_comb = p3_add_93840_comb + p2_add_93127;
  assign p3_add_93939_comb = p3_add_93839_comb + p2_add_93126;
  assign p3_add_93938_comb = p3_add_93838_comb + p2_add_93125;
  assign p3_add_93937_comb = p3_add_93837_comb + p2_add_93124;
  assign p3_add_93936_comb = p3_add_93836_comb + p2_add_93123;
  assign p3_add_93935_comb = p3_add_93835_comb + p2_add_93122;
  assign p3_add_93934_comb = p3_add_93834_comb + p2_add_93121;
  assign p3_add_93933_comb = p3_add_93833_comb + p2_add_93120;
  assign p3_add_93932_comb = p3_add_93832_comb + p2_add_93119;
  assign p3_add_93931_comb = p3_add_93831_comb + p2_add_93118;
  assign p3_add_93930_comb = p3_add_93830_comb + p2_add_93117;
  assign p3_add_93929_comb = p3_add_93829_comb + p2_add_93116;
  assign p3_add_93928_comb = p3_add_93828_comb + p2_add_93115;
  assign p3_add_93927_comb = p3_add_93827_comb + p2_add_93114;
  assign p3_add_93926_comb = p3_add_93826_comb + p2_add_93113;

  // Registers for pipe stage 3:
  reg [31:0] p3_add_94025;
  reg [31:0] p3_add_94024;
  reg [31:0] p3_add_94023;
  reg [31:0] p3_add_94022;
  reg [31:0] p3_add_94021;
  reg [31:0] p3_add_94020;
  reg [31:0] p3_add_94019;
  reg [31:0] p3_add_94018;
  reg [31:0] p3_add_94017;
  reg [31:0] p3_add_94016;
  reg [31:0] p3_add_94015;
  reg [31:0] p3_add_94014;
  reg [31:0] p3_add_94013;
  reg [31:0] p3_add_94012;
  reg [31:0] p3_add_94011;
  reg [31:0] p3_add_94010;
  reg [31:0] p3_add_94009;
  reg [31:0] p3_add_94008;
  reg [31:0] p3_add_94007;
  reg [31:0] p3_add_94006;
  reg [31:0] p3_add_94005;
  reg [31:0] p3_add_94004;
  reg [31:0] p3_add_94003;
  reg [31:0] p3_add_94002;
  reg [31:0] p3_add_94001;
  reg [31:0] p3_add_94000;
  reg [31:0] p3_add_93999;
  reg [31:0] p3_add_93998;
  reg [31:0] p3_add_93997;
  reg [31:0] p3_add_93996;
  reg [31:0] p3_add_93995;
  reg [31:0] p3_add_93994;
  reg [31:0] p3_add_93993;
  reg [31:0] p3_add_93992;
  reg [31:0] p3_add_93991;
  reg [31:0] p3_add_93990;
  reg [31:0] p3_add_93989;
  reg [31:0] p3_add_93988;
  reg [31:0] p3_add_93987;
  reg [31:0] p3_add_93986;
  reg [31:0] p3_add_93985;
  reg [31:0] p3_add_93984;
  reg [31:0] p3_add_93983;
  reg [31:0] p3_add_93982;
  reg [31:0] p3_add_93981;
  reg [31:0] p3_add_93980;
  reg [31:0] p3_add_93979;
  reg [31:0] p3_add_93978;
  reg [31:0] p3_add_93977;
  reg [31:0] p3_add_93976;
  reg [31:0] p3_add_93975;
  reg [31:0] p3_add_93974;
  reg [31:0] p3_add_93973;
  reg [31:0] p3_add_93972;
  reg [31:0] p3_add_93971;
  reg [31:0] p3_add_93970;
  reg [31:0] p3_add_93969;
  reg [31:0] p3_add_93968;
  reg [31:0] p3_add_93967;
  reg [31:0] p3_add_93966;
  reg [31:0] p3_add_93965;
  reg [31:0] p3_add_93964;
  reg [31:0] p3_add_93963;
  reg [31:0] p3_add_93962;
  reg [31:0] p3_add_93961;
  reg [31:0] p3_add_93960;
  reg [31:0] p3_add_93959;
  reg [31:0] p3_add_93958;
  reg [31:0] p3_add_93957;
  reg [31:0] p3_add_93956;
  reg [31:0] p3_add_93955;
  reg [31:0] p3_add_93954;
  reg [31:0] p3_add_93953;
  reg [31:0] p3_add_93952;
  reg [31:0] p3_add_93951;
  reg [31:0] p3_add_93950;
  reg [31:0] p3_add_93949;
  reg [31:0] p3_add_93948;
  reg [31:0] p3_add_93947;
  reg [31:0] p3_add_93946;
  reg [31:0] p3_add_93945;
  reg [31:0] p3_add_93944;
  reg [31:0] p3_add_93943;
  reg [31:0] p3_add_93942;
  reg [31:0] p3_add_93941;
  reg [31:0] p3_add_93940;
  reg [31:0] p3_add_93939;
  reg [31:0] p3_add_93938;
  reg [31:0] p3_add_93937;
  reg [31:0] p3_add_93936;
  reg [31:0] p3_add_93935;
  reg [31:0] p3_add_93934;
  reg [31:0] p3_add_93933;
  reg [31:0] p3_add_93932;
  reg [31:0] p3_add_93931;
  reg [31:0] p3_add_93930;
  reg [31:0] p3_add_93929;
  reg [31:0] p3_add_93928;
  reg [31:0] p3_add_93927;
  reg [31:0] p3_add_93926;
  always_ff @ (posedge clk) begin
    p3_add_94025 <= p3_add_94025_comb;
    p3_add_94024 <= p3_add_94024_comb;
    p3_add_94023 <= p3_add_94023_comb;
    p3_add_94022 <= p3_add_94022_comb;
    p3_add_94021 <= p3_add_94021_comb;
    p3_add_94020 <= p3_add_94020_comb;
    p3_add_94019 <= p3_add_94019_comb;
    p3_add_94018 <= p3_add_94018_comb;
    p3_add_94017 <= p3_add_94017_comb;
    p3_add_94016 <= p3_add_94016_comb;
    p3_add_94015 <= p3_add_94015_comb;
    p3_add_94014 <= p3_add_94014_comb;
    p3_add_94013 <= p3_add_94013_comb;
    p3_add_94012 <= p3_add_94012_comb;
    p3_add_94011 <= p3_add_94011_comb;
    p3_add_94010 <= p3_add_94010_comb;
    p3_add_94009 <= p3_add_94009_comb;
    p3_add_94008 <= p3_add_94008_comb;
    p3_add_94007 <= p3_add_94007_comb;
    p3_add_94006 <= p3_add_94006_comb;
    p3_add_94005 <= p3_add_94005_comb;
    p3_add_94004 <= p3_add_94004_comb;
    p3_add_94003 <= p3_add_94003_comb;
    p3_add_94002 <= p3_add_94002_comb;
    p3_add_94001 <= p3_add_94001_comb;
    p3_add_94000 <= p3_add_94000_comb;
    p3_add_93999 <= p3_add_93999_comb;
    p3_add_93998 <= p3_add_93998_comb;
    p3_add_93997 <= p3_add_93997_comb;
    p3_add_93996 <= p3_add_93996_comb;
    p3_add_93995 <= p3_add_93995_comb;
    p3_add_93994 <= p3_add_93994_comb;
    p3_add_93993 <= p3_add_93993_comb;
    p3_add_93992 <= p3_add_93992_comb;
    p3_add_93991 <= p3_add_93991_comb;
    p3_add_93990 <= p3_add_93990_comb;
    p3_add_93989 <= p3_add_93989_comb;
    p3_add_93988 <= p3_add_93988_comb;
    p3_add_93987 <= p3_add_93987_comb;
    p3_add_93986 <= p3_add_93986_comb;
    p3_add_93985 <= p3_add_93985_comb;
    p3_add_93984 <= p3_add_93984_comb;
    p3_add_93983 <= p3_add_93983_comb;
    p3_add_93982 <= p3_add_93982_comb;
    p3_add_93981 <= p3_add_93981_comb;
    p3_add_93980 <= p3_add_93980_comb;
    p3_add_93979 <= p3_add_93979_comb;
    p3_add_93978 <= p3_add_93978_comb;
    p3_add_93977 <= p3_add_93977_comb;
    p3_add_93976 <= p3_add_93976_comb;
    p3_add_93975 <= p3_add_93975_comb;
    p3_add_93974 <= p3_add_93974_comb;
    p3_add_93973 <= p3_add_93973_comb;
    p3_add_93972 <= p3_add_93972_comb;
    p3_add_93971 <= p3_add_93971_comb;
    p3_add_93970 <= p3_add_93970_comb;
    p3_add_93969 <= p3_add_93969_comb;
    p3_add_93968 <= p3_add_93968_comb;
    p3_add_93967 <= p3_add_93967_comb;
    p3_add_93966 <= p3_add_93966_comb;
    p3_add_93965 <= p3_add_93965_comb;
    p3_add_93964 <= p3_add_93964_comb;
    p3_add_93963 <= p3_add_93963_comb;
    p3_add_93962 <= p3_add_93962_comb;
    p3_add_93961 <= p3_add_93961_comb;
    p3_add_93960 <= p3_add_93960_comb;
    p3_add_93959 <= p3_add_93959_comb;
    p3_add_93958 <= p3_add_93958_comb;
    p3_add_93957 <= p3_add_93957_comb;
    p3_add_93956 <= p3_add_93956_comb;
    p3_add_93955 <= p3_add_93955_comb;
    p3_add_93954 <= p3_add_93954_comb;
    p3_add_93953 <= p3_add_93953_comb;
    p3_add_93952 <= p3_add_93952_comb;
    p3_add_93951 <= p3_add_93951_comb;
    p3_add_93950 <= p3_add_93950_comb;
    p3_add_93949 <= p3_add_93949_comb;
    p3_add_93948 <= p3_add_93948_comb;
    p3_add_93947 <= p3_add_93947_comb;
    p3_add_93946 <= p3_add_93946_comb;
    p3_add_93945 <= p3_add_93945_comb;
    p3_add_93944 <= p3_add_93944_comb;
    p3_add_93943 <= p3_add_93943_comb;
    p3_add_93942 <= p3_add_93942_comb;
    p3_add_93941 <= p3_add_93941_comb;
    p3_add_93940 <= p3_add_93940_comb;
    p3_add_93939 <= p3_add_93939_comb;
    p3_add_93938 <= p3_add_93938_comb;
    p3_add_93937 <= p3_add_93937_comb;
    p3_add_93936 <= p3_add_93936_comb;
    p3_add_93935 <= p3_add_93935_comb;
    p3_add_93934 <= p3_add_93934_comb;
    p3_add_93933 <= p3_add_93933_comb;
    p3_add_93932 <= p3_add_93932_comb;
    p3_add_93931 <= p3_add_93931_comb;
    p3_add_93930 <= p3_add_93930_comb;
    p3_add_93929 <= p3_add_93929_comb;
    p3_add_93928 <= p3_add_93928_comb;
    p3_add_93927 <= p3_add_93927_comb;
    p3_add_93926 <= p3_add_93926_comb;
  end

  // ===== Pipe stage 4:

  // Registers for pipe stage 4:
  reg [31:0] p4_add_94025;
  reg [31:0] p4_add_94024;
  reg [31:0] p4_add_94023;
  reg [31:0] p4_add_94022;
  reg [31:0] p4_add_94021;
  reg [31:0] p4_add_94020;
  reg [31:0] p4_add_94019;
  reg [31:0] p4_add_94018;
  reg [31:0] p4_add_94017;
  reg [31:0] p4_add_94016;
  reg [31:0] p4_add_94015;
  reg [31:0] p4_add_94014;
  reg [31:0] p4_add_94013;
  reg [31:0] p4_add_94012;
  reg [31:0] p4_add_94011;
  reg [31:0] p4_add_94010;
  reg [31:0] p4_add_94009;
  reg [31:0] p4_add_94008;
  reg [31:0] p4_add_94007;
  reg [31:0] p4_add_94006;
  reg [31:0] p4_add_94005;
  reg [31:0] p4_add_94004;
  reg [31:0] p4_add_94003;
  reg [31:0] p4_add_94002;
  reg [31:0] p4_add_94001;
  reg [31:0] p4_add_94000;
  reg [31:0] p4_add_93999;
  reg [31:0] p4_add_93998;
  reg [31:0] p4_add_93997;
  reg [31:0] p4_add_93996;
  reg [31:0] p4_add_93995;
  reg [31:0] p4_add_93994;
  reg [31:0] p4_add_93993;
  reg [31:0] p4_add_93992;
  reg [31:0] p4_add_93991;
  reg [31:0] p4_add_93990;
  reg [31:0] p4_add_93989;
  reg [31:0] p4_add_93988;
  reg [31:0] p4_add_93987;
  reg [31:0] p4_add_93986;
  reg [31:0] p4_add_93985;
  reg [31:0] p4_add_93984;
  reg [31:0] p4_add_93983;
  reg [31:0] p4_add_93982;
  reg [31:0] p4_add_93981;
  reg [31:0] p4_add_93980;
  reg [31:0] p4_add_93979;
  reg [31:0] p4_add_93978;
  reg [31:0] p4_add_93977;
  reg [31:0] p4_add_93976;
  reg [31:0] p4_add_93975;
  reg [31:0] p4_add_93974;
  reg [31:0] p4_add_93973;
  reg [31:0] p4_add_93972;
  reg [31:0] p4_add_93971;
  reg [31:0] p4_add_93970;
  reg [31:0] p4_add_93969;
  reg [31:0] p4_add_93968;
  reg [31:0] p4_add_93967;
  reg [31:0] p4_add_93966;
  reg [31:0] p4_add_93965;
  reg [31:0] p4_add_93964;
  reg [31:0] p4_add_93963;
  reg [31:0] p4_add_93962;
  reg [31:0] p4_add_93961;
  reg [31:0] p4_add_93960;
  reg [31:0] p4_add_93959;
  reg [31:0] p4_add_93958;
  reg [31:0] p4_add_93957;
  reg [31:0] p4_add_93956;
  reg [31:0] p4_add_93955;
  reg [31:0] p4_add_93954;
  reg [31:0] p4_add_93953;
  reg [31:0] p4_add_93952;
  reg [31:0] p4_add_93951;
  reg [31:0] p4_add_93950;
  reg [31:0] p4_add_93949;
  reg [31:0] p4_add_93948;
  reg [31:0] p4_add_93947;
  reg [31:0] p4_add_93946;
  reg [31:0] p4_add_93945;
  reg [31:0] p4_add_93944;
  reg [31:0] p4_add_93943;
  reg [31:0] p4_add_93942;
  reg [31:0] p4_add_93941;
  reg [31:0] p4_add_93940;
  reg [31:0] p4_add_93939;
  reg [31:0] p4_add_93938;
  reg [31:0] p4_add_93937;
  reg [31:0] p4_add_93936;
  reg [31:0] p4_add_93935;
  reg [31:0] p4_add_93934;
  reg [31:0] p4_add_93933;
  reg [31:0] p4_add_93932;
  reg [31:0] p4_add_93931;
  reg [31:0] p4_add_93930;
  reg [31:0] p4_add_93929;
  reg [31:0] p4_add_93928;
  reg [31:0] p4_add_93927;
  reg [31:0] p4_add_93926;
  always_ff @ (posedge clk) begin
    p4_add_94025 <= p3_add_94025;
    p4_add_94024 <= p3_add_94024;
    p4_add_94023 <= p3_add_94023;
    p4_add_94022 <= p3_add_94022;
    p4_add_94021 <= p3_add_94021;
    p4_add_94020 <= p3_add_94020;
    p4_add_94019 <= p3_add_94019;
    p4_add_94018 <= p3_add_94018;
    p4_add_94017 <= p3_add_94017;
    p4_add_94016 <= p3_add_94016;
    p4_add_94015 <= p3_add_94015;
    p4_add_94014 <= p3_add_94014;
    p4_add_94013 <= p3_add_94013;
    p4_add_94012 <= p3_add_94012;
    p4_add_94011 <= p3_add_94011;
    p4_add_94010 <= p3_add_94010;
    p4_add_94009 <= p3_add_94009;
    p4_add_94008 <= p3_add_94008;
    p4_add_94007 <= p3_add_94007;
    p4_add_94006 <= p3_add_94006;
    p4_add_94005 <= p3_add_94005;
    p4_add_94004 <= p3_add_94004;
    p4_add_94003 <= p3_add_94003;
    p4_add_94002 <= p3_add_94002;
    p4_add_94001 <= p3_add_94001;
    p4_add_94000 <= p3_add_94000;
    p4_add_93999 <= p3_add_93999;
    p4_add_93998 <= p3_add_93998;
    p4_add_93997 <= p3_add_93997;
    p4_add_93996 <= p3_add_93996;
    p4_add_93995 <= p3_add_93995;
    p4_add_93994 <= p3_add_93994;
    p4_add_93993 <= p3_add_93993;
    p4_add_93992 <= p3_add_93992;
    p4_add_93991 <= p3_add_93991;
    p4_add_93990 <= p3_add_93990;
    p4_add_93989 <= p3_add_93989;
    p4_add_93988 <= p3_add_93988;
    p4_add_93987 <= p3_add_93987;
    p4_add_93986 <= p3_add_93986;
    p4_add_93985 <= p3_add_93985;
    p4_add_93984 <= p3_add_93984;
    p4_add_93983 <= p3_add_93983;
    p4_add_93982 <= p3_add_93982;
    p4_add_93981 <= p3_add_93981;
    p4_add_93980 <= p3_add_93980;
    p4_add_93979 <= p3_add_93979;
    p4_add_93978 <= p3_add_93978;
    p4_add_93977 <= p3_add_93977;
    p4_add_93976 <= p3_add_93976;
    p4_add_93975 <= p3_add_93975;
    p4_add_93974 <= p3_add_93974;
    p4_add_93973 <= p3_add_93973;
    p4_add_93972 <= p3_add_93972;
    p4_add_93971 <= p3_add_93971;
    p4_add_93970 <= p3_add_93970;
    p4_add_93969 <= p3_add_93969;
    p4_add_93968 <= p3_add_93968;
    p4_add_93967 <= p3_add_93967;
    p4_add_93966 <= p3_add_93966;
    p4_add_93965 <= p3_add_93965;
    p4_add_93964 <= p3_add_93964;
    p4_add_93963 <= p3_add_93963;
    p4_add_93962 <= p3_add_93962;
    p4_add_93961 <= p3_add_93961;
    p4_add_93960 <= p3_add_93960;
    p4_add_93959 <= p3_add_93959;
    p4_add_93958 <= p3_add_93958;
    p4_add_93957 <= p3_add_93957;
    p4_add_93956 <= p3_add_93956;
    p4_add_93955 <= p3_add_93955;
    p4_add_93954 <= p3_add_93954;
    p4_add_93953 <= p3_add_93953;
    p4_add_93952 <= p3_add_93952;
    p4_add_93951 <= p3_add_93951;
    p4_add_93950 <= p3_add_93950;
    p4_add_93949 <= p3_add_93949;
    p4_add_93948 <= p3_add_93948;
    p4_add_93947 <= p3_add_93947;
    p4_add_93946 <= p3_add_93946;
    p4_add_93945 <= p3_add_93945;
    p4_add_93944 <= p3_add_93944;
    p4_add_93943 <= p3_add_93943;
    p4_add_93942 <= p3_add_93942;
    p4_add_93941 <= p3_add_93941;
    p4_add_93940 <= p3_add_93940;
    p4_add_93939 <= p3_add_93939;
    p4_add_93938 <= p3_add_93938;
    p4_add_93937 <= p3_add_93937;
    p4_add_93936 <= p3_add_93936;
    p4_add_93935 <= p3_add_93935;
    p4_add_93934 <= p3_add_93934;
    p4_add_93933 <= p3_add_93933;
    p4_add_93932 <= p3_add_93932;
    p4_add_93931 <= p3_add_93931;
    p4_add_93930 <= p3_add_93930;
    p4_add_93929 <= p3_add_93929;
    p4_add_93928 <= p3_add_93928;
    p4_add_93927 <= p3_add_93927;
    p4_add_93926 <= p3_add_93926;
  end

  // ===== Pipe stage 5:
  wire [3499:0] p5_tuple_94852_comb;
  wire p5_tuple_index_94856_comb;
  wire p5_tuple_index_94859_comb;
  wire p5_tuple_index_94862_comb;
  wire p5_tuple_index_94865_comb;
  wire p5_tuple_index_94868_comb;
  wire p5_tuple_index_94871_comb;
  wire p5_tuple_index_94874_comb;
  wire p5_tuple_index_94877_comb;
  wire p5_tuple_index_94880_comb;
  wire p5_tuple_index_94883_comb;
  wire p5_tuple_index_94886_comb;
  wire p5_tuple_index_94889_comb;
  wire p5_tuple_index_94892_comb;
  wire p5_tuple_index_94895_comb;
  wire p5_tuple_index_94898_comb;
  wire p5_tuple_index_94901_comb;
  wire p5_tuple_index_94904_comb;
  wire p5_tuple_index_94907_comb;
  wire p5_tuple_index_94910_comb;
  wire p5_tuple_index_94913_comb;
  wire p5_tuple_index_94916_comb;
  wire p5_tuple_index_94919_comb;
  wire p5_tuple_index_94922_comb;
  wire p5_tuple_index_94925_comb;
  wire p5_tuple_index_94928_comb;
  wire p5_tuple_index_94931_comb;
  wire p5_tuple_index_94934_comb;
  wire p5_tuple_index_94937_comb;
  wire p5_tuple_index_94940_comb;
  wire p5_tuple_index_94943_comb;
  wire p5_tuple_index_94946_comb;
  wire p5_tuple_index_94949_comb;
  wire p5_tuple_index_94952_comb;
  wire p5_tuple_index_94955_comb;
  wire p5_tuple_index_94958_comb;
  wire p5_tuple_index_94961_comb;
  wire p5_tuple_index_94964_comb;
  wire p5_tuple_index_94967_comb;
  wire p5_tuple_index_94970_comb;
  wire p5_tuple_index_94973_comb;
  wire p5_tuple_index_94976_comb;
  wire p5_tuple_index_94979_comb;
  wire p5_tuple_index_94982_comb;
  wire p5_tuple_index_94985_comb;
  wire p5_tuple_index_94988_comb;
  wire p5_tuple_index_94991_comb;
  wire p5_tuple_index_94994_comb;
  wire p5_tuple_index_94997_comb;
  wire p5_tuple_index_95000_comb;
  wire p5_tuple_index_95003_comb;
  wire p5_tuple_index_95006_comb;
  wire p5_tuple_index_95009_comb;
  wire p5_tuple_index_95012_comb;
  wire p5_tuple_index_95015_comb;
  wire p5_tuple_index_95018_comb;
  wire p5_tuple_index_95021_comb;
  wire p5_tuple_index_95024_comb;
  wire p5_tuple_index_95027_comb;
  wire p5_tuple_index_95030_comb;
  wire p5_tuple_index_95033_comb;
  wire p5_tuple_index_95036_comb;
  wire p5_tuple_index_95039_comb;
  wire p5_tuple_index_95042_comb;
  wire p5_tuple_index_95045_comb;
  wire p5_tuple_index_95048_comb;
  wire p5_tuple_index_95051_comb;
  wire p5_tuple_index_95054_comb;
  wire p5_tuple_index_95057_comb;
  wire p5_tuple_index_95060_comb;
  wire p5_tuple_index_95063_comb;
  wire p5_tuple_index_95066_comb;
  wire p5_tuple_index_95069_comb;
  wire p5_tuple_index_95072_comb;
  wire p5_tuple_index_95075_comb;
  wire p5_tuple_index_95078_comb;
  wire p5_tuple_index_95081_comb;
  wire p5_tuple_index_95084_comb;
  wire p5_tuple_index_95087_comb;
  wire p5_tuple_index_95090_comb;
  wire p5_tuple_index_95093_comb;
  wire p5_tuple_index_95096_comb;
  wire p5_tuple_index_95099_comb;
  wire p5_tuple_index_95102_comb;
  wire p5_tuple_index_95105_comb;
  wire p5_tuple_index_95108_comb;
  wire p5_tuple_index_95111_comb;
  wire p5_tuple_index_95114_comb;
  wire p5_tuple_index_95117_comb;
  wire p5_tuple_index_95120_comb;
  wire p5_tuple_index_95123_comb;
  wire p5_tuple_index_95126_comb;
  wire p5_tuple_index_95129_comb;
  wire p5_tuple_index_95132_comb;
  wire p5_tuple_index_95135_comb;
  wire p5_tuple_index_95138_comb;
  wire p5_tuple_index_95141_comb;
  wire p5_tuple_index_95144_comb;
  wire p5_tuple_index_95147_comb;
  wire p5_tuple_index_95150_comb;
  wire p5_tuple_index_95153_comb;
  wire p5_tuple_index_95156_comb;
  wire p5_tuple_index_95159_comb;
  wire p5_tuple_index_95162_comb;
  wire p5_tuple_index_95165_comb;
  wire p5_tuple_index_95168_comb;
  wire p5_tuple_index_95171_comb;
  wire p5_tuple_index_95174_comb;
  wire p5_tuple_index_95177_comb;
  wire p5_tuple_index_95180_comb;
  wire p5_tuple_index_95183_comb;
  wire p5_tuple_index_95186_comb;
  wire p5_tuple_index_95189_comb;
  wire p5_tuple_index_95192_comb;
  wire p5_tuple_index_95195_comb;
  wire p5_tuple_index_95198_comb;
  wire p5_tuple_index_95201_comb;
  wire p5_tuple_index_95204_comb;
  wire p5_tuple_index_95207_comb;
  wire p5_tuple_index_95210_comb;
  wire p5_tuple_index_95213_comb;
  wire p5_tuple_index_95216_comb;
  wire p5_tuple_index_95219_comb;
  wire p5_tuple_index_95222_comb;
  wire p5_tuple_index_95225_comb;
  wire p5_tuple_index_95228_comb;
  wire p5_tuple_index_95231_comb;
  wire p5_tuple_index_95234_comb;
  wire p5_tuple_index_95237_comb;
  wire p5_tuple_index_95240_comb;
  wire p5_tuple_index_95243_comb;
  wire p5_tuple_index_95246_comb;
  wire p5_tuple_index_95249_comb;
  wire p5_tuple_index_95252_comb;
  wire p5_tuple_index_95255_comb;
  wire p5_tuple_index_95258_comb;
  wire p5_tuple_index_95261_comb;
  wire p5_tuple_index_95264_comb;
  wire p5_tuple_index_95267_comb;
  wire p5_tuple_index_95270_comb;
  wire p5_tuple_index_95273_comb;
  wire p5_tuple_index_95276_comb;
  wire p5_tuple_index_95279_comb;
  wire p5_tuple_index_95282_comb;
  wire p5_tuple_index_95285_comb;
  wire p5_tuple_index_95288_comb;
  wire p5_tuple_index_95291_comb;
  wire p5_tuple_index_95294_comb;
  wire p5_tuple_index_95297_comb;
  wire p5_tuple_index_95300_comb;
  wire p5_tuple_index_95303_comb;
  wire p5_tuple_index_95306_comb;
  wire p5_tuple_index_95309_comb;
  wire p5_tuple_index_95312_comb;
  wire p5_tuple_index_95315_comb;
  wire p5_tuple_index_95318_comb;
  wire p5_tuple_index_95321_comb;
  wire p5_tuple_index_95324_comb;
  wire p5_tuple_index_95327_comb;
  wire p5_tuple_index_95330_comb;
  wire p5_tuple_index_95333_comb;
  wire p5_tuple_index_95336_comb;
  wire p5_tuple_index_95339_comb;
  wire p5_tuple_index_95342_comb;
  wire p5_tuple_index_95345_comb;
  wire p5_tuple_index_95348_comb;
  wire p5_tuple_index_95351_comb;
  wire p5_tuple_index_95354_comb;
  wire p5_tuple_index_95357_comb;
  wire p5_tuple_index_95360_comb;
  wire p5_tuple_index_95363_comb;
  wire p5_tuple_index_95366_comb;
  wire p5_tuple_index_95369_comb;
  wire p5_tuple_index_95372_comb;
  wire p5_tuple_index_95375_comb;
  wire p5_tuple_index_95378_comb;
  wire p5_tuple_index_95381_comb;
  wire p5_tuple_index_95384_comb;
  wire p5_tuple_index_95387_comb;
  wire p5_tuple_index_95390_comb;
  wire p5_tuple_index_95393_comb;
  wire p5_tuple_index_95396_comb;
  wire p5_tuple_index_95399_comb;
  wire p5_tuple_index_95402_comb;
  wire p5_tuple_index_95405_comb;
  wire p5_tuple_index_95408_comb;
  wire p5_tuple_index_95411_comb;
  wire p5_tuple_index_95414_comb;
  wire p5_tuple_index_95417_comb;
  wire p5_tuple_index_95420_comb;
  wire p5_tuple_index_95423_comb;
  wire p5_tuple_index_95426_comb;
  wire p5_tuple_index_95429_comb;
  wire p5_tuple_index_95432_comb;
  wire p5_tuple_index_95435_comb;
  wire p5_tuple_index_95438_comb;
  wire p5_tuple_index_95441_comb;
  wire p5_tuple_index_95444_comb;
  wire p5_tuple_index_95447_comb;
  wire p5_tuple_index_95450_comb;
  wire p5_tuple_index_95453_comb;
  wire [32:0] p5_tuple_index_95456_comb;
  wire [32:0] p5_tuple_index_95459_comb;
  wire [32:0] p5_tuple_index_95462_comb;
  wire [32:0] p5_tuple_index_95465_comb;
  wire [32:0] p5_tuple_index_95468_comb;
  wire [32:0] p5_tuple_index_95471_comb;
  wire [32:0] p5_tuple_index_95474_comb;
  wire [32:0] p5_tuple_index_95477_comb;
  wire [32:0] p5_tuple_index_95480_comb;
  wire [32:0] p5_tuple_index_95483_comb;
  wire [32:0] p5_tuple_index_95486_comb;
  wire [32:0] p5_tuple_index_95489_comb;
  wire [32:0] p5_tuple_index_95492_comb;
  wire [32:0] p5_tuple_index_95495_comb;
  wire [32:0] p5_tuple_index_95498_comb;
  wire [32:0] p5_tuple_index_95501_comb;
  wire [32:0] p5_tuple_index_95504_comb;
  wire [32:0] p5_tuple_index_95507_comb;
  wire [32:0] p5_tuple_index_95510_comb;
  wire [32:0] p5_tuple_index_95513_comb;
  wire [32:0] p5_tuple_index_95516_comb;
  wire [32:0] p5_tuple_index_95519_comb;
  wire [32:0] p5_tuple_index_95522_comb;
  wire [32:0] p5_tuple_index_95525_comb;
  wire [32:0] p5_tuple_index_95528_comb;
  wire [32:0] p5_tuple_index_95531_comb;
  wire [32:0] p5_tuple_index_95534_comb;
  wire [32:0] p5_tuple_index_95537_comb;
  wire [32:0] p5_tuple_index_95540_comb;
  wire [32:0] p5_tuple_index_95543_comb;
  wire [32:0] p5_tuple_index_95546_comb;
  wire [32:0] p5_tuple_index_95549_comb;
  wire [32:0] p5_tuple_index_95552_comb;
  wire [32:0] p5_tuple_index_95555_comb;
  wire [32:0] p5_tuple_index_95558_comb;
  wire [32:0] p5_tuple_index_95561_comb;
  wire [32:0] p5_tuple_index_95564_comb;
  wire [32:0] p5_tuple_index_95567_comb;
  wire [32:0] p5_tuple_index_95570_comb;
  wire [32:0] p5_tuple_index_95573_comb;
  wire [32:0] p5_tuple_index_95576_comb;
  wire [32:0] p5_tuple_index_95579_comb;
  wire [32:0] p5_tuple_index_95582_comb;
  wire [32:0] p5_tuple_index_95585_comb;
  wire [32:0] p5_tuple_index_95588_comb;
  wire [32:0] p5_tuple_index_95591_comb;
  wire [32:0] p5_tuple_index_95594_comb;
  wire [32:0] p5_tuple_index_95597_comb;
  wire [32:0] p5_tuple_index_95600_comb;
  wire [32:0] p5_tuple_index_95603_comb;
  wire [32:0] p5_tuple_index_95606_comb;
  wire [32:0] p5_tuple_index_95609_comb;
  wire [32:0] p5_tuple_index_95612_comb;
  wire [32:0] p5_tuple_index_95615_comb;
  wire [32:0] p5_tuple_index_95618_comb;
  wire [32:0] p5_tuple_index_95621_comb;
  wire [32:0] p5_tuple_index_95624_comb;
  wire [32:0] p5_tuple_index_95627_comb;
  wire [32:0] p5_tuple_index_95630_comb;
  wire [32:0] p5_tuple_index_95633_comb;
  wire [32:0] p5_tuple_index_95636_comb;
  wire [32:0] p5_tuple_index_95639_comb;
  wire [32:0] p5_tuple_index_95642_comb;
  wire [32:0] p5_tuple_index_95645_comb;
  wire [32:0] p5_tuple_index_95648_comb;
  wire [32:0] p5_tuple_index_95651_comb;
  wire [32:0] p5_tuple_index_95654_comb;
  wire [32:0] p5_tuple_index_95657_comb;
  wire [32:0] p5_tuple_index_95660_comb;
  wire [32:0] p5_tuple_index_95663_comb;
  wire [32:0] p5_tuple_index_95666_comb;
  wire [32:0] p5_tuple_index_95669_comb;
  wire [32:0] p5_tuple_index_95672_comb;
  wire [32:0] p5_tuple_index_95675_comb;
  wire [32:0] p5_tuple_index_95678_comb;
  wire [32:0] p5_tuple_index_95681_comb;
  wire [32:0] p5_tuple_index_95684_comb;
  wire [32:0] p5_tuple_index_95687_comb;
  wire [32:0] p5_tuple_index_95690_comb;
  wire [32:0] p5_tuple_index_95693_comb;
  wire [32:0] p5_tuple_index_95696_comb;
  wire [32:0] p5_tuple_index_95699_comb;
  wire [32:0] p5_tuple_index_95702_comb;
  wire [32:0] p5_tuple_index_95705_comb;
  wire [32:0] p5_tuple_index_95708_comb;
  wire [32:0] p5_tuple_index_95711_comb;
  wire [32:0] p5_tuple_index_95714_comb;
  wire [32:0] p5_tuple_index_95717_comb;
  wire [32:0] p5_tuple_index_95720_comb;
  wire [32:0] p5_tuple_index_95723_comb;
  wire [32:0] p5_tuple_index_95726_comb;
  wire [32:0] p5_tuple_index_95729_comb;
  wire [32:0] p5_tuple_index_95732_comb;
  wire [32:0] p5_tuple_index_95735_comb;
  wire [32:0] p5_tuple_index_95738_comb;
  wire [32:0] p5_tuple_index_95741_comb;
  wire [32:0] p5_tuple_index_95744_comb;
  wire [32:0] p5_tuple_index_95747_comb;
  wire [32:0] p5_tuple_index_95750_comb;
  wire [32:0] p5_tuple_index_95753_comb;
  assign p5_tuple_94852_comb = {1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, {p4_add_93926, 1'h1}, {p4_add_93927, 1'h1}, {p4_add_93928, 1'h1}, {p4_add_93929, 1'h1}, {p4_add_93930, 1'h1}, {p4_add_93931, 1'h1}, {p4_add_93932, 1'h1}, {p4_add_93933, 1'h1}, {p4_add_93934, 1'h1}, {p4_add_93935, 1'h1}, {p4_add_93936, 1'h1}, {p4_add_93937, 1'h1}, {p4_add_93938, 1'h1}, {p4_add_93939, 1'h1}, {p4_add_93940, 1'h1}, {p4_add_93941, 1'h1}, {p4_add_93942, 1'h1}, {p4_add_93943, 1'h1}, {p4_add_93944, 1'h1}, {p4_add_93945, 1'h1}, {p4_add_93946, 1'h1}, {p4_add_93947, 1'h1}, {p4_add_93948, 1'h1}, {p4_add_93949, 1'h1}, {p4_add_93950, 1'h1}, {p4_add_93951, 1'h1}, {p4_add_93952, 1'h1}, {p4_add_93953, 1'h1}, {p4_add_93954, 1'h1}, {p4_add_93955, 1'h1}, {p4_add_93956, 1'h1}, {p4_add_93957, 1'h1}, {p4_add_93958, 1'h1}, {p4_add_93959, 1'h1}, {p4_add_93960, 1'h1}, {p4_add_93961, 1'h1}, {p4_add_93962, 1'h1}, {p4_add_93963, 1'h1}, {p4_add_93964, 1'h1}, {p4_add_93965, 1'h1}, {p4_add_93966, 1'h1}, {p4_add_93967, 1'h1}, {p4_add_93968, 1'h1}, {p4_add_93969, 1'h1}, {p4_add_93970, 1'h1}, {p4_add_93971, 1'h1}, {p4_add_93972, 1'h1}, {p4_add_93973, 1'h1}, {p4_add_93974, 1'h1}, {p4_add_93975, 1'h1}, {p4_add_93976, 1'h1}, {p4_add_93977, 1'h1}, {p4_add_93978, 1'h1}, {p4_add_93979, 1'h1}, {p4_add_93980, 1'h1}, {p4_add_93981, 1'h1}, {p4_add_93982, 1'h1}, {p4_add_93983, 1'h1}, {p4_add_93984, 1'h1}, {p4_add_93985, 1'h1}, {p4_add_93986, 1'h1}, {p4_add_93987, 1'h1}, {p4_add_93988, 1'h1}, {p4_add_93989, 1'h1}, {p4_add_93990, 1'h1}, {p4_add_93991, 1'h1}, {p4_add_93992, 1'h1}, {p4_add_93993, 1'h1}, {p4_add_93994, 1'h1}, {p4_add_93995, 1'h1}, {p4_add_93996, 1'h1}, {p4_add_93997, 1'h1}, {p4_add_93998, 1'h1}, {p4_add_93999, 1'h1}, {p4_add_94000, 1'h1}, {p4_add_94001, 1'h1}, {p4_add_94002, 1'h1}, {p4_add_94003, 1'h1}, {p4_add_94004, 1'h1}, {p4_add_94005, 1'h1}, {p4_add_94006, 1'h1}, {p4_add_94007, 1'h1}, {p4_add_94008, 1'h1}, {p4_add_94009, 1'h1}, {p4_add_94010, 1'h1}, {p4_add_94011, 1'h1}, {p4_add_94012, 1'h1}, {p4_add_94013, 1'h1}, {p4_add_94014, 1'h1}, {p4_add_94015, 1'h1}, {p4_add_94016, 1'h1}, {p4_add_94017, 1'h1}, {p4_add_94018, 1'h1}, {p4_add_94019, 1'h1}, {p4_add_94020, 1'h1}, {p4_add_94021, 1'h1}, {p4_add_94022, 1'h1}, {p4_add_94023, 1'h1}, {p4_add_94024, 1'h1}, {p4_add_94025, 1'h1}};
  assign p5_tuple_index_94856_comb = p5_tuple_94852_comb[3499:3499];
  assign p5_tuple_index_94859_comb = p5_tuple_94852_comb[3498:3498];
  assign p5_tuple_index_94862_comb = p5_tuple_94852_comb[3497:3497];
  assign p5_tuple_index_94865_comb = p5_tuple_94852_comb[3496:3496];
  assign p5_tuple_index_94868_comb = p5_tuple_94852_comb[3495:3495];
  assign p5_tuple_index_94871_comb = p5_tuple_94852_comb[3494:3494];
  assign p5_tuple_index_94874_comb = p5_tuple_94852_comb[3493:3493];
  assign p5_tuple_index_94877_comb = p5_tuple_94852_comb[3492:3492];
  assign p5_tuple_index_94880_comb = p5_tuple_94852_comb[3491:3491];
  assign p5_tuple_index_94883_comb = p5_tuple_94852_comb[3490:3490];
  assign p5_tuple_index_94886_comb = p5_tuple_94852_comb[3489:3489];
  assign p5_tuple_index_94889_comb = p5_tuple_94852_comb[3488:3488];
  assign p5_tuple_index_94892_comb = p5_tuple_94852_comb[3487:3487];
  assign p5_tuple_index_94895_comb = p5_tuple_94852_comb[3486:3486];
  assign p5_tuple_index_94898_comb = p5_tuple_94852_comb[3485:3485];
  assign p5_tuple_index_94901_comb = p5_tuple_94852_comb[3484:3484];
  assign p5_tuple_index_94904_comb = p5_tuple_94852_comb[3483:3483];
  assign p5_tuple_index_94907_comb = p5_tuple_94852_comb[3482:3482];
  assign p5_tuple_index_94910_comb = p5_tuple_94852_comb[3481:3481];
  assign p5_tuple_index_94913_comb = p5_tuple_94852_comb[3480:3480];
  assign p5_tuple_index_94916_comb = p5_tuple_94852_comb[3479:3479];
  assign p5_tuple_index_94919_comb = p5_tuple_94852_comb[3478:3478];
  assign p5_tuple_index_94922_comb = p5_tuple_94852_comb[3477:3477];
  assign p5_tuple_index_94925_comb = p5_tuple_94852_comb[3476:3476];
  assign p5_tuple_index_94928_comb = p5_tuple_94852_comb[3475:3475];
  assign p5_tuple_index_94931_comb = p5_tuple_94852_comb[3474:3474];
  assign p5_tuple_index_94934_comb = p5_tuple_94852_comb[3473:3473];
  assign p5_tuple_index_94937_comb = p5_tuple_94852_comb[3472:3472];
  assign p5_tuple_index_94940_comb = p5_tuple_94852_comb[3471:3471];
  assign p5_tuple_index_94943_comb = p5_tuple_94852_comb[3470:3470];
  assign p5_tuple_index_94946_comb = p5_tuple_94852_comb[3469:3469];
  assign p5_tuple_index_94949_comb = p5_tuple_94852_comb[3468:3468];
  assign p5_tuple_index_94952_comb = p5_tuple_94852_comb[3467:3467];
  assign p5_tuple_index_94955_comb = p5_tuple_94852_comb[3466:3466];
  assign p5_tuple_index_94958_comb = p5_tuple_94852_comb[3465:3465];
  assign p5_tuple_index_94961_comb = p5_tuple_94852_comb[3464:3464];
  assign p5_tuple_index_94964_comb = p5_tuple_94852_comb[3463:3463];
  assign p5_tuple_index_94967_comb = p5_tuple_94852_comb[3462:3462];
  assign p5_tuple_index_94970_comb = p5_tuple_94852_comb[3461:3461];
  assign p5_tuple_index_94973_comb = p5_tuple_94852_comb[3460:3460];
  assign p5_tuple_index_94976_comb = p5_tuple_94852_comb[3459:3459];
  assign p5_tuple_index_94979_comb = p5_tuple_94852_comb[3458:3458];
  assign p5_tuple_index_94982_comb = p5_tuple_94852_comb[3457:3457];
  assign p5_tuple_index_94985_comb = p5_tuple_94852_comb[3456:3456];
  assign p5_tuple_index_94988_comb = p5_tuple_94852_comb[3455:3455];
  assign p5_tuple_index_94991_comb = p5_tuple_94852_comb[3454:3454];
  assign p5_tuple_index_94994_comb = p5_tuple_94852_comb[3453:3453];
  assign p5_tuple_index_94997_comb = p5_tuple_94852_comb[3452:3452];
  assign p5_tuple_index_95000_comb = p5_tuple_94852_comb[3451:3451];
  assign p5_tuple_index_95003_comb = p5_tuple_94852_comb[3450:3450];
  assign p5_tuple_index_95006_comb = p5_tuple_94852_comb[3449:3449];
  assign p5_tuple_index_95009_comb = p5_tuple_94852_comb[3448:3448];
  assign p5_tuple_index_95012_comb = p5_tuple_94852_comb[3447:3447];
  assign p5_tuple_index_95015_comb = p5_tuple_94852_comb[3446:3446];
  assign p5_tuple_index_95018_comb = p5_tuple_94852_comb[3445:3445];
  assign p5_tuple_index_95021_comb = p5_tuple_94852_comb[3444:3444];
  assign p5_tuple_index_95024_comb = p5_tuple_94852_comb[3443:3443];
  assign p5_tuple_index_95027_comb = p5_tuple_94852_comb[3442:3442];
  assign p5_tuple_index_95030_comb = p5_tuple_94852_comb[3441:3441];
  assign p5_tuple_index_95033_comb = p5_tuple_94852_comb[3440:3440];
  assign p5_tuple_index_95036_comb = p5_tuple_94852_comb[3439:3439];
  assign p5_tuple_index_95039_comb = p5_tuple_94852_comb[3438:3438];
  assign p5_tuple_index_95042_comb = p5_tuple_94852_comb[3437:3437];
  assign p5_tuple_index_95045_comb = p5_tuple_94852_comb[3436:3436];
  assign p5_tuple_index_95048_comb = p5_tuple_94852_comb[3435:3435];
  assign p5_tuple_index_95051_comb = p5_tuple_94852_comb[3434:3434];
  assign p5_tuple_index_95054_comb = p5_tuple_94852_comb[3433:3433];
  assign p5_tuple_index_95057_comb = p5_tuple_94852_comb[3432:3432];
  assign p5_tuple_index_95060_comb = p5_tuple_94852_comb[3431:3431];
  assign p5_tuple_index_95063_comb = p5_tuple_94852_comb[3430:3430];
  assign p5_tuple_index_95066_comb = p5_tuple_94852_comb[3429:3429];
  assign p5_tuple_index_95069_comb = p5_tuple_94852_comb[3428:3428];
  assign p5_tuple_index_95072_comb = p5_tuple_94852_comb[3427:3427];
  assign p5_tuple_index_95075_comb = p5_tuple_94852_comb[3426:3426];
  assign p5_tuple_index_95078_comb = p5_tuple_94852_comb[3425:3425];
  assign p5_tuple_index_95081_comb = p5_tuple_94852_comb[3424:3424];
  assign p5_tuple_index_95084_comb = p5_tuple_94852_comb[3423:3423];
  assign p5_tuple_index_95087_comb = p5_tuple_94852_comb[3422:3422];
  assign p5_tuple_index_95090_comb = p5_tuple_94852_comb[3421:3421];
  assign p5_tuple_index_95093_comb = p5_tuple_94852_comb[3420:3420];
  assign p5_tuple_index_95096_comb = p5_tuple_94852_comb[3419:3419];
  assign p5_tuple_index_95099_comb = p5_tuple_94852_comb[3418:3418];
  assign p5_tuple_index_95102_comb = p5_tuple_94852_comb[3417:3417];
  assign p5_tuple_index_95105_comb = p5_tuple_94852_comb[3416:3416];
  assign p5_tuple_index_95108_comb = p5_tuple_94852_comb[3415:3415];
  assign p5_tuple_index_95111_comb = p5_tuple_94852_comb[3414:3414];
  assign p5_tuple_index_95114_comb = p5_tuple_94852_comb[3413:3413];
  assign p5_tuple_index_95117_comb = p5_tuple_94852_comb[3412:3412];
  assign p5_tuple_index_95120_comb = p5_tuple_94852_comb[3411:3411];
  assign p5_tuple_index_95123_comb = p5_tuple_94852_comb[3410:3410];
  assign p5_tuple_index_95126_comb = p5_tuple_94852_comb[3409:3409];
  assign p5_tuple_index_95129_comb = p5_tuple_94852_comb[3408:3408];
  assign p5_tuple_index_95132_comb = p5_tuple_94852_comb[3407:3407];
  assign p5_tuple_index_95135_comb = p5_tuple_94852_comb[3406:3406];
  assign p5_tuple_index_95138_comb = p5_tuple_94852_comb[3405:3405];
  assign p5_tuple_index_95141_comb = p5_tuple_94852_comb[3404:3404];
  assign p5_tuple_index_95144_comb = p5_tuple_94852_comb[3403:3403];
  assign p5_tuple_index_95147_comb = p5_tuple_94852_comb[3402:3402];
  assign p5_tuple_index_95150_comb = p5_tuple_94852_comb[3401:3401];
  assign p5_tuple_index_95153_comb = p5_tuple_94852_comb[3400:3400];
  assign p5_tuple_index_95156_comb = p5_tuple_94852_comb[3399:3399];
  assign p5_tuple_index_95159_comb = p5_tuple_94852_comb[3398:3398];
  assign p5_tuple_index_95162_comb = p5_tuple_94852_comb[3397:3397];
  assign p5_tuple_index_95165_comb = p5_tuple_94852_comb[3396:3396];
  assign p5_tuple_index_95168_comb = p5_tuple_94852_comb[3395:3395];
  assign p5_tuple_index_95171_comb = p5_tuple_94852_comb[3394:3394];
  assign p5_tuple_index_95174_comb = p5_tuple_94852_comb[3393:3393];
  assign p5_tuple_index_95177_comb = p5_tuple_94852_comb[3392:3392];
  assign p5_tuple_index_95180_comb = p5_tuple_94852_comb[3391:3391];
  assign p5_tuple_index_95183_comb = p5_tuple_94852_comb[3390:3390];
  assign p5_tuple_index_95186_comb = p5_tuple_94852_comb[3389:3389];
  assign p5_tuple_index_95189_comb = p5_tuple_94852_comb[3388:3388];
  assign p5_tuple_index_95192_comb = p5_tuple_94852_comb[3387:3387];
  assign p5_tuple_index_95195_comb = p5_tuple_94852_comb[3386:3386];
  assign p5_tuple_index_95198_comb = p5_tuple_94852_comb[3385:3385];
  assign p5_tuple_index_95201_comb = p5_tuple_94852_comb[3384:3384];
  assign p5_tuple_index_95204_comb = p5_tuple_94852_comb[3383:3383];
  assign p5_tuple_index_95207_comb = p5_tuple_94852_comb[3382:3382];
  assign p5_tuple_index_95210_comb = p5_tuple_94852_comb[3381:3381];
  assign p5_tuple_index_95213_comb = p5_tuple_94852_comb[3380:3380];
  assign p5_tuple_index_95216_comb = p5_tuple_94852_comb[3379:3379];
  assign p5_tuple_index_95219_comb = p5_tuple_94852_comb[3378:3378];
  assign p5_tuple_index_95222_comb = p5_tuple_94852_comb[3377:3377];
  assign p5_tuple_index_95225_comb = p5_tuple_94852_comb[3376:3376];
  assign p5_tuple_index_95228_comb = p5_tuple_94852_comb[3375:3375];
  assign p5_tuple_index_95231_comb = p5_tuple_94852_comb[3374:3374];
  assign p5_tuple_index_95234_comb = p5_tuple_94852_comb[3373:3373];
  assign p5_tuple_index_95237_comb = p5_tuple_94852_comb[3372:3372];
  assign p5_tuple_index_95240_comb = p5_tuple_94852_comb[3371:3371];
  assign p5_tuple_index_95243_comb = p5_tuple_94852_comb[3370:3370];
  assign p5_tuple_index_95246_comb = p5_tuple_94852_comb[3369:3369];
  assign p5_tuple_index_95249_comb = p5_tuple_94852_comb[3368:3368];
  assign p5_tuple_index_95252_comb = p5_tuple_94852_comb[3367:3367];
  assign p5_tuple_index_95255_comb = p5_tuple_94852_comb[3366:3366];
  assign p5_tuple_index_95258_comb = p5_tuple_94852_comb[3365:3365];
  assign p5_tuple_index_95261_comb = p5_tuple_94852_comb[3364:3364];
  assign p5_tuple_index_95264_comb = p5_tuple_94852_comb[3363:3363];
  assign p5_tuple_index_95267_comb = p5_tuple_94852_comb[3362:3362];
  assign p5_tuple_index_95270_comb = p5_tuple_94852_comb[3361:3361];
  assign p5_tuple_index_95273_comb = p5_tuple_94852_comb[3360:3360];
  assign p5_tuple_index_95276_comb = p5_tuple_94852_comb[3359:3359];
  assign p5_tuple_index_95279_comb = p5_tuple_94852_comb[3358:3358];
  assign p5_tuple_index_95282_comb = p5_tuple_94852_comb[3357:3357];
  assign p5_tuple_index_95285_comb = p5_tuple_94852_comb[3356:3356];
  assign p5_tuple_index_95288_comb = p5_tuple_94852_comb[3355:3355];
  assign p5_tuple_index_95291_comb = p5_tuple_94852_comb[3354:3354];
  assign p5_tuple_index_95294_comb = p5_tuple_94852_comb[3353:3353];
  assign p5_tuple_index_95297_comb = p5_tuple_94852_comb[3352:3352];
  assign p5_tuple_index_95300_comb = p5_tuple_94852_comb[3351:3351];
  assign p5_tuple_index_95303_comb = p5_tuple_94852_comb[3350:3350];
  assign p5_tuple_index_95306_comb = p5_tuple_94852_comb[3349:3349];
  assign p5_tuple_index_95309_comb = p5_tuple_94852_comb[3348:3348];
  assign p5_tuple_index_95312_comb = p5_tuple_94852_comb[3347:3347];
  assign p5_tuple_index_95315_comb = p5_tuple_94852_comb[3346:3346];
  assign p5_tuple_index_95318_comb = p5_tuple_94852_comb[3345:3345];
  assign p5_tuple_index_95321_comb = p5_tuple_94852_comb[3344:3344];
  assign p5_tuple_index_95324_comb = p5_tuple_94852_comb[3343:3343];
  assign p5_tuple_index_95327_comb = p5_tuple_94852_comb[3342:3342];
  assign p5_tuple_index_95330_comb = p5_tuple_94852_comb[3341:3341];
  assign p5_tuple_index_95333_comb = p5_tuple_94852_comb[3340:3340];
  assign p5_tuple_index_95336_comb = p5_tuple_94852_comb[3339:3339];
  assign p5_tuple_index_95339_comb = p5_tuple_94852_comb[3338:3338];
  assign p5_tuple_index_95342_comb = p5_tuple_94852_comb[3337:3337];
  assign p5_tuple_index_95345_comb = p5_tuple_94852_comb[3336:3336];
  assign p5_tuple_index_95348_comb = p5_tuple_94852_comb[3335:3335];
  assign p5_tuple_index_95351_comb = p5_tuple_94852_comb[3334:3334];
  assign p5_tuple_index_95354_comb = p5_tuple_94852_comb[3333:3333];
  assign p5_tuple_index_95357_comb = p5_tuple_94852_comb[3332:3332];
  assign p5_tuple_index_95360_comb = p5_tuple_94852_comb[3331:3331];
  assign p5_tuple_index_95363_comb = p5_tuple_94852_comb[3330:3330];
  assign p5_tuple_index_95366_comb = p5_tuple_94852_comb[3329:3329];
  assign p5_tuple_index_95369_comb = p5_tuple_94852_comb[3328:3328];
  assign p5_tuple_index_95372_comb = p5_tuple_94852_comb[3327:3327];
  assign p5_tuple_index_95375_comb = p5_tuple_94852_comb[3326:3326];
  assign p5_tuple_index_95378_comb = p5_tuple_94852_comb[3325:3325];
  assign p5_tuple_index_95381_comb = p5_tuple_94852_comb[3324:3324];
  assign p5_tuple_index_95384_comb = p5_tuple_94852_comb[3323:3323];
  assign p5_tuple_index_95387_comb = p5_tuple_94852_comb[3322:3322];
  assign p5_tuple_index_95390_comb = p5_tuple_94852_comb[3321:3321];
  assign p5_tuple_index_95393_comb = p5_tuple_94852_comb[3320:3320];
  assign p5_tuple_index_95396_comb = p5_tuple_94852_comb[3319:3319];
  assign p5_tuple_index_95399_comb = p5_tuple_94852_comb[3318:3318];
  assign p5_tuple_index_95402_comb = p5_tuple_94852_comb[3317:3317];
  assign p5_tuple_index_95405_comb = p5_tuple_94852_comb[3316:3316];
  assign p5_tuple_index_95408_comb = p5_tuple_94852_comb[3315:3315];
  assign p5_tuple_index_95411_comb = p5_tuple_94852_comb[3314:3314];
  assign p5_tuple_index_95414_comb = p5_tuple_94852_comb[3313:3313];
  assign p5_tuple_index_95417_comb = p5_tuple_94852_comb[3312:3312];
  assign p5_tuple_index_95420_comb = p5_tuple_94852_comb[3311:3311];
  assign p5_tuple_index_95423_comb = p5_tuple_94852_comb[3310:3310];
  assign p5_tuple_index_95426_comb = p5_tuple_94852_comb[3309:3309];
  assign p5_tuple_index_95429_comb = p5_tuple_94852_comb[3308:3308];
  assign p5_tuple_index_95432_comb = p5_tuple_94852_comb[3307:3307];
  assign p5_tuple_index_95435_comb = p5_tuple_94852_comb[3306:3306];
  assign p5_tuple_index_95438_comb = p5_tuple_94852_comb[3305:3305];
  assign p5_tuple_index_95441_comb = p5_tuple_94852_comb[3304:3304];
  assign p5_tuple_index_95444_comb = p5_tuple_94852_comb[3303:3303];
  assign p5_tuple_index_95447_comb = p5_tuple_94852_comb[3302:3302];
  assign p5_tuple_index_95450_comb = p5_tuple_94852_comb[3301:3301];
  assign p5_tuple_index_95453_comb = p5_tuple_94852_comb[3300:3300];
  assign p5_tuple_index_95456_comb = p5_tuple_94852_comb[3299:3267];
  assign p5_tuple_index_95459_comb = p5_tuple_94852_comb[3266:3234];
  assign p5_tuple_index_95462_comb = p5_tuple_94852_comb[3233:3201];
  assign p5_tuple_index_95465_comb = p5_tuple_94852_comb[3200:3168];
  assign p5_tuple_index_95468_comb = p5_tuple_94852_comb[3167:3135];
  assign p5_tuple_index_95471_comb = p5_tuple_94852_comb[3134:3102];
  assign p5_tuple_index_95474_comb = p5_tuple_94852_comb[3101:3069];
  assign p5_tuple_index_95477_comb = p5_tuple_94852_comb[3068:3036];
  assign p5_tuple_index_95480_comb = p5_tuple_94852_comb[3035:3003];
  assign p5_tuple_index_95483_comb = p5_tuple_94852_comb[3002:2970];
  assign p5_tuple_index_95486_comb = p5_tuple_94852_comb[2969:2937];
  assign p5_tuple_index_95489_comb = p5_tuple_94852_comb[2936:2904];
  assign p5_tuple_index_95492_comb = p5_tuple_94852_comb[2903:2871];
  assign p5_tuple_index_95495_comb = p5_tuple_94852_comb[2870:2838];
  assign p5_tuple_index_95498_comb = p5_tuple_94852_comb[2837:2805];
  assign p5_tuple_index_95501_comb = p5_tuple_94852_comb[2804:2772];
  assign p5_tuple_index_95504_comb = p5_tuple_94852_comb[2771:2739];
  assign p5_tuple_index_95507_comb = p5_tuple_94852_comb[2738:2706];
  assign p5_tuple_index_95510_comb = p5_tuple_94852_comb[2705:2673];
  assign p5_tuple_index_95513_comb = p5_tuple_94852_comb[2672:2640];
  assign p5_tuple_index_95516_comb = p5_tuple_94852_comb[2639:2607];
  assign p5_tuple_index_95519_comb = p5_tuple_94852_comb[2606:2574];
  assign p5_tuple_index_95522_comb = p5_tuple_94852_comb[2573:2541];
  assign p5_tuple_index_95525_comb = p5_tuple_94852_comb[2540:2508];
  assign p5_tuple_index_95528_comb = p5_tuple_94852_comb[2507:2475];
  assign p5_tuple_index_95531_comb = p5_tuple_94852_comb[2474:2442];
  assign p5_tuple_index_95534_comb = p5_tuple_94852_comb[2441:2409];
  assign p5_tuple_index_95537_comb = p5_tuple_94852_comb[2408:2376];
  assign p5_tuple_index_95540_comb = p5_tuple_94852_comb[2375:2343];
  assign p5_tuple_index_95543_comb = p5_tuple_94852_comb[2342:2310];
  assign p5_tuple_index_95546_comb = p5_tuple_94852_comb[2309:2277];
  assign p5_tuple_index_95549_comb = p5_tuple_94852_comb[2276:2244];
  assign p5_tuple_index_95552_comb = p5_tuple_94852_comb[2243:2211];
  assign p5_tuple_index_95555_comb = p5_tuple_94852_comb[2210:2178];
  assign p5_tuple_index_95558_comb = p5_tuple_94852_comb[2177:2145];
  assign p5_tuple_index_95561_comb = p5_tuple_94852_comb[2144:2112];
  assign p5_tuple_index_95564_comb = p5_tuple_94852_comb[2111:2079];
  assign p5_tuple_index_95567_comb = p5_tuple_94852_comb[2078:2046];
  assign p5_tuple_index_95570_comb = p5_tuple_94852_comb[2045:2013];
  assign p5_tuple_index_95573_comb = p5_tuple_94852_comb[2012:1980];
  assign p5_tuple_index_95576_comb = p5_tuple_94852_comb[1979:1947];
  assign p5_tuple_index_95579_comb = p5_tuple_94852_comb[1946:1914];
  assign p5_tuple_index_95582_comb = p5_tuple_94852_comb[1913:1881];
  assign p5_tuple_index_95585_comb = p5_tuple_94852_comb[1880:1848];
  assign p5_tuple_index_95588_comb = p5_tuple_94852_comb[1847:1815];
  assign p5_tuple_index_95591_comb = p5_tuple_94852_comb[1814:1782];
  assign p5_tuple_index_95594_comb = p5_tuple_94852_comb[1781:1749];
  assign p5_tuple_index_95597_comb = p5_tuple_94852_comb[1748:1716];
  assign p5_tuple_index_95600_comb = p5_tuple_94852_comb[1715:1683];
  assign p5_tuple_index_95603_comb = p5_tuple_94852_comb[1682:1650];
  assign p5_tuple_index_95606_comb = p5_tuple_94852_comb[1649:1617];
  assign p5_tuple_index_95609_comb = p5_tuple_94852_comb[1616:1584];
  assign p5_tuple_index_95612_comb = p5_tuple_94852_comb[1583:1551];
  assign p5_tuple_index_95615_comb = p5_tuple_94852_comb[1550:1518];
  assign p5_tuple_index_95618_comb = p5_tuple_94852_comb[1517:1485];
  assign p5_tuple_index_95621_comb = p5_tuple_94852_comb[1484:1452];
  assign p5_tuple_index_95624_comb = p5_tuple_94852_comb[1451:1419];
  assign p5_tuple_index_95627_comb = p5_tuple_94852_comb[1418:1386];
  assign p5_tuple_index_95630_comb = p5_tuple_94852_comb[1385:1353];
  assign p5_tuple_index_95633_comb = p5_tuple_94852_comb[1352:1320];
  assign p5_tuple_index_95636_comb = p5_tuple_94852_comb[1319:1287];
  assign p5_tuple_index_95639_comb = p5_tuple_94852_comb[1286:1254];
  assign p5_tuple_index_95642_comb = p5_tuple_94852_comb[1253:1221];
  assign p5_tuple_index_95645_comb = p5_tuple_94852_comb[1220:1188];
  assign p5_tuple_index_95648_comb = p5_tuple_94852_comb[1187:1155];
  assign p5_tuple_index_95651_comb = p5_tuple_94852_comb[1154:1122];
  assign p5_tuple_index_95654_comb = p5_tuple_94852_comb[1121:1089];
  assign p5_tuple_index_95657_comb = p5_tuple_94852_comb[1088:1056];
  assign p5_tuple_index_95660_comb = p5_tuple_94852_comb[1055:1023];
  assign p5_tuple_index_95663_comb = p5_tuple_94852_comb[1022:990];
  assign p5_tuple_index_95666_comb = p5_tuple_94852_comb[989:957];
  assign p5_tuple_index_95669_comb = p5_tuple_94852_comb[956:924];
  assign p5_tuple_index_95672_comb = p5_tuple_94852_comb[923:891];
  assign p5_tuple_index_95675_comb = p5_tuple_94852_comb[890:858];
  assign p5_tuple_index_95678_comb = p5_tuple_94852_comb[857:825];
  assign p5_tuple_index_95681_comb = p5_tuple_94852_comb[824:792];
  assign p5_tuple_index_95684_comb = p5_tuple_94852_comb[791:759];
  assign p5_tuple_index_95687_comb = p5_tuple_94852_comb[758:726];
  assign p5_tuple_index_95690_comb = p5_tuple_94852_comb[725:693];
  assign p5_tuple_index_95693_comb = p5_tuple_94852_comb[692:660];
  assign p5_tuple_index_95696_comb = p5_tuple_94852_comb[659:627];
  assign p5_tuple_index_95699_comb = p5_tuple_94852_comb[626:594];
  assign p5_tuple_index_95702_comb = p5_tuple_94852_comb[593:561];
  assign p5_tuple_index_95705_comb = p5_tuple_94852_comb[560:528];
  assign p5_tuple_index_95708_comb = p5_tuple_94852_comb[527:495];
  assign p5_tuple_index_95711_comb = p5_tuple_94852_comb[494:462];
  assign p5_tuple_index_95714_comb = p5_tuple_94852_comb[461:429];
  assign p5_tuple_index_95717_comb = p5_tuple_94852_comb[428:396];
  assign p5_tuple_index_95720_comb = p5_tuple_94852_comb[395:363];
  assign p5_tuple_index_95723_comb = p5_tuple_94852_comb[362:330];
  assign p5_tuple_index_95726_comb = p5_tuple_94852_comb[329:297];
  assign p5_tuple_index_95729_comb = p5_tuple_94852_comb[296:264];
  assign p5_tuple_index_95732_comb = p5_tuple_94852_comb[263:231];
  assign p5_tuple_index_95735_comb = p5_tuple_94852_comb[230:198];
  assign p5_tuple_index_95738_comb = p5_tuple_94852_comb[197:165];
  assign p5_tuple_index_95741_comb = p5_tuple_94852_comb[164:132];
  assign p5_tuple_index_95744_comb = p5_tuple_94852_comb[131:99];
  assign p5_tuple_index_95747_comb = p5_tuple_94852_comb[98:66];
  assign p5_tuple_index_95750_comb = p5_tuple_94852_comb[65:33];
  assign p5_tuple_index_95753_comb = p5_tuple_94852_comb[32:0];

  // Registers for pipe stage 5:
  reg p5_tuple_94852_index1;
  reg p5_tuple_94852_index2;
  reg p5_tuple_94852_index3;
  reg p5_tuple_94852_index4;
  reg p5_tuple_94852_index5;
  reg p5_tuple_94852_index6;
  reg p5_tuple_94852_index7;
  reg p5_tuple_94852_index8;
  reg p5_tuple_94852_index9;
  reg p5_tuple_94852_index10;
  reg p5_tuple_94852_index11;
  reg p5_tuple_94852_index12;
  reg p5_tuple_94852_index13;
  reg p5_tuple_94852_index14;
  reg p5_tuple_94852_index15;
  reg p5_tuple_94852_index16;
  reg p5_tuple_94852_index17;
  reg p5_tuple_94852_index18;
  reg p5_tuple_94852_index19;
  reg p5_tuple_94852_index20;
  reg p5_tuple_94852_index21;
  reg p5_tuple_94852_index22;
  reg p5_tuple_94852_index23;
  reg p5_tuple_94852_index24;
  reg p5_tuple_94852_index25;
  reg p5_tuple_94852_index26;
  reg p5_tuple_94852_index27;
  reg p5_tuple_94852_index28;
  reg p5_tuple_94852_index29;
  reg p5_tuple_94852_index30;
  reg p5_tuple_94852_index31;
  reg p5_tuple_94852_index32;
  reg p5_tuple_94852_index33;
  reg p5_tuple_94852_index34;
  reg p5_tuple_94852_index35;
  reg p5_tuple_94852_index36;
  reg p5_tuple_94852_index37;
  reg p5_tuple_94852_index38;
  reg p5_tuple_94852_index39;
  reg p5_tuple_94852_index40;
  reg p5_tuple_94852_index41;
  reg p5_tuple_94852_index42;
  reg p5_tuple_94852_index43;
  reg p5_tuple_94852_index44;
  reg p5_tuple_94852_index45;
  reg p5_tuple_94852_index46;
  reg p5_tuple_94852_index47;
  reg p5_tuple_94852_index48;
  reg p5_tuple_94852_index49;
  reg p5_tuple_94852_index50;
  reg p5_tuple_94852_index51;
  reg p5_tuple_94852_index52;
  reg p5_tuple_94852_index53;
  reg p5_tuple_94852_index54;
  reg p5_tuple_94852_index55;
  reg p5_tuple_94852_index56;
  reg p5_tuple_94852_index57;
  reg p5_tuple_94852_index58;
  reg p5_tuple_94852_index59;
  reg p5_tuple_94852_index60;
  reg p5_tuple_94852_index61;
  reg p5_tuple_94852_index62;
  reg p5_tuple_94852_index63;
  reg p5_tuple_94852_index64;
  reg p5_tuple_94852_index65;
  reg p5_tuple_94852_index66;
  reg p5_tuple_94852_index67;
  reg p5_tuple_94852_index68;
  reg p5_tuple_94852_index69;
  reg p5_tuple_94852_index70;
  reg p5_tuple_94852_index71;
  reg p5_tuple_94852_index72;
  reg p5_tuple_94852_index73;
  reg p5_tuple_94852_index74;
  reg p5_tuple_94852_index75;
  reg p5_tuple_94852_index76;
  reg p5_tuple_94852_index77;
  reg p5_tuple_94852_index78;
  reg p5_tuple_94852_index79;
  reg p5_tuple_94852_index80;
  reg p5_tuple_94852_index81;
  reg p5_tuple_94852_index82;
  reg p5_tuple_94852_index83;
  reg p5_tuple_94852_index84;
  reg p5_tuple_94852_index85;
  reg p5_tuple_94852_index86;
  reg p5_tuple_94852_index87;
  reg p5_tuple_94852_index88;
  reg p5_tuple_94852_index89;
  reg p5_tuple_94852_index90;
  reg p5_tuple_94852_index91;
  reg p5_tuple_94852_index92;
  reg p5_tuple_94852_index93;
  reg p5_tuple_94852_index94;
  reg p5_tuple_94852_index95;
  reg p5_tuple_94852_index96;
  reg p5_tuple_94852_index97;
  reg p5_tuple_94852_index98;
  reg p5_tuple_94852_index99;
  reg p5_tuple_94852_index100;
  reg p5_tuple_94852_index101;
  reg p5_tuple_94852_index102;
  reg p5_tuple_94852_index103;
  reg p5_tuple_94852_index104;
  reg p5_tuple_94852_index105;
  reg p5_tuple_94852_index106;
  reg p5_tuple_94852_index107;
  reg p5_tuple_94852_index108;
  reg p5_tuple_94852_index109;
  reg p5_tuple_94852_index110;
  reg p5_tuple_94852_index111;
  reg p5_tuple_94852_index112;
  reg p5_tuple_94852_index113;
  reg p5_tuple_94852_index114;
  reg p5_tuple_94852_index115;
  reg p5_tuple_94852_index116;
  reg p5_tuple_94852_index117;
  reg p5_tuple_94852_index118;
  reg p5_tuple_94852_index119;
  reg p5_tuple_94852_index120;
  reg p5_tuple_94852_index121;
  reg p5_tuple_94852_index122;
  reg p5_tuple_94852_index123;
  reg p5_tuple_94852_index124;
  reg p5_tuple_94852_index125;
  reg p5_tuple_94852_index126;
  reg p5_tuple_94852_index127;
  reg p5_tuple_94852_index128;
  reg p5_tuple_94852_index129;
  reg p5_tuple_94852_index130;
  reg p5_tuple_94852_index131;
  reg p5_tuple_94852_index132;
  reg p5_tuple_94852_index133;
  reg p5_tuple_94852_index134;
  reg p5_tuple_94852_index135;
  reg p5_tuple_94852_index136;
  reg p5_tuple_94852_index137;
  reg p5_tuple_94852_index138;
  reg p5_tuple_94852_index139;
  reg p5_tuple_94852_index140;
  reg p5_tuple_94852_index141;
  reg p5_tuple_94852_index142;
  reg p5_tuple_94852_index143;
  reg p5_tuple_94852_index144;
  reg p5_tuple_94852_index145;
  reg p5_tuple_94852_index146;
  reg p5_tuple_94852_index147;
  reg p5_tuple_94852_index148;
  reg p5_tuple_94852_index149;
  reg p5_tuple_94852_index150;
  reg p5_tuple_94852_index151;
  reg p5_tuple_94852_index152;
  reg p5_tuple_94852_index153;
  reg p5_tuple_94852_index154;
  reg p5_tuple_94852_index155;
  reg p5_tuple_94852_index156;
  reg p5_tuple_94852_index157;
  reg p5_tuple_94852_index158;
  reg p5_tuple_94852_index159;
  reg p5_tuple_94852_index160;
  reg p5_tuple_94852_index161;
  reg p5_tuple_94852_index162;
  reg p5_tuple_94852_index163;
  reg p5_tuple_94852_index164;
  reg p5_tuple_94852_index165;
  reg p5_tuple_94852_index166;
  reg p5_tuple_94852_index167;
  reg p5_tuple_94852_index168;
  reg p5_tuple_94852_index169;
  reg p5_tuple_94852_index170;
  reg p5_tuple_94852_index171;
  reg p5_tuple_94852_index172;
  reg p5_tuple_94852_index173;
  reg p5_tuple_94852_index174;
  reg p5_tuple_94852_index175;
  reg p5_tuple_94852_index176;
  reg p5_tuple_94852_index177;
  reg p5_tuple_94852_index178;
  reg p5_tuple_94852_index179;
  reg p5_tuple_94852_index180;
  reg p5_tuple_94852_index181;
  reg p5_tuple_94852_index182;
  reg p5_tuple_94852_index183;
  reg p5_tuple_94852_index184;
  reg p5_tuple_94852_index185;
  reg p5_tuple_94852_index186;
  reg p5_tuple_94852_index187;
  reg p5_tuple_94852_index188;
  reg p5_tuple_94852_index189;
  reg p5_tuple_94852_index190;
  reg p5_tuple_94852_index191;
  reg p5_tuple_94852_index192;
  reg p5_tuple_94852_index193;
  reg p5_tuple_94852_index194;
  reg p5_tuple_94852_index195;
  reg p5_tuple_94852_index196;
  reg p5_tuple_94852_index197;
  reg p5_tuple_94852_index198;
  reg p5_tuple_94852_index199;
  reg p5_tuple_94852_index200;
  reg [32:0] p5_tuple_94852_index201;
  reg [32:0] p5_tuple_94852_index202;
  reg [32:0] p5_tuple_94852_index203;
  reg [32:0] p5_tuple_94852_index204;
  reg [32:0] p5_tuple_94852_index205;
  reg [32:0] p5_tuple_94852_index206;
  reg [32:0] p5_tuple_94852_index207;
  reg [32:0] p5_tuple_94852_index208;
  reg [32:0] p5_tuple_94852_index209;
  reg [32:0] p5_tuple_94852_index210;
  reg [32:0] p5_tuple_94852_index211;
  reg [32:0] p5_tuple_94852_index212;
  reg [32:0] p5_tuple_94852_index213;
  reg [32:0] p5_tuple_94852_index214;
  reg [32:0] p5_tuple_94852_index215;
  reg [32:0] p5_tuple_94852_index216;
  reg [32:0] p5_tuple_94852_index217;
  reg [32:0] p5_tuple_94852_index218;
  reg [32:0] p5_tuple_94852_index219;
  reg [32:0] p5_tuple_94852_index220;
  reg [32:0] p5_tuple_94852_index221;
  reg [32:0] p5_tuple_94852_index222;
  reg [32:0] p5_tuple_94852_index223;
  reg [32:0] p5_tuple_94852_index224;
  reg [32:0] p5_tuple_94852_index225;
  reg [32:0] p5_tuple_94852_index226;
  reg [32:0] p5_tuple_94852_index227;
  reg [32:0] p5_tuple_94852_index228;
  reg [32:0] p5_tuple_94852_index229;
  reg [32:0] p5_tuple_94852_index230;
  reg [32:0] p5_tuple_94852_index231;
  reg [32:0] p5_tuple_94852_index232;
  reg [32:0] p5_tuple_94852_index233;
  reg [32:0] p5_tuple_94852_index234;
  reg [32:0] p5_tuple_94852_index235;
  reg [32:0] p5_tuple_94852_index236;
  reg [32:0] p5_tuple_94852_index237;
  reg [32:0] p5_tuple_94852_index238;
  reg [32:0] p5_tuple_94852_index239;
  reg [32:0] p5_tuple_94852_index240;
  reg [32:0] p5_tuple_94852_index241;
  reg [32:0] p5_tuple_94852_index242;
  reg [32:0] p5_tuple_94852_index243;
  reg [32:0] p5_tuple_94852_index244;
  reg [32:0] p5_tuple_94852_index245;
  reg [32:0] p5_tuple_94852_index246;
  reg [32:0] p5_tuple_94852_index247;
  reg [32:0] p5_tuple_94852_index248;
  reg [32:0] p5_tuple_94852_index249;
  reg [32:0] p5_tuple_94852_index250;
  reg [32:0] p5_tuple_94852_index251;
  reg [32:0] p5_tuple_94852_index252;
  reg [32:0] p5_tuple_94852_index253;
  reg [32:0] p5_tuple_94852_index254;
  reg [32:0] p5_tuple_94852_index255;
  reg [32:0] p5_tuple_94852_index256;
  reg [32:0] p5_tuple_94852_index257;
  reg [32:0] p5_tuple_94852_index258;
  reg [32:0] p5_tuple_94852_index259;
  reg [32:0] p5_tuple_94852_index260;
  reg [32:0] p5_tuple_94852_index261;
  reg [32:0] p5_tuple_94852_index262;
  reg [32:0] p5_tuple_94852_index263;
  reg [32:0] p5_tuple_94852_index264;
  reg [32:0] p5_tuple_94852_index265;
  reg [32:0] p5_tuple_94852_index266;
  reg [32:0] p5_tuple_94852_index267;
  reg [32:0] p5_tuple_94852_index268;
  reg [32:0] p5_tuple_94852_index269;
  reg [32:0] p5_tuple_94852_index270;
  reg [32:0] p5_tuple_94852_index271;
  reg [32:0] p5_tuple_94852_index272;
  reg [32:0] p5_tuple_94852_index273;
  reg [32:0] p5_tuple_94852_index274;
  reg [32:0] p5_tuple_94852_index275;
  reg [32:0] p5_tuple_94852_index276;
  reg [32:0] p5_tuple_94852_index277;
  reg [32:0] p5_tuple_94852_index278;
  reg [32:0] p5_tuple_94852_index279;
  reg [32:0] p5_tuple_94852_index280;
  reg [32:0] p5_tuple_94852_index281;
  reg [32:0] p5_tuple_94852_index282;
  reg [32:0] p5_tuple_94852_index283;
  reg [32:0] p5_tuple_94852_index284;
  reg [32:0] p5_tuple_94852_index285;
  reg [32:0] p5_tuple_94852_index286;
  reg [32:0] p5_tuple_94852_index287;
  reg [32:0] p5_tuple_94852_index288;
  reg [32:0] p5_tuple_94852_index289;
  reg [32:0] p5_tuple_94852_index290;
  reg [32:0] p5_tuple_94852_index291;
  reg [32:0] p5_tuple_94852_index292;
  reg [32:0] p5_tuple_94852_index293;
  reg [32:0] p5_tuple_94852_index294;
  reg [32:0] p5_tuple_94852_index295;
  reg [32:0] p5_tuple_94852_index296;
  reg [32:0] p5_tuple_94852_index297;
  reg [32:0] p5_tuple_94852_index298;
  reg [32:0] p5_tuple_94852_index299;
  reg [32:0] p5_tuple_94852_index300;
  always_ff @ (posedge clk) begin
    p5_tuple_94852_index1 <= p5_tuple_index_94856_comb;
    p5_tuple_94852_index2 <= p5_tuple_index_94859_comb;
    p5_tuple_94852_index3 <= p5_tuple_index_94862_comb;
    p5_tuple_94852_index4 <= p5_tuple_index_94865_comb;
    p5_tuple_94852_index5 <= p5_tuple_index_94868_comb;
    p5_tuple_94852_index6 <= p5_tuple_index_94871_comb;
    p5_tuple_94852_index7 <= p5_tuple_index_94874_comb;
    p5_tuple_94852_index8 <= p5_tuple_index_94877_comb;
    p5_tuple_94852_index9 <= p5_tuple_index_94880_comb;
    p5_tuple_94852_index10 <= p5_tuple_index_94883_comb;
    p5_tuple_94852_index11 <= p5_tuple_index_94886_comb;
    p5_tuple_94852_index12 <= p5_tuple_index_94889_comb;
    p5_tuple_94852_index13 <= p5_tuple_index_94892_comb;
    p5_tuple_94852_index14 <= p5_tuple_index_94895_comb;
    p5_tuple_94852_index15 <= p5_tuple_index_94898_comb;
    p5_tuple_94852_index16 <= p5_tuple_index_94901_comb;
    p5_tuple_94852_index17 <= p5_tuple_index_94904_comb;
    p5_tuple_94852_index18 <= p5_tuple_index_94907_comb;
    p5_tuple_94852_index19 <= p5_tuple_index_94910_comb;
    p5_tuple_94852_index20 <= p5_tuple_index_94913_comb;
    p5_tuple_94852_index21 <= p5_tuple_index_94916_comb;
    p5_tuple_94852_index22 <= p5_tuple_index_94919_comb;
    p5_tuple_94852_index23 <= p5_tuple_index_94922_comb;
    p5_tuple_94852_index24 <= p5_tuple_index_94925_comb;
    p5_tuple_94852_index25 <= p5_tuple_index_94928_comb;
    p5_tuple_94852_index26 <= p5_tuple_index_94931_comb;
    p5_tuple_94852_index27 <= p5_tuple_index_94934_comb;
    p5_tuple_94852_index28 <= p5_tuple_index_94937_comb;
    p5_tuple_94852_index29 <= p5_tuple_index_94940_comb;
    p5_tuple_94852_index30 <= p5_tuple_index_94943_comb;
    p5_tuple_94852_index31 <= p5_tuple_index_94946_comb;
    p5_tuple_94852_index32 <= p5_tuple_index_94949_comb;
    p5_tuple_94852_index33 <= p5_tuple_index_94952_comb;
    p5_tuple_94852_index34 <= p5_tuple_index_94955_comb;
    p5_tuple_94852_index35 <= p5_tuple_index_94958_comb;
    p5_tuple_94852_index36 <= p5_tuple_index_94961_comb;
    p5_tuple_94852_index37 <= p5_tuple_index_94964_comb;
    p5_tuple_94852_index38 <= p5_tuple_index_94967_comb;
    p5_tuple_94852_index39 <= p5_tuple_index_94970_comb;
    p5_tuple_94852_index40 <= p5_tuple_index_94973_comb;
    p5_tuple_94852_index41 <= p5_tuple_index_94976_comb;
    p5_tuple_94852_index42 <= p5_tuple_index_94979_comb;
    p5_tuple_94852_index43 <= p5_tuple_index_94982_comb;
    p5_tuple_94852_index44 <= p5_tuple_index_94985_comb;
    p5_tuple_94852_index45 <= p5_tuple_index_94988_comb;
    p5_tuple_94852_index46 <= p5_tuple_index_94991_comb;
    p5_tuple_94852_index47 <= p5_tuple_index_94994_comb;
    p5_tuple_94852_index48 <= p5_tuple_index_94997_comb;
    p5_tuple_94852_index49 <= p5_tuple_index_95000_comb;
    p5_tuple_94852_index50 <= p5_tuple_index_95003_comb;
    p5_tuple_94852_index51 <= p5_tuple_index_95006_comb;
    p5_tuple_94852_index52 <= p5_tuple_index_95009_comb;
    p5_tuple_94852_index53 <= p5_tuple_index_95012_comb;
    p5_tuple_94852_index54 <= p5_tuple_index_95015_comb;
    p5_tuple_94852_index55 <= p5_tuple_index_95018_comb;
    p5_tuple_94852_index56 <= p5_tuple_index_95021_comb;
    p5_tuple_94852_index57 <= p5_tuple_index_95024_comb;
    p5_tuple_94852_index58 <= p5_tuple_index_95027_comb;
    p5_tuple_94852_index59 <= p5_tuple_index_95030_comb;
    p5_tuple_94852_index60 <= p5_tuple_index_95033_comb;
    p5_tuple_94852_index61 <= p5_tuple_index_95036_comb;
    p5_tuple_94852_index62 <= p5_tuple_index_95039_comb;
    p5_tuple_94852_index63 <= p5_tuple_index_95042_comb;
    p5_tuple_94852_index64 <= p5_tuple_index_95045_comb;
    p5_tuple_94852_index65 <= p5_tuple_index_95048_comb;
    p5_tuple_94852_index66 <= p5_tuple_index_95051_comb;
    p5_tuple_94852_index67 <= p5_tuple_index_95054_comb;
    p5_tuple_94852_index68 <= p5_tuple_index_95057_comb;
    p5_tuple_94852_index69 <= p5_tuple_index_95060_comb;
    p5_tuple_94852_index70 <= p5_tuple_index_95063_comb;
    p5_tuple_94852_index71 <= p5_tuple_index_95066_comb;
    p5_tuple_94852_index72 <= p5_tuple_index_95069_comb;
    p5_tuple_94852_index73 <= p5_tuple_index_95072_comb;
    p5_tuple_94852_index74 <= p5_tuple_index_95075_comb;
    p5_tuple_94852_index75 <= p5_tuple_index_95078_comb;
    p5_tuple_94852_index76 <= p5_tuple_index_95081_comb;
    p5_tuple_94852_index77 <= p5_tuple_index_95084_comb;
    p5_tuple_94852_index78 <= p5_tuple_index_95087_comb;
    p5_tuple_94852_index79 <= p5_tuple_index_95090_comb;
    p5_tuple_94852_index80 <= p5_tuple_index_95093_comb;
    p5_tuple_94852_index81 <= p5_tuple_index_95096_comb;
    p5_tuple_94852_index82 <= p5_tuple_index_95099_comb;
    p5_tuple_94852_index83 <= p5_tuple_index_95102_comb;
    p5_tuple_94852_index84 <= p5_tuple_index_95105_comb;
    p5_tuple_94852_index85 <= p5_tuple_index_95108_comb;
    p5_tuple_94852_index86 <= p5_tuple_index_95111_comb;
    p5_tuple_94852_index87 <= p5_tuple_index_95114_comb;
    p5_tuple_94852_index88 <= p5_tuple_index_95117_comb;
    p5_tuple_94852_index89 <= p5_tuple_index_95120_comb;
    p5_tuple_94852_index90 <= p5_tuple_index_95123_comb;
    p5_tuple_94852_index91 <= p5_tuple_index_95126_comb;
    p5_tuple_94852_index92 <= p5_tuple_index_95129_comb;
    p5_tuple_94852_index93 <= p5_tuple_index_95132_comb;
    p5_tuple_94852_index94 <= p5_tuple_index_95135_comb;
    p5_tuple_94852_index95 <= p5_tuple_index_95138_comb;
    p5_tuple_94852_index96 <= p5_tuple_index_95141_comb;
    p5_tuple_94852_index97 <= p5_tuple_index_95144_comb;
    p5_tuple_94852_index98 <= p5_tuple_index_95147_comb;
    p5_tuple_94852_index99 <= p5_tuple_index_95150_comb;
    p5_tuple_94852_index100 <= p5_tuple_index_95153_comb;
    p5_tuple_94852_index101 <= p5_tuple_index_95156_comb;
    p5_tuple_94852_index102 <= p5_tuple_index_95159_comb;
    p5_tuple_94852_index103 <= p5_tuple_index_95162_comb;
    p5_tuple_94852_index104 <= p5_tuple_index_95165_comb;
    p5_tuple_94852_index105 <= p5_tuple_index_95168_comb;
    p5_tuple_94852_index106 <= p5_tuple_index_95171_comb;
    p5_tuple_94852_index107 <= p5_tuple_index_95174_comb;
    p5_tuple_94852_index108 <= p5_tuple_index_95177_comb;
    p5_tuple_94852_index109 <= p5_tuple_index_95180_comb;
    p5_tuple_94852_index110 <= p5_tuple_index_95183_comb;
    p5_tuple_94852_index111 <= p5_tuple_index_95186_comb;
    p5_tuple_94852_index112 <= p5_tuple_index_95189_comb;
    p5_tuple_94852_index113 <= p5_tuple_index_95192_comb;
    p5_tuple_94852_index114 <= p5_tuple_index_95195_comb;
    p5_tuple_94852_index115 <= p5_tuple_index_95198_comb;
    p5_tuple_94852_index116 <= p5_tuple_index_95201_comb;
    p5_tuple_94852_index117 <= p5_tuple_index_95204_comb;
    p5_tuple_94852_index118 <= p5_tuple_index_95207_comb;
    p5_tuple_94852_index119 <= p5_tuple_index_95210_comb;
    p5_tuple_94852_index120 <= p5_tuple_index_95213_comb;
    p5_tuple_94852_index121 <= p5_tuple_index_95216_comb;
    p5_tuple_94852_index122 <= p5_tuple_index_95219_comb;
    p5_tuple_94852_index123 <= p5_tuple_index_95222_comb;
    p5_tuple_94852_index124 <= p5_tuple_index_95225_comb;
    p5_tuple_94852_index125 <= p5_tuple_index_95228_comb;
    p5_tuple_94852_index126 <= p5_tuple_index_95231_comb;
    p5_tuple_94852_index127 <= p5_tuple_index_95234_comb;
    p5_tuple_94852_index128 <= p5_tuple_index_95237_comb;
    p5_tuple_94852_index129 <= p5_tuple_index_95240_comb;
    p5_tuple_94852_index130 <= p5_tuple_index_95243_comb;
    p5_tuple_94852_index131 <= p5_tuple_index_95246_comb;
    p5_tuple_94852_index132 <= p5_tuple_index_95249_comb;
    p5_tuple_94852_index133 <= p5_tuple_index_95252_comb;
    p5_tuple_94852_index134 <= p5_tuple_index_95255_comb;
    p5_tuple_94852_index135 <= p5_tuple_index_95258_comb;
    p5_tuple_94852_index136 <= p5_tuple_index_95261_comb;
    p5_tuple_94852_index137 <= p5_tuple_index_95264_comb;
    p5_tuple_94852_index138 <= p5_tuple_index_95267_comb;
    p5_tuple_94852_index139 <= p5_tuple_index_95270_comb;
    p5_tuple_94852_index140 <= p5_tuple_index_95273_comb;
    p5_tuple_94852_index141 <= p5_tuple_index_95276_comb;
    p5_tuple_94852_index142 <= p5_tuple_index_95279_comb;
    p5_tuple_94852_index143 <= p5_tuple_index_95282_comb;
    p5_tuple_94852_index144 <= p5_tuple_index_95285_comb;
    p5_tuple_94852_index145 <= p5_tuple_index_95288_comb;
    p5_tuple_94852_index146 <= p5_tuple_index_95291_comb;
    p5_tuple_94852_index147 <= p5_tuple_index_95294_comb;
    p5_tuple_94852_index148 <= p5_tuple_index_95297_comb;
    p5_tuple_94852_index149 <= p5_tuple_index_95300_comb;
    p5_tuple_94852_index150 <= p5_tuple_index_95303_comb;
    p5_tuple_94852_index151 <= p5_tuple_index_95306_comb;
    p5_tuple_94852_index152 <= p5_tuple_index_95309_comb;
    p5_tuple_94852_index153 <= p5_tuple_index_95312_comb;
    p5_tuple_94852_index154 <= p5_tuple_index_95315_comb;
    p5_tuple_94852_index155 <= p5_tuple_index_95318_comb;
    p5_tuple_94852_index156 <= p5_tuple_index_95321_comb;
    p5_tuple_94852_index157 <= p5_tuple_index_95324_comb;
    p5_tuple_94852_index158 <= p5_tuple_index_95327_comb;
    p5_tuple_94852_index159 <= p5_tuple_index_95330_comb;
    p5_tuple_94852_index160 <= p5_tuple_index_95333_comb;
    p5_tuple_94852_index161 <= p5_tuple_index_95336_comb;
    p5_tuple_94852_index162 <= p5_tuple_index_95339_comb;
    p5_tuple_94852_index163 <= p5_tuple_index_95342_comb;
    p5_tuple_94852_index164 <= p5_tuple_index_95345_comb;
    p5_tuple_94852_index165 <= p5_tuple_index_95348_comb;
    p5_tuple_94852_index166 <= p5_tuple_index_95351_comb;
    p5_tuple_94852_index167 <= p5_tuple_index_95354_comb;
    p5_tuple_94852_index168 <= p5_tuple_index_95357_comb;
    p5_tuple_94852_index169 <= p5_tuple_index_95360_comb;
    p5_tuple_94852_index170 <= p5_tuple_index_95363_comb;
    p5_tuple_94852_index171 <= p5_tuple_index_95366_comb;
    p5_tuple_94852_index172 <= p5_tuple_index_95369_comb;
    p5_tuple_94852_index173 <= p5_tuple_index_95372_comb;
    p5_tuple_94852_index174 <= p5_tuple_index_95375_comb;
    p5_tuple_94852_index175 <= p5_tuple_index_95378_comb;
    p5_tuple_94852_index176 <= p5_tuple_index_95381_comb;
    p5_tuple_94852_index177 <= p5_tuple_index_95384_comb;
    p5_tuple_94852_index178 <= p5_tuple_index_95387_comb;
    p5_tuple_94852_index179 <= p5_tuple_index_95390_comb;
    p5_tuple_94852_index180 <= p5_tuple_index_95393_comb;
    p5_tuple_94852_index181 <= p5_tuple_index_95396_comb;
    p5_tuple_94852_index182 <= p5_tuple_index_95399_comb;
    p5_tuple_94852_index183 <= p5_tuple_index_95402_comb;
    p5_tuple_94852_index184 <= p5_tuple_index_95405_comb;
    p5_tuple_94852_index185 <= p5_tuple_index_95408_comb;
    p5_tuple_94852_index186 <= p5_tuple_index_95411_comb;
    p5_tuple_94852_index187 <= p5_tuple_index_95414_comb;
    p5_tuple_94852_index188 <= p5_tuple_index_95417_comb;
    p5_tuple_94852_index189 <= p5_tuple_index_95420_comb;
    p5_tuple_94852_index190 <= p5_tuple_index_95423_comb;
    p5_tuple_94852_index191 <= p5_tuple_index_95426_comb;
    p5_tuple_94852_index192 <= p5_tuple_index_95429_comb;
    p5_tuple_94852_index193 <= p5_tuple_index_95432_comb;
    p5_tuple_94852_index194 <= p5_tuple_index_95435_comb;
    p5_tuple_94852_index195 <= p5_tuple_index_95438_comb;
    p5_tuple_94852_index196 <= p5_tuple_index_95441_comb;
    p5_tuple_94852_index197 <= p5_tuple_index_95444_comb;
    p5_tuple_94852_index198 <= p5_tuple_index_95447_comb;
    p5_tuple_94852_index199 <= p5_tuple_index_95450_comb;
    p5_tuple_94852_index200 <= p5_tuple_index_95453_comb;
    p5_tuple_94852_index201 <= p5_tuple_index_95456_comb;
    p5_tuple_94852_index202 <= p5_tuple_index_95459_comb;
    p5_tuple_94852_index203 <= p5_tuple_index_95462_comb;
    p5_tuple_94852_index204 <= p5_tuple_index_95465_comb;
    p5_tuple_94852_index205 <= p5_tuple_index_95468_comb;
    p5_tuple_94852_index206 <= p5_tuple_index_95471_comb;
    p5_tuple_94852_index207 <= p5_tuple_index_95474_comb;
    p5_tuple_94852_index208 <= p5_tuple_index_95477_comb;
    p5_tuple_94852_index209 <= p5_tuple_index_95480_comb;
    p5_tuple_94852_index210 <= p5_tuple_index_95483_comb;
    p5_tuple_94852_index211 <= p5_tuple_index_95486_comb;
    p5_tuple_94852_index212 <= p5_tuple_index_95489_comb;
    p5_tuple_94852_index213 <= p5_tuple_index_95492_comb;
    p5_tuple_94852_index214 <= p5_tuple_index_95495_comb;
    p5_tuple_94852_index215 <= p5_tuple_index_95498_comb;
    p5_tuple_94852_index216 <= p5_tuple_index_95501_comb;
    p5_tuple_94852_index217 <= p5_tuple_index_95504_comb;
    p5_tuple_94852_index218 <= p5_tuple_index_95507_comb;
    p5_tuple_94852_index219 <= p5_tuple_index_95510_comb;
    p5_tuple_94852_index220 <= p5_tuple_index_95513_comb;
    p5_tuple_94852_index221 <= p5_tuple_index_95516_comb;
    p5_tuple_94852_index222 <= p5_tuple_index_95519_comb;
    p5_tuple_94852_index223 <= p5_tuple_index_95522_comb;
    p5_tuple_94852_index224 <= p5_tuple_index_95525_comb;
    p5_tuple_94852_index225 <= p5_tuple_index_95528_comb;
    p5_tuple_94852_index226 <= p5_tuple_index_95531_comb;
    p5_tuple_94852_index227 <= p5_tuple_index_95534_comb;
    p5_tuple_94852_index228 <= p5_tuple_index_95537_comb;
    p5_tuple_94852_index229 <= p5_tuple_index_95540_comb;
    p5_tuple_94852_index230 <= p5_tuple_index_95543_comb;
    p5_tuple_94852_index231 <= p5_tuple_index_95546_comb;
    p5_tuple_94852_index232 <= p5_tuple_index_95549_comb;
    p5_tuple_94852_index233 <= p5_tuple_index_95552_comb;
    p5_tuple_94852_index234 <= p5_tuple_index_95555_comb;
    p5_tuple_94852_index235 <= p5_tuple_index_95558_comb;
    p5_tuple_94852_index236 <= p5_tuple_index_95561_comb;
    p5_tuple_94852_index237 <= p5_tuple_index_95564_comb;
    p5_tuple_94852_index238 <= p5_tuple_index_95567_comb;
    p5_tuple_94852_index239 <= p5_tuple_index_95570_comb;
    p5_tuple_94852_index240 <= p5_tuple_index_95573_comb;
    p5_tuple_94852_index241 <= p5_tuple_index_95576_comb;
    p5_tuple_94852_index242 <= p5_tuple_index_95579_comb;
    p5_tuple_94852_index243 <= p5_tuple_index_95582_comb;
    p5_tuple_94852_index244 <= p5_tuple_index_95585_comb;
    p5_tuple_94852_index245 <= p5_tuple_index_95588_comb;
    p5_tuple_94852_index246 <= p5_tuple_index_95591_comb;
    p5_tuple_94852_index247 <= p5_tuple_index_95594_comb;
    p5_tuple_94852_index248 <= p5_tuple_index_95597_comb;
    p5_tuple_94852_index249 <= p5_tuple_index_95600_comb;
    p5_tuple_94852_index250 <= p5_tuple_index_95603_comb;
    p5_tuple_94852_index251 <= p5_tuple_index_95606_comb;
    p5_tuple_94852_index252 <= p5_tuple_index_95609_comb;
    p5_tuple_94852_index253 <= p5_tuple_index_95612_comb;
    p5_tuple_94852_index254 <= p5_tuple_index_95615_comb;
    p5_tuple_94852_index255 <= p5_tuple_index_95618_comb;
    p5_tuple_94852_index256 <= p5_tuple_index_95621_comb;
    p5_tuple_94852_index257 <= p5_tuple_index_95624_comb;
    p5_tuple_94852_index258 <= p5_tuple_index_95627_comb;
    p5_tuple_94852_index259 <= p5_tuple_index_95630_comb;
    p5_tuple_94852_index260 <= p5_tuple_index_95633_comb;
    p5_tuple_94852_index261 <= p5_tuple_index_95636_comb;
    p5_tuple_94852_index262 <= p5_tuple_index_95639_comb;
    p5_tuple_94852_index263 <= p5_tuple_index_95642_comb;
    p5_tuple_94852_index264 <= p5_tuple_index_95645_comb;
    p5_tuple_94852_index265 <= p5_tuple_index_95648_comb;
    p5_tuple_94852_index266 <= p5_tuple_index_95651_comb;
    p5_tuple_94852_index267 <= p5_tuple_index_95654_comb;
    p5_tuple_94852_index268 <= p5_tuple_index_95657_comb;
    p5_tuple_94852_index269 <= p5_tuple_index_95660_comb;
    p5_tuple_94852_index270 <= p5_tuple_index_95663_comb;
    p5_tuple_94852_index271 <= p5_tuple_index_95666_comb;
    p5_tuple_94852_index272 <= p5_tuple_index_95669_comb;
    p5_tuple_94852_index273 <= p5_tuple_index_95672_comb;
    p5_tuple_94852_index274 <= p5_tuple_index_95675_comb;
    p5_tuple_94852_index275 <= p5_tuple_index_95678_comb;
    p5_tuple_94852_index276 <= p5_tuple_index_95681_comb;
    p5_tuple_94852_index277 <= p5_tuple_index_95684_comb;
    p5_tuple_94852_index278 <= p5_tuple_index_95687_comb;
    p5_tuple_94852_index279 <= p5_tuple_index_95690_comb;
    p5_tuple_94852_index280 <= p5_tuple_index_95693_comb;
    p5_tuple_94852_index281 <= p5_tuple_index_95696_comb;
    p5_tuple_94852_index282 <= p5_tuple_index_95699_comb;
    p5_tuple_94852_index283 <= p5_tuple_index_95702_comb;
    p5_tuple_94852_index284 <= p5_tuple_index_95705_comb;
    p5_tuple_94852_index285 <= p5_tuple_index_95708_comb;
    p5_tuple_94852_index286 <= p5_tuple_index_95711_comb;
    p5_tuple_94852_index287 <= p5_tuple_index_95714_comb;
    p5_tuple_94852_index288 <= p5_tuple_index_95717_comb;
    p5_tuple_94852_index289 <= p5_tuple_index_95720_comb;
    p5_tuple_94852_index290 <= p5_tuple_index_95723_comb;
    p5_tuple_94852_index291 <= p5_tuple_index_95726_comb;
    p5_tuple_94852_index292 <= p5_tuple_index_95729_comb;
    p5_tuple_94852_index293 <= p5_tuple_index_95732_comb;
    p5_tuple_94852_index294 <= p5_tuple_index_95735_comb;
    p5_tuple_94852_index295 <= p5_tuple_index_95738_comb;
    p5_tuple_94852_index296 <= p5_tuple_index_95741_comb;
    p5_tuple_94852_index297 <= p5_tuple_index_95744_comb;
    p5_tuple_94852_index298 <= p5_tuple_index_95747_comb;
    p5_tuple_94852_index299 <= p5_tuple_index_95750_comb;
    p5_tuple_94852_index300 <= p5_tuple_index_95753_comb;
  end

  // ===== Pipe stage 6:
  assign out = {p5_tuple_94852_index1, p5_tuple_94852_index2, p5_tuple_94852_index3, p5_tuple_94852_index4, p5_tuple_94852_index5, p5_tuple_94852_index6, p5_tuple_94852_index7, p5_tuple_94852_index8, p5_tuple_94852_index9, p5_tuple_94852_index10, p5_tuple_94852_index11, p5_tuple_94852_index12, p5_tuple_94852_index13, p5_tuple_94852_index14, p5_tuple_94852_index15, p5_tuple_94852_index16, p5_tuple_94852_index17, p5_tuple_94852_index18, p5_tuple_94852_index19, p5_tuple_94852_index20, p5_tuple_94852_index21, p5_tuple_94852_index22, p5_tuple_94852_index23, p5_tuple_94852_index24, p5_tuple_94852_index25, p5_tuple_94852_index26, p5_tuple_94852_index27, p5_tuple_94852_index28, p5_tuple_94852_index29, p5_tuple_94852_index30, p5_tuple_94852_index31, p5_tuple_94852_index32, p5_tuple_94852_index33, p5_tuple_94852_index34, p5_tuple_94852_index35, p5_tuple_94852_index36, p5_tuple_94852_index37, p5_tuple_94852_index38, p5_tuple_94852_index39, p5_tuple_94852_index40, p5_tuple_94852_index41, p5_tuple_94852_index42, p5_tuple_94852_index43, p5_tuple_94852_index44, p5_tuple_94852_index45, p5_tuple_94852_index46, p5_tuple_94852_index47, p5_tuple_94852_index48, p5_tuple_94852_index49, p5_tuple_94852_index50, p5_tuple_94852_index51, p5_tuple_94852_index52, p5_tuple_94852_index53, p5_tuple_94852_index54, p5_tuple_94852_index55, p5_tuple_94852_index56, p5_tuple_94852_index57, p5_tuple_94852_index58, p5_tuple_94852_index59, p5_tuple_94852_index60, p5_tuple_94852_index61, p5_tuple_94852_index62, p5_tuple_94852_index63, p5_tuple_94852_index64, p5_tuple_94852_index65, p5_tuple_94852_index66, p5_tuple_94852_index67, p5_tuple_94852_index68, p5_tuple_94852_index69, p5_tuple_94852_index70, p5_tuple_94852_index71, p5_tuple_94852_index72, p5_tuple_94852_index73, p5_tuple_94852_index74, p5_tuple_94852_index75, p5_tuple_94852_index76, p5_tuple_94852_index77, p5_tuple_94852_index78, p5_tuple_94852_index79, p5_tuple_94852_index80, p5_tuple_94852_index81, p5_tuple_94852_index82, p5_tuple_94852_index83, p5_tuple_94852_index84, p5_tuple_94852_index85, p5_tuple_94852_index86, p5_tuple_94852_index87, p5_tuple_94852_index88, p5_tuple_94852_index89, p5_tuple_94852_index90, p5_tuple_94852_index91, p5_tuple_94852_index92, p5_tuple_94852_index93, p5_tuple_94852_index94, p5_tuple_94852_index95, p5_tuple_94852_index96, p5_tuple_94852_index97, p5_tuple_94852_index98, p5_tuple_94852_index99, p5_tuple_94852_index100, p5_tuple_94852_index101, p5_tuple_94852_index102, p5_tuple_94852_index103, p5_tuple_94852_index104, p5_tuple_94852_index105, p5_tuple_94852_index106, p5_tuple_94852_index107, p5_tuple_94852_index108, p5_tuple_94852_index109, p5_tuple_94852_index110, p5_tuple_94852_index111, p5_tuple_94852_index112, p5_tuple_94852_index113, p5_tuple_94852_index114, p5_tuple_94852_index115, p5_tuple_94852_index116, p5_tuple_94852_index117, p5_tuple_94852_index118, p5_tuple_94852_index119, p5_tuple_94852_index120, p5_tuple_94852_index121, p5_tuple_94852_index122, p5_tuple_94852_index123, p5_tuple_94852_index124, p5_tuple_94852_index125, p5_tuple_94852_index126, p5_tuple_94852_index127, p5_tuple_94852_index128, p5_tuple_94852_index129, p5_tuple_94852_index130, p5_tuple_94852_index131, p5_tuple_94852_index132, p5_tuple_94852_index133, p5_tuple_94852_index134, p5_tuple_94852_index135, p5_tuple_94852_index136, p5_tuple_94852_index137, p5_tuple_94852_index138, p5_tuple_94852_index139, p5_tuple_94852_index140, p5_tuple_94852_index141, p5_tuple_94852_index142, p5_tuple_94852_index143, p5_tuple_94852_index144, p5_tuple_94852_index145, p5_tuple_94852_index146, p5_tuple_94852_index147, p5_tuple_94852_index148, p5_tuple_94852_index149, p5_tuple_94852_index150, p5_tuple_94852_index151, p5_tuple_94852_index152, p5_tuple_94852_index153, p5_tuple_94852_index154, p5_tuple_94852_index155, p5_tuple_94852_index156, p5_tuple_94852_index157, p5_tuple_94852_index158, p5_tuple_94852_index159, p5_tuple_94852_index160, p5_tuple_94852_index161, p5_tuple_94852_index162, p5_tuple_94852_index163, p5_tuple_94852_index164, p5_tuple_94852_index165, p5_tuple_94852_index166, p5_tuple_94852_index167, p5_tuple_94852_index168, p5_tuple_94852_index169, p5_tuple_94852_index170, p5_tuple_94852_index171, p5_tuple_94852_index172, p5_tuple_94852_index173, p5_tuple_94852_index174, p5_tuple_94852_index175, p5_tuple_94852_index176, p5_tuple_94852_index177, p5_tuple_94852_index178, p5_tuple_94852_index179, p5_tuple_94852_index180, p5_tuple_94852_index181, p5_tuple_94852_index182, p5_tuple_94852_index183, p5_tuple_94852_index184, p5_tuple_94852_index185, p5_tuple_94852_index186, p5_tuple_94852_index187, p5_tuple_94852_index188, p5_tuple_94852_index189, p5_tuple_94852_index190, p5_tuple_94852_index191, p5_tuple_94852_index192, p5_tuple_94852_index193, p5_tuple_94852_index194, p5_tuple_94852_index195, p5_tuple_94852_index196, p5_tuple_94852_index197, p5_tuple_94852_index198, p5_tuple_94852_index199, p5_tuple_94852_index200, p5_tuple_94852_index201, p5_tuple_94852_index202, p5_tuple_94852_index203, p5_tuple_94852_index204, p5_tuple_94852_index205, p5_tuple_94852_index206, p5_tuple_94852_index207, p5_tuple_94852_index208, p5_tuple_94852_index209, p5_tuple_94852_index210, p5_tuple_94852_index211, p5_tuple_94852_index212, p5_tuple_94852_index213, p5_tuple_94852_index214, p5_tuple_94852_index215, p5_tuple_94852_index216, p5_tuple_94852_index217, p5_tuple_94852_index218, p5_tuple_94852_index219, p5_tuple_94852_index220, p5_tuple_94852_index221, p5_tuple_94852_index222, p5_tuple_94852_index223, p5_tuple_94852_index224, p5_tuple_94852_index225, p5_tuple_94852_index226, p5_tuple_94852_index227, p5_tuple_94852_index228, p5_tuple_94852_index229, p5_tuple_94852_index230, p5_tuple_94852_index231, p5_tuple_94852_index232, p5_tuple_94852_index233, p5_tuple_94852_index234, p5_tuple_94852_index235, p5_tuple_94852_index236, p5_tuple_94852_index237, p5_tuple_94852_index238, p5_tuple_94852_index239, p5_tuple_94852_index240, p5_tuple_94852_index241, p5_tuple_94852_index242, p5_tuple_94852_index243, p5_tuple_94852_index244, p5_tuple_94852_index245, p5_tuple_94852_index246, p5_tuple_94852_index247, p5_tuple_94852_index248, p5_tuple_94852_index249, p5_tuple_94852_index250, p5_tuple_94852_index251, p5_tuple_94852_index252, p5_tuple_94852_index253, p5_tuple_94852_index254, p5_tuple_94852_index255, p5_tuple_94852_index256, p5_tuple_94852_index257, p5_tuple_94852_index258, p5_tuple_94852_index259, p5_tuple_94852_index260, p5_tuple_94852_index261, p5_tuple_94852_index262, p5_tuple_94852_index263, p5_tuple_94852_index264, p5_tuple_94852_index265, p5_tuple_94852_index266, p5_tuple_94852_index267, p5_tuple_94852_index268, p5_tuple_94852_index269, p5_tuple_94852_index270, p5_tuple_94852_index271, p5_tuple_94852_index272, p5_tuple_94852_index273, p5_tuple_94852_index274, p5_tuple_94852_index275, p5_tuple_94852_index276, p5_tuple_94852_index277, p5_tuple_94852_index278, p5_tuple_94852_index279, p5_tuple_94852_index280, p5_tuple_94852_index281, p5_tuple_94852_index282, p5_tuple_94852_index283, p5_tuple_94852_index284, p5_tuple_94852_index285, p5_tuple_94852_index286, p5_tuple_94852_index287, p5_tuple_94852_index288, p5_tuple_94852_index289, p5_tuple_94852_index290, p5_tuple_94852_index291, p5_tuple_94852_index292, p5_tuple_94852_index293, p5_tuple_94852_index294, p5_tuple_94852_index295, p5_tuple_94852_index296, p5_tuple_94852_index297, p5_tuple_94852_index298, p5_tuple_94852_index299, p5_tuple_94852_index300};
endmodule
