module matrix_mul_10_pipeline(
  input wire clk,
  input wire [31:0] TestBlock__A_op0,
  input wire [31:0] TestBlock__A_op1,
  input wire [31:0] TestBlock__A_op2,
  input wire [31:0] TestBlock__A_op3,
  input wire [31:0] TestBlock__A_op4,
  input wire [31:0] TestBlock__A_op5,
  input wire [31:0] TestBlock__A_op6,
  input wire [31:0] TestBlock__A_op7,
  input wire [31:0] TestBlock__A_op8,
  input wire [31:0] TestBlock__A_op9,
  input wire [31:0] TestBlock__A_op10,
  input wire [31:0] TestBlock__A_op11,
  input wire [31:0] TestBlock__A_op12,
  input wire [31:0] TestBlock__A_op13,
  input wire [31:0] TestBlock__A_op14,
  input wire [31:0] TestBlock__A_op15,
  input wire [31:0] TestBlock__A_op16,
  input wire [31:0] TestBlock__A_op17,
  input wire [31:0] TestBlock__A_op18,
  input wire [31:0] TestBlock__A_op19,
  input wire [31:0] TestBlock__A_op20,
  input wire [31:0] TestBlock__A_op21,
  input wire [31:0] TestBlock__A_op22,
  input wire [31:0] TestBlock__A_op23,
  input wire [31:0] TestBlock__A_op24,
  input wire [31:0] TestBlock__A_op25,
  input wire [31:0] TestBlock__A_op26,
  input wire [31:0] TestBlock__A_op27,
  input wire [31:0] TestBlock__A_op28,
  input wire [31:0] TestBlock__A_op29,
  input wire [31:0] TestBlock__A_op30,
  input wire [31:0] TestBlock__A_op31,
  input wire [31:0] TestBlock__A_op32,
  input wire [31:0] TestBlock__A_op33,
  input wire [31:0] TestBlock__A_op34,
  input wire [31:0] TestBlock__A_op35,
  input wire [31:0] TestBlock__A_op36,
  input wire [31:0] TestBlock__A_op37,
  input wire [31:0] TestBlock__A_op38,
  input wire [31:0] TestBlock__A_op39,
  input wire [31:0] TestBlock__A_op40,
  input wire [31:0] TestBlock__A_op41,
  input wire [31:0] TestBlock__A_op42,
  input wire [31:0] TestBlock__A_op43,
  input wire [31:0] TestBlock__A_op44,
  input wire [31:0] TestBlock__A_op45,
  input wire [31:0] TestBlock__A_op46,
  input wire [31:0] TestBlock__A_op47,
  input wire [31:0] TestBlock__A_op48,
  input wire [31:0] TestBlock__A_op49,
  input wire [31:0] TestBlock__A_op50,
  input wire [31:0] TestBlock__A_op51,
  input wire [31:0] TestBlock__A_op52,
  input wire [31:0] TestBlock__A_op53,
  input wire [31:0] TestBlock__A_op54,
  input wire [31:0] TestBlock__A_op55,
  input wire [31:0] TestBlock__A_op56,
  input wire [31:0] TestBlock__A_op57,
  input wire [31:0] TestBlock__A_op58,
  input wire [31:0] TestBlock__A_op59,
  input wire [31:0] TestBlock__A_op60,
  input wire [31:0] TestBlock__A_op61,
  input wire [31:0] TestBlock__A_op62,
  input wire [31:0] TestBlock__A_op63,
  input wire [31:0] TestBlock__A_op64,
  input wire [31:0] TestBlock__A_op65,
  input wire [31:0] TestBlock__A_op66,
  input wire [31:0] TestBlock__A_op67,
  input wire [31:0] TestBlock__A_op68,
  input wire [31:0] TestBlock__A_op69,
  input wire [31:0] TestBlock__A_op70,
  input wire [31:0] TestBlock__A_op71,
  input wire [31:0] TestBlock__A_op72,
  input wire [31:0] TestBlock__A_op73,
  input wire [31:0] TestBlock__A_op74,
  input wire [31:0] TestBlock__A_op75,
  input wire [31:0] TestBlock__A_op76,
  input wire [31:0] TestBlock__A_op77,
  input wire [31:0] TestBlock__A_op78,
  input wire [31:0] TestBlock__A_op79,
  input wire [31:0] TestBlock__A_op80,
  input wire [31:0] TestBlock__A_op81,
  input wire [31:0] TestBlock__A_op82,
  input wire [31:0] TestBlock__A_op83,
  input wire [31:0] TestBlock__A_op84,
  input wire [31:0] TestBlock__A_op85,
  input wire [31:0] TestBlock__A_op86,
  input wire [31:0] TestBlock__A_op87,
  input wire [31:0] TestBlock__A_op88,
  input wire [31:0] TestBlock__A_op89,
  input wire [31:0] TestBlock__A_op90,
  input wire [31:0] TestBlock__A_op91,
  input wire [31:0] TestBlock__A_op92,
  input wire [31:0] TestBlock__A_op93,
  input wire [31:0] TestBlock__A_op94,
  input wire [31:0] TestBlock__A_op95,
  input wire [31:0] TestBlock__A_op96,
  input wire [31:0] TestBlock__A_op97,
  input wire [31:0] TestBlock__A_op98,
  input wire [31:0] TestBlock__A_op99,
  input wire [31:0] TestBlock__B_op0,
  input wire [31:0] TestBlock__B_op1,
  input wire [31:0] TestBlock__B_op2,
  input wire [31:0] TestBlock__B_op3,
  input wire [31:0] TestBlock__B_op4,
  input wire [31:0] TestBlock__B_op5,
  input wire [31:0] TestBlock__B_op6,
  input wire [31:0] TestBlock__B_op7,
  input wire [31:0] TestBlock__B_op8,
  input wire [31:0] TestBlock__B_op9,
  input wire [31:0] TestBlock__B_op10,
  input wire [31:0] TestBlock__B_op11,
  input wire [31:0] TestBlock__B_op12,
  input wire [31:0] TestBlock__B_op13,
  input wire [31:0] TestBlock__B_op14,
  input wire [31:0] TestBlock__B_op15,
  input wire [31:0] TestBlock__B_op16,
  input wire [31:0] TestBlock__B_op17,
  input wire [31:0] TestBlock__B_op18,
  input wire [31:0] TestBlock__B_op19,
  input wire [31:0] TestBlock__B_op20,
  input wire [31:0] TestBlock__B_op21,
  input wire [31:0] TestBlock__B_op22,
  input wire [31:0] TestBlock__B_op23,
  input wire [31:0] TestBlock__B_op24,
  input wire [31:0] TestBlock__B_op25,
  input wire [31:0] TestBlock__B_op26,
  input wire [31:0] TestBlock__B_op27,
  input wire [31:0] TestBlock__B_op28,
  input wire [31:0] TestBlock__B_op29,
  input wire [31:0] TestBlock__B_op30,
  input wire [31:0] TestBlock__B_op31,
  input wire [31:0] TestBlock__B_op32,
  input wire [31:0] TestBlock__B_op33,
  input wire [31:0] TestBlock__B_op34,
  input wire [31:0] TestBlock__B_op35,
  input wire [31:0] TestBlock__B_op36,
  input wire [31:0] TestBlock__B_op37,
  input wire [31:0] TestBlock__B_op38,
  input wire [31:0] TestBlock__B_op39,
  input wire [31:0] TestBlock__B_op40,
  input wire [31:0] TestBlock__B_op41,
  input wire [31:0] TestBlock__B_op42,
  input wire [31:0] TestBlock__B_op43,
  input wire [31:0] TestBlock__B_op44,
  input wire [31:0] TestBlock__B_op45,
  input wire [31:0] TestBlock__B_op46,
  input wire [31:0] TestBlock__B_op47,
  input wire [31:0] TestBlock__B_op48,
  input wire [31:0] TestBlock__B_op49,
  input wire [31:0] TestBlock__B_op50,
  input wire [31:0] TestBlock__B_op51,
  input wire [31:0] TestBlock__B_op52,
  input wire [31:0] TestBlock__B_op53,
  input wire [31:0] TestBlock__B_op54,
  input wire [31:0] TestBlock__B_op55,
  input wire [31:0] TestBlock__B_op56,
  input wire [31:0] TestBlock__B_op57,
  input wire [31:0] TestBlock__B_op58,
  input wire [31:0] TestBlock__B_op59,
  input wire [31:0] TestBlock__B_op60,
  input wire [31:0] TestBlock__B_op61,
  input wire [31:0] TestBlock__B_op62,
  input wire [31:0] TestBlock__B_op63,
  input wire [31:0] TestBlock__B_op64,
  input wire [31:0] TestBlock__B_op65,
  input wire [31:0] TestBlock__B_op66,
  input wire [31:0] TestBlock__B_op67,
  input wire [31:0] TestBlock__B_op68,
  input wire [31:0] TestBlock__B_op69,
  input wire [31:0] TestBlock__B_op70,
  input wire [31:0] TestBlock__B_op71,
  input wire [31:0] TestBlock__B_op72,
  input wire [31:0] TestBlock__B_op73,
  input wire [31:0] TestBlock__B_op74,
  input wire [31:0] TestBlock__B_op75,
  input wire [31:0] TestBlock__B_op76,
  input wire [31:0] TestBlock__B_op77,
  input wire [31:0] TestBlock__B_op78,
  input wire [31:0] TestBlock__B_op79,
  input wire [31:0] TestBlock__B_op80,
  input wire [31:0] TestBlock__B_op81,
  input wire [31:0] TestBlock__B_op82,
  input wire [31:0] TestBlock__B_op83,
  input wire [31:0] TestBlock__B_op84,
  input wire [31:0] TestBlock__B_op85,
  input wire [31:0] TestBlock__B_op86,
  input wire [31:0] TestBlock__B_op87,
  input wire [31:0] TestBlock__B_op88,
  input wire [31:0] TestBlock__B_op89,
  input wire [31:0] TestBlock__B_op90,
  input wire [31:0] TestBlock__B_op91,
  input wire [31:0] TestBlock__B_op92,
  input wire [31:0] TestBlock__B_op93,
  input wire [31:0] TestBlock__B_op94,
  input wire [31:0] TestBlock__B_op95,
  input wire [31:0] TestBlock__B_op96,
  input wire [31:0] TestBlock__B_op97,
  input wire [31:0] TestBlock__B_op98,
  input wire [31:0] TestBlock__B_op99,
  output wire [3499:0] out
);
  // lint_off SIGNED_TYPE
  // lint_off MULTIPLY
  function automatic [31:0] smul32b_32b_x_32b (input reg [31:0] lhs, input reg [31:0] rhs);
    reg signed [31:0] signed_lhs;
    reg signed [31:0] signed_rhs;
    reg signed [31:0] signed_result;
    begin
      signed_lhs = $signed(lhs);
      signed_rhs = $signed(rhs);
      signed_result = signed_lhs * signed_rhs;
      smul32b_32b_x_32b = $unsigned(signed_result);
    end
  endfunction
  // lint_on MULTIPLY
  // lint_on SIGNED_TYPE

  // ===== Pipe stage 0:

  // Registers for pipe stage 0:
  reg [31:0] p0_TestBlock__A_op0;
  reg [31:0] p0_TestBlock__A_op1;
  reg [31:0] p0_TestBlock__A_op2;
  reg [31:0] p0_TestBlock__A_op3;
  reg [31:0] p0_TestBlock__A_op4;
  reg [31:0] p0_TestBlock__A_op5;
  reg [31:0] p0_TestBlock__A_op6;
  reg [31:0] p0_TestBlock__A_op7;
  reg [31:0] p0_TestBlock__A_op8;
  reg [31:0] p0_TestBlock__A_op9;
  reg [31:0] p0_TestBlock__A_op10;
  reg [31:0] p0_TestBlock__A_op11;
  reg [31:0] p0_TestBlock__A_op12;
  reg [31:0] p0_TestBlock__A_op13;
  reg [31:0] p0_TestBlock__A_op14;
  reg [31:0] p0_TestBlock__A_op15;
  reg [31:0] p0_TestBlock__A_op16;
  reg [31:0] p0_TestBlock__A_op17;
  reg [31:0] p0_TestBlock__A_op18;
  reg [31:0] p0_TestBlock__A_op19;
  reg [31:0] p0_TestBlock__A_op20;
  reg [31:0] p0_TestBlock__A_op21;
  reg [31:0] p0_TestBlock__A_op22;
  reg [31:0] p0_TestBlock__A_op23;
  reg [31:0] p0_TestBlock__A_op24;
  reg [31:0] p0_TestBlock__A_op25;
  reg [31:0] p0_TestBlock__A_op26;
  reg [31:0] p0_TestBlock__A_op27;
  reg [31:0] p0_TestBlock__A_op28;
  reg [31:0] p0_TestBlock__A_op29;
  reg [31:0] p0_TestBlock__A_op30;
  reg [31:0] p0_TestBlock__A_op31;
  reg [31:0] p0_TestBlock__A_op32;
  reg [31:0] p0_TestBlock__A_op33;
  reg [31:0] p0_TestBlock__A_op34;
  reg [31:0] p0_TestBlock__A_op35;
  reg [31:0] p0_TestBlock__A_op36;
  reg [31:0] p0_TestBlock__A_op37;
  reg [31:0] p0_TestBlock__A_op38;
  reg [31:0] p0_TestBlock__A_op39;
  reg [31:0] p0_TestBlock__A_op40;
  reg [31:0] p0_TestBlock__A_op41;
  reg [31:0] p0_TestBlock__A_op42;
  reg [31:0] p0_TestBlock__A_op43;
  reg [31:0] p0_TestBlock__A_op44;
  reg [31:0] p0_TestBlock__A_op45;
  reg [31:0] p0_TestBlock__A_op46;
  reg [31:0] p0_TestBlock__A_op47;
  reg [31:0] p0_TestBlock__A_op48;
  reg [31:0] p0_TestBlock__A_op49;
  reg [31:0] p0_TestBlock__A_op50;
  reg [31:0] p0_TestBlock__A_op51;
  reg [31:0] p0_TestBlock__A_op52;
  reg [31:0] p0_TestBlock__A_op53;
  reg [31:0] p0_TestBlock__A_op54;
  reg [31:0] p0_TestBlock__A_op55;
  reg [31:0] p0_TestBlock__A_op56;
  reg [31:0] p0_TestBlock__A_op57;
  reg [31:0] p0_TestBlock__A_op58;
  reg [31:0] p0_TestBlock__A_op59;
  reg [31:0] p0_TestBlock__A_op60;
  reg [31:0] p0_TestBlock__A_op61;
  reg [31:0] p0_TestBlock__A_op62;
  reg [31:0] p0_TestBlock__A_op63;
  reg [31:0] p0_TestBlock__A_op64;
  reg [31:0] p0_TestBlock__A_op65;
  reg [31:0] p0_TestBlock__A_op66;
  reg [31:0] p0_TestBlock__A_op67;
  reg [31:0] p0_TestBlock__A_op68;
  reg [31:0] p0_TestBlock__A_op69;
  reg [31:0] p0_TestBlock__A_op70;
  reg [31:0] p0_TestBlock__A_op71;
  reg [31:0] p0_TestBlock__A_op72;
  reg [31:0] p0_TestBlock__A_op73;
  reg [31:0] p0_TestBlock__A_op74;
  reg [31:0] p0_TestBlock__A_op75;
  reg [31:0] p0_TestBlock__A_op76;
  reg [31:0] p0_TestBlock__A_op77;
  reg [31:0] p0_TestBlock__A_op78;
  reg [31:0] p0_TestBlock__A_op79;
  reg [31:0] p0_TestBlock__A_op80;
  reg [31:0] p0_TestBlock__A_op81;
  reg [31:0] p0_TestBlock__A_op82;
  reg [31:0] p0_TestBlock__A_op83;
  reg [31:0] p0_TestBlock__A_op84;
  reg [31:0] p0_TestBlock__A_op85;
  reg [31:0] p0_TestBlock__A_op86;
  reg [31:0] p0_TestBlock__A_op87;
  reg [31:0] p0_TestBlock__A_op88;
  reg [31:0] p0_TestBlock__A_op89;
  reg [31:0] p0_TestBlock__A_op90;
  reg [31:0] p0_TestBlock__A_op91;
  reg [31:0] p0_TestBlock__A_op92;
  reg [31:0] p0_TestBlock__A_op93;
  reg [31:0] p0_TestBlock__A_op94;
  reg [31:0] p0_TestBlock__A_op95;
  reg [31:0] p0_TestBlock__A_op96;
  reg [31:0] p0_TestBlock__A_op97;
  reg [31:0] p0_TestBlock__A_op98;
  reg [31:0] p0_TestBlock__A_op99;
  reg [31:0] p0_TestBlock__B_op0;
  reg [31:0] p0_TestBlock__B_op1;
  reg [31:0] p0_TestBlock__B_op2;
  reg [31:0] p0_TestBlock__B_op3;
  reg [31:0] p0_TestBlock__B_op4;
  reg [31:0] p0_TestBlock__B_op5;
  reg [31:0] p0_TestBlock__B_op6;
  reg [31:0] p0_TestBlock__B_op7;
  reg [31:0] p0_TestBlock__B_op8;
  reg [31:0] p0_TestBlock__B_op9;
  reg [31:0] p0_TestBlock__B_op10;
  reg [31:0] p0_TestBlock__B_op11;
  reg [31:0] p0_TestBlock__B_op12;
  reg [31:0] p0_TestBlock__B_op13;
  reg [31:0] p0_TestBlock__B_op14;
  reg [31:0] p0_TestBlock__B_op15;
  reg [31:0] p0_TestBlock__B_op16;
  reg [31:0] p0_TestBlock__B_op17;
  reg [31:0] p0_TestBlock__B_op18;
  reg [31:0] p0_TestBlock__B_op19;
  reg [31:0] p0_TestBlock__B_op20;
  reg [31:0] p0_TestBlock__B_op21;
  reg [31:0] p0_TestBlock__B_op22;
  reg [31:0] p0_TestBlock__B_op23;
  reg [31:0] p0_TestBlock__B_op24;
  reg [31:0] p0_TestBlock__B_op25;
  reg [31:0] p0_TestBlock__B_op26;
  reg [31:0] p0_TestBlock__B_op27;
  reg [31:0] p0_TestBlock__B_op28;
  reg [31:0] p0_TestBlock__B_op29;
  reg [31:0] p0_TestBlock__B_op30;
  reg [31:0] p0_TestBlock__B_op31;
  reg [31:0] p0_TestBlock__B_op32;
  reg [31:0] p0_TestBlock__B_op33;
  reg [31:0] p0_TestBlock__B_op34;
  reg [31:0] p0_TestBlock__B_op35;
  reg [31:0] p0_TestBlock__B_op36;
  reg [31:0] p0_TestBlock__B_op37;
  reg [31:0] p0_TestBlock__B_op38;
  reg [31:0] p0_TestBlock__B_op39;
  reg [31:0] p0_TestBlock__B_op40;
  reg [31:0] p0_TestBlock__B_op41;
  reg [31:0] p0_TestBlock__B_op42;
  reg [31:0] p0_TestBlock__B_op43;
  reg [31:0] p0_TestBlock__B_op44;
  reg [31:0] p0_TestBlock__B_op45;
  reg [31:0] p0_TestBlock__B_op46;
  reg [31:0] p0_TestBlock__B_op47;
  reg [31:0] p0_TestBlock__B_op48;
  reg [31:0] p0_TestBlock__B_op49;
  reg [31:0] p0_TestBlock__B_op50;
  reg [31:0] p0_TestBlock__B_op51;
  reg [31:0] p0_TestBlock__B_op52;
  reg [31:0] p0_TestBlock__B_op53;
  reg [31:0] p0_TestBlock__B_op54;
  reg [31:0] p0_TestBlock__B_op55;
  reg [31:0] p0_TestBlock__B_op56;
  reg [31:0] p0_TestBlock__B_op57;
  reg [31:0] p0_TestBlock__B_op58;
  reg [31:0] p0_TestBlock__B_op59;
  reg [31:0] p0_TestBlock__B_op60;
  reg [31:0] p0_TestBlock__B_op61;
  reg [31:0] p0_TestBlock__B_op62;
  reg [31:0] p0_TestBlock__B_op63;
  reg [31:0] p0_TestBlock__B_op64;
  reg [31:0] p0_TestBlock__B_op65;
  reg [31:0] p0_TestBlock__B_op66;
  reg [31:0] p0_TestBlock__B_op67;
  reg [31:0] p0_TestBlock__B_op68;
  reg [31:0] p0_TestBlock__B_op69;
  reg [31:0] p0_TestBlock__B_op70;
  reg [31:0] p0_TestBlock__B_op71;
  reg [31:0] p0_TestBlock__B_op72;
  reg [31:0] p0_TestBlock__B_op73;
  reg [31:0] p0_TestBlock__B_op74;
  reg [31:0] p0_TestBlock__B_op75;
  reg [31:0] p0_TestBlock__B_op76;
  reg [31:0] p0_TestBlock__B_op77;
  reg [31:0] p0_TestBlock__B_op78;
  reg [31:0] p0_TestBlock__B_op79;
  reg [31:0] p0_TestBlock__B_op80;
  reg [31:0] p0_TestBlock__B_op81;
  reg [31:0] p0_TestBlock__B_op82;
  reg [31:0] p0_TestBlock__B_op83;
  reg [31:0] p0_TestBlock__B_op84;
  reg [31:0] p0_TestBlock__B_op85;
  reg [31:0] p0_TestBlock__B_op86;
  reg [31:0] p0_TestBlock__B_op87;
  reg [31:0] p0_TestBlock__B_op88;
  reg [31:0] p0_TestBlock__B_op89;
  reg [31:0] p0_TestBlock__B_op90;
  reg [31:0] p0_TestBlock__B_op91;
  reg [31:0] p0_TestBlock__B_op92;
  reg [31:0] p0_TestBlock__B_op93;
  reg [31:0] p0_TestBlock__B_op94;
  reg [31:0] p0_TestBlock__B_op95;
  reg [31:0] p0_TestBlock__B_op96;
  reg [31:0] p0_TestBlock__B_op97;
  reg [31:0] p0_TestBlock__B_op98;
  reg [31:0] p0_TestBlock__B_op99;
  always_ff @ (posedge clk) begin
    p0_TestBlock__A_op0 <= TestBlock__A_op0;
    p0_TestBlock__A_op1 <= TestBlock__A_op1;
    p0_TestBlock__A_op2 <= TestBlock__A_op2;
    p0_TestBlock__A_op3 <= TestBlock__A_op3;
    p0_TestBlock__A_op4 <= TestBlock__A_op4;
    p0_TestBlock__A_op5 <= TestBlock__A_op5;
    p0_TestBlock__A_op6 <= TestBlock__A_op6;
    p0_TestBlock__A_op7 <= TestBlock__A_op7;
    p0_TestBlock__A_op8 <= TestBlock__A_op8;
    p0_TestBlock__A_op9 <= TestBlock__A_op9;
    p0_TestBlock__A_op10 <= TestBlock__A_op10;
    p0_TestBlock__A_op11 <= TestBlock__A_op11;
    p0_TestBlock__A_op12 <= TestBlock__A_op12;
    p0_TestBlock__A_op13 <= TestBlock__A_op13;
    p0_TestBlock__A_op14 <= TestBlock__A_op14;
    p0_TestBlock__A_op15 <= TestBlock__A_op15;
    p0_TestBlock__A_op16 <= TestBlock__A_op16;
    p0_TestBlock__A_op17 <= TestBlock__A_op17;
    p0_TestBlock__A_op18 <= TestBlock__A_op18;
    p0_TestBlock__A_op19 <= TestBlock__A_op19;
    p0_TestBlock__A_op20 <= TestBlock__A_op20;
    p0_TestBlock__A_op21 <= TestBlock__A_op21;
    p0_TestBlock__A_op22 <= TestBlock__A_op22;
    p0_TestBlock__A_op23 <= TestBlock__A_op23;
    p0_TestBlock__A_op24 <= TestBlock__A_op24;
    p0_TestBlock__A_op25 <= TestBlock__A_op25;
    p0_TestBlock__A_op26 <= TestBlock__A_op26;
    p0_TestBlock__A_op27 <= TestBlock__A_op27;
    p0_TestBlock__A_op28 <= TestBlock__A_op28;
    p0_TestBlock__A_op29 <= TestBlock__A_op29;
    p0_TestBlock__A_op30 <= TestBlock__A_op30;
    p0_TestBlock__A_op31 <= TestBlock__A_op31;
    p0_TestBlock__A_op32 <= TestBlock__A_op32;
    p0_TestBlock__A_op33 <= TestBlock__A_op33;
    p0_TestBlock__A_op34 <= TestBlock__A_op34;
    p0_TestBlock__A_op35 <= TestBlock__A_op35;
    p0_TestBlock__A_op36 <= TestBlock__A_op36;
    p0_TestBlock__A_op37 <= TestBlock__A_op37;
    p0_TestBlock__A_op38 <= TestBlock__A_op38;
    p0_TestBlock__A_op39 <= TestBlock__A_op39;
    p0_TestBlock__A_op40 <= TestBlock__A_op40;
    p0_TestBlock__A_op41 <= TestBlock__A_op41;
    p0_TestBlock__A_op42 <= TestBlock__A_op42;
    p0_TestBlock__A_op43 <= TestBlock__A_op43;
    p0_TestBlock__A_op44 <= TestBlock__A_op44;
    p0_TestBlock__A_op45 <= TestBlock__A_op45;
    p0_TestBlock__A_op46 <= TestBlock__A_op46;
    p0_TestBlock__A_op47 <= TestBlock__A_op47;
    p0_TestBlock__A_op48 <= TestBlock__A_op48;
    p0_TestBlock__A_op49 <= TestBlock__A_op49;
    p0_TestBlock__A_op50 <= TestBlock__A_op50;
    p0_TestBlock__A_op51 <= TestBlock__A_op51;
    p0_TestBlock__A_op52 <= TestBlock__A_op52;
    p0_TestBlock__A_op53 <= TestBlock__A_op53;
    p0_TestBlock__A_op54 <= TestBlock__A_op54;
    p0_TestBlock__A_op55 <= TestBlock__A_op55;
    p0_TestBlock__A_op56 <= TestBlock__A_op56;
    p0_TestBlock__A_op57 <= TestBlock__A_op57;
    p0_TestBlock__A_op58 <= TestBlock__A_op58;
    p0_TestBlock__A_op59 <= TestBlock__A_op59;
    p0_TestBlock__A_op60 <= TestBlock__A_op60;
    p0_TestBlock__A_op61 <= TestBlock__A_op61;
    p0_TestBlock__A_op62 <= TestBlock__A_op62;
    p0_TestBlock__A_op63 <= TestBlock__A_op63;
    p0_TestBlock__A_op64 <= TestBlock__A_op64;
    p0_TestBlock__A_op65 <= TestBlock__A_op65;
    p0_TestBlock__A_op66 <= TestBlock__A_op66;
    p0_TestBlock__A_op67 <= TestBlock__A_op67;
    p0_TestBlock__A_op68 <= TestBlock__A_op68;
    p0_TestBlock__A_op69 <= TestBlock__A_op69;
    p0_TestBlock__A_op70 <= TestBlock__A_op70;
    p0_TestBlock__A_op71 <= TestBlock__A_op71;
    p0_TestBlock__A_op72 <= TestBlock__A_op72;
    p0_TestBlock__A_op73 <= TestBlock__A_op73;
    p0_TestBlock__A_op74 <= TestBlock__A_op74;
    p0_TestBlock__A_op75 <= TestBlock__A_op75;
    p0_TestBlock__A_op76 <= TestBlock__A_op76;
    p0_TestBlock__A_op77 <= TestBlock__A_op77;
    p0_TestBlock__A_op78 <= TestBlock__A_op78;
    p0_TestBlock__A_op79 <= TestBlock__A_op79;
    p0_TestBlock__A_op80 <= TestBlock__A_op80;
    p0_TestBlock__A_op81 <= TestBlock__A_op81;
    p0_TestBlock__A_op82 <= TestBlock__A_op82;
    p0_TestBlock__A_op83 <= TestBlock__A_op83;
    p0_TestBlock__A_op84 <= TestBlock__A_op84;
    p0_TestBlock__A_op85 <= TestBlock__A_op85;
    p0_TestBlock__A_op86 <= TestBlock__A_op86;
    p0_TestBlock__A_op87 <= TestBlock__A_op87;
    p0_TestBlock__A_op88 <= TestBlock__A_op88;
    p0_TestBlock__A_op89 <= TestBlock__A_op89;
    p0_TestBlock__A_op90 <= TestBlock__A_op90;
    p0_TestBlock__A_op91 <= TestBlock__A_op91;
    p0_TestBlock__A_op92 <= TestBlock__A_op92;
    p0_TestBlock__A_op93 <= TestBlock__A_op93;
    p0_TestBlock__A_op94 <= TestBlock__A_op94;
    p0_TestBlock__A_op95 <= TestBlock__A_op95;
    p0_TestBlock__A_op96 <= TestBlock__A_op96;
    p0_TestBlock__A_op97 <= TestBlock__A_op97;
    p0_TestBlock__A_op98 <= TestBlock__A_op98;
    p0_TestBlock__A_op99 <= TestBlock__A_op99;
    p0_TestBlock__B_op0 <= TestBlock__B_op0;
    p0_TestBlock__B_op1 <= TestBlock__B_op1;
    p0_TestBlock__B_op2 <= TestBlock__B_op2;
    p0_TestBlock__B_op3 <= TestBlock__B_op3;
    p0_TestBlock__B_op4 <= TestBlock__B_op4;
    p0_TestBlock__B_op5 <= TestBlock__B_op5;
    p0_TestBlock__B_op6 <= TestBlock__B_op6;
    p0_TestBlock__B_op7 <= TestBlock__B_op7;
    p0_TestBlock__B_op8 <= TestBlock__B_op8;
    p0_TestBlock__B_op9 <= TestBlock__B_op9;
    p0_TestBlock__B_op10 <= TestBlock__B_op10;
    p0_TestBlock__B_op11 <= TestBlock__B_op11;
    p0_TestBlock__B_op12 <= TestBlock__B_op12;
    p0_TestBlock__B_op13 <= TestBlock__B_op13;
    p0_TestBlock__B_op14 <= TestBlock__B_op14;
    p0_TestBlock__B_op15 <= TestBlock__B_op15;
    p0_TestBlock__B_op16 <= TestBlock__B_op16;
    p0_TestBlock__B_op17 <= TestBlock__B_op17;
    p0_TestBlock__B_op18 <= TestBlock__B_op18;
    p0_TestBlock__B_op19 <= TestBlock__B_op19;
    p0_TestBlock__B_op20 <= TestBlock__B_op20;
    p0_TestBlock__B_op21 <= TestBlock__B_op21;
    p0_TestBlock__B_op22 <= TestBlock__B_op22;
    p0_TestBlock__B_op23 <= TestBlock__B_op23;
    p0_TestBlock__B_op24 <= TestBlock__B_op24;
    p0_TestBlock__B_op25 <= TestBlock__B_op25;
    p0_TestBlock__B_op26 <= TestBlock__B_op26;
    p0_TestBlock__B_op27 <= TestBlock__B_op27;
    p0_TestBlock__B_op28 <= TestBlock__B_op28;
    p0_TestBlock__B_op29 <= TestBlock__B_op29;
    p0_TestBlock__B_op30 <= TestBlock__B_op30;
    p0_TestBlock__B_op31 <= TestBlock__B_op31;
    p0_TestBlock__B_op32 <= TestBlock__B_op32;
    p0_TestBlock__B_op33 <= TestBlock__B_op33;
    p0_TestBlock__B_op34 <= TestBlock__B_op34;
    p0_TestBlock__B_op35 <= TestBlock__B_op35;
    p0_TestBlock__B_op36 <= TestBlock__B_op36;
    p0_TestBlock__B_op37 <= TestBlock__B_op37;
    p0_TestBlock__B_op38 <= TestBlock__B_op38;
    p0_TestBlock__B_op39 <= TestBlock__B_op39;
    p0_TestBlock__B_op40 <= TestBlock__B_op40;
    p0_TestBlock__B_op41 <= TestBlock__B_op41;
    p0_TestBlock__B_op42 <= TestBlock__B_op42;
    p0_TestBlock__B_op43 <= TestBlock__B_op43;
    p0_TestBlock__B_op44 <= TestBlock__B_op44;
    p0_TestBlock__B_op45 <= TestBlock__B_op45;
    p0_TestBlock__B_op46 <= TestBlock__B_op46;
    p0_TestBlock__B_op47 <= TestBlock__B_op47;
    p0_TestBlock__B_op48 <= TestBlock__B_op48;
    p0_TestBlock__B_op49 <= TestBlock__B_op49;
    p0_TestBlock__B_op50 <= TestBlock__B_op50;
    p0_TestBlock__B_op51 <= TestBlock__B_op51;
    p0_TestBlock__B_op52 <= TestBlock__B_op52;
    p0_TestBlock__B_op53 <= TestBlock__B_op53;
    p0_TestBlock__B_op54 <= TestBlock__B_op54;
    p0_TestBlock__B_op55 <= TestBlock__B_op55;
    p0_TestBlock__B_op56 <= TestBlock__B_op56;
    p0_TestBlock__B_op57 <= TestBlock__B_op57;
    p0_TestBlock__B_op58 <= TestBlock__B_op58;
    p0_TestBlock__B_op59 <= TestBlock__B_op59;
    p0_TestBlock__B_op60 <= TestBlock__B_op60;
    p0_TestBlock__B_op61 <= TestBlock__B_op61;
    p0_TestBlock__B_op62 <= TestBlock__B_op62;
    p0_TestBlock__B_op63 <= TestBlock__B_op63;
    p0_TestBlock__B_op64 <= TestBlock__B_op64;
    p0_TestBlock__B_op65 <= TestBlock__B_op65;
    p0_TestBlock__B_op66 <= TestBlock__B_op66;
    p0_TestBlock__B_op67 <= TestBlock__B_op67;
    p0_TestBlock__B_op68 <= TestBlock__B_op68;
    p0_TestBlock__B_op69 <= TestBlock__B_op69;
    p0_TestBlock__B_op70 <= TestBlock__B_op70;
    p0_TestBlock__B_op71 <= TestBlock__B_op71;
    p0_TestBlock__B_op72 <= TestBlock__B_op72;
    p0_TestBlock__B_op73 <= TestBlock__B_op73;
    p0_TestBlock__B_op74 <= TestBlock__B_op74;
    p0_TestBlock__B_op75 <= TestBlock__B_op75;
    p0_TestBlock__B_op76 <= TestBlock__B_op76;
    p0_TestBlock__B_op77 <= TestBlock__B_op77;
    p0_TestBlock__B_op78 <= TestBlock__B_op78;
    p0_TestBlock__B_op79 <= TestBlock__B_op79;
    p0_TestBlock__B_op80 <= TestBlock__B_op80;
    p0_TestBlock__B_op81 <= TestBlock__B_op81;
    p0_TestBlock__B_op82 <= TestBlock__B_op82;
    p0_TestBlock__B_op83 <= TestBlock__B_op83;
    p0_TestBlock__B_op84 <= TestBlock__B_op84;
    p0_TestBlock__B_op85 <= TestBlock__B_op85;
    p0_TestBlock__B_op86 <= TestBlock__B_op86;
    p0_TestBlock__B_op87 <= TestBlock__B_op87;
    p0_TestBlock__B_op88 <= TestBlock__B_op88;
    p0_TestBlock__B_op89 <= TestBlock__B_op89;
    p0_TestBlock__B_op90 <= TestBlock__B_op90;
    p0_TestBlock__B_op91 <= TestBlock__B_op91;
    p0_TestBlock__B_op92 <= TestBlock__B_op92;
    p0_TestBlock__B_op93 <= TestBlock__B_op93;
    p0_TestBlock__B_op94 <= TestBlock__B_op94;
    p0_TestBlock__B_op95 <= TestBlock__B_op95;
    p0_TestBlock__B_op96 <= TestBlock__B_op96;
    p0_TestBlock__B_op97 <= TestBlock__B_op97;
    p0_TestBlock__B_op98 <= TestBlock__B_op98;
    p0_TestBlock__B_op99 <= TestBlock__B_op99;
  end

  // ===== Pipe stage 1:
  wire [31:0] p1_smul_75972_comb;
  wire [31:0] p1_smul_75973_comb;
  wire [31:0] p1_smul_75974_comb;
  wire [31:0] p1_smul_75975_comb;
  wire [31:0] p1_smul_75976_comb;
  wire [31:0] p1_smul_75977_comb;
  wire [31:0] p1_smul_75978_comb;
  wire [31:0] p1_smul_75979_comb;
  wire [31:0] p1_smul_75980_comb;
  wire [31:0] p1_smul_75981_comb;
  wire [31:0] p1_smul_75982_comb;
  wire [31:0] p1_smul_75983_comb;
  wire [31:0] p1_smul_75984_comb;
  wire [31:0] p1_smul_75985_comb;
  wire [31:0] p1_smul_75986_comb;
  wire [31:0] p1_smul_75987_comb;
  wire [31:0] p1_smul_75988_comb;
  wire [31:0] p1_smul_75989_comb;
  wire [31:0] p1_smul_75990_comb;
  wire [31:0] p1_smul_75991_comb;
  wire [31:0] p1_smul_75992_comb;
  wire [31:0] p1_smul_75993_comb;
  wire [31:0] p1_smul_75994_comb;
  wire [31:0] p1_smul_75995_comb;
  wire [31:0] p1_smul_75996_comb;
  wire [31:0] p1_smul_75997_comb;
  wire [31:0] p1_smul_75998_comb;
  wire [31:0] p1_smul_75999_comb;
  wire [31:0] p1_smul_76000_comb;
  wire [31:0] p1_smul_76001_comb;
  wire [31:0] p1_smul_76002_comb;
  wire [31:0] p1_smul_76003_comb;
  wire [31:0] p1_smul_76004_comb;
  wire [31:0] p1_smul_76005_comb;
  wire [31:0] p1_smul_76006_comb;
  wire [31:0] p1_smul_76007_comb;
  wire [31:0] p1_smul_76008_comb;
  wire [31:0] p1_smul_76009_comb;
  wire [31:0] p1_smul_76010_comb;
  wire [31:0] p1_smul_76011_comb;
  wire [31:0] p1_smul_76012_comb;
  wire [31:0] p1_smul_76013_comb;
  wire [31:0] p1_smul_76014_comb;
  wire [31:0] p1_smul_76015_comb;
  wire [31:0] p1_smul_76016_comb;
  wire [31:0] p1_smul_76017_comb;
  wire [31:0] p1_smul_76018_comb;
  wire [31:0] p1_smul_76019_comb;
  wire [31:0] p1_smul_76020_comb;
  wire [31:0] p1_smul_76021_comb;
  wire [31:0] p1_smul_76022_comb;
  wire [31:0] p1_smul_76023_comb;
  wire [31:0] p1_smul_76024_comb;
  wire [31:0] p1_smul_76025_comb;
  wire [31:0] p1_smul_76026_comb;
  wire [31:0] p1_smul_76027_comb;
  wire [31:0] p1_smul_76028_comb;
  wire [31:0] p1_smul_76029_comb;
  wire [31:0] p1_smul_76030_comb;
  wire [31:0] p1_smul_76031_comb;
  wire [31:0] p1_smul_76032_comb;
  wire [31:0] p1_smul_76033_comb;
  wire [31:0] p1_smul_76034_comb;
  wire [31:0] p1_smul_76035_comb;
  wire [31:0] p1_smul_76036_comb;
  wire [31:0] p1_smul_76037_comb;
  wire [31:0] p1_smul_76038_comb;
  wire [31:0] p1_smul_76039_comb;
  wire [31:0] p1_smul_76040_comb;
  wire [31:0] p1_smul_76041_comb;
  wire [31:0] p1_smul_76042_comb;
  wire [31:0] p1_smul_76043_comb;
  wire [31:0] p1_smul_76044_comb;
  wire [31:0] p1_smul_76045_comb;
  wire [31:0] p1_smul_76046_comb;
  wire [31:0] p1_smul_76047_comb;
  wire [31:0] p1_smul_76048_comb;
  wire [31:0] p1_smul_76049_comb;
  wire [31:0] p1_smul_76050_comb;
  wire [31:0] p1_smul_76051_comb;
  wire [31:0] p1_smul_76052_comb;
  wire [31:0] p1_smul_76053_comb;
  wire [31:0] p1_smul_76054_comb;
  wire [31:0] p1_smul_76055_comb;
  wire [31:0] p1_smul_76056_comb;
  wire [31:0] p1_smul_76057_comb;
  wire [31:0] p1_smul_76058_comb;
  wire [31:0] p1_smul_76059_comb;
  wire [31:0] p1_smul_76060_comb;
  wire [31:0] p1_smul_76061_comb;
  wire [31:0] p1_smul_76062_comb;
  wire [31:0] p1_smul_76063_comb;
  wire [31:0] p1_smul_76064_comb;
  wire [31:0] p1_smul_76065_comb;
  wire [31:0] p1_smul_76066_comb;
  wire [31:0] p1_smul_76067_comb;
  wire [31:0] p1_smul_76068_comb;
  wire [31:0] p1_smul_76069_comb;
  wire [31:0] p1_smul_76070_comb;
  wire [31:0] p1_smul_76071_comb;
  wire [31:0] p1_smul_76072_comb;
  wire [31:0] p1_smul_76073_comb;
  wire [31:0] p1_smul_76074_comb;
  wire [31:0] p1_smul_76075_comb;
  wire [31:0] p1_smul_76076_comb;
  wire [31:0] p1_smul_76077_comb;
  wire [31:0] p1_smul_76078_comb;
  wire [31:0] p1_smul_76079_comb;
  wire [31:0] p1_smul_76080_comb;
  wire [31:0] p1_smul_76081_comb;
  wire [31:0] p1_smul_76082_comb;
  wire [31:0] p1_smul_76083_comb;
  wire [31:0] p1_smul_76084_comb;
  wire [31:0] p1_smul_76085_comb;
  wire [31:0] p1_smul_76086_comb;
  wire [31:0] p1_smul_76087_comb;
  wire [31:0] p1_smul_76088_comb;
  wire [31:0] p1_smul_76089_comb;
  wire [31:0] p1_smul_76090_comb;
  wire [31:0] p1_smul_76091_comb;
  wire [31:0] p1_smul_76092_comb;
  wire [31:0] p1_smul_76093_comb;
  wire [31:0] p1_smul_76094_comb;
  wire [31:0] p1_smul_76095_comb;
  wire [31:0] p1_smul_76096_comb;
  wire [31:0] p1_smul_76097_comb;
  wire [31:0] p1_smul_76098_comb;
  wire [31:0] p1_smul_76099_comb;
  wire [31:0] p1_smul_76100_comb;
  wire [31:0] p1_smul_76101_comb;
  wire [31:0] p1_smul_76102_comb;
  wire [31:0] p1_smul_76103_comb;
  wire [31:0] p1_smul_76104_comb;
  wire [31:0] p1_smul_76105_comb;
  wire [31:0] p1_smul_76106_comb;
  wire [31:0] p1_smul_76107_comb;
  wire [31:0] p1_smul_76108_comb;
  wire [31:0] p1_smul_76109_comb;
  wire [31:0] p1_smul_76110_comb;
  wire [31:0] p1_smul_76111_comb;
  wire [31:0] p1_smul_76112_comb;
  wire [31:0] p1_smul_76113_comb;
  wire [31:0] p1_smul_76114_comb;
  wire [31:0] p1_smul_76115_comb;
  wire [31:0] p1_smul_76116_comb;
  wire [31:0] p1_smul_76117_comb;
  wire [31:0] p1_smul_76118_comb;
  wire [31:0] p1_smul_76119_comb;
  wire [31:0] p1_smul_76120_comb;
  wire [31:0] p1_smul_76121_comb;
  wire [31:0] p1_smul_76122_comb;
  wire [31:0] p1_smul_76123_comb;
  wire [31:0] p1_smul_76124_comb;
  wire [31:0] p1_smul_76125_comb;
  wire [31:0] p1_smul_76126_comb;
  wire [31:0] p1_smul_76127_comb;
  wire [31:0] p1_smul_76128_comb;
  wire [31:0] p1_smul_76129_comb;
  wire [31:0] p1_smul_76130_comb;
  wire [31:0] p1_smul_76131_comb;
  wire [31:0] p1_smul_76132_comb;
  wire [31:0] p1_smul_76133_comb;
  wire [31:0] p1_smul_76134_comb;
  wire [31:0] p1_smul_76135_comb;
  wire [31:0] p1_smul_76136_comb;
  wire [31:0] p1_smul_76137_comb;
  wire [31:0] p1_smul_76138_comb;
  wire [31:0] p1_smul_76139_comb;
  wire [31:0] p1_smul_76140_comb;
  wire [31:0] p1_smul_76141_comb;
  wire [31:0] p1_smul_76142_comb;
  wire [31:0] p1_smul_76143_comb;
  wire [31:0] p1_smul_76144_comb;
  wire [31:0] p1_smul_76145_comb;
  wire [31:0] p1_smul_76146_comb;
  wire [31:0] p1_smul_76147_comb;
  wire [31:0] p1_smul_76148_comb;
  wire [31:0] p1_smul_76149_comb;
  wire [31:0] p1_smul_76150_comb;
  wire [31:0] p1_smul_76151_comb;
  wire [31:0] p1_smul_76152_comb;
  wire [31:0] p1_smul_76153_comb;
  wire [31:0] p1_smul_76154_comb;
  wire [31:0] p1_smul_76155_comb;
  wire [31:0] p1_smul_76156_comb;
  wire [31:0] p1_smul_76157_comb;
  wire [31:0] p1_smul_76158_comb;
  wire [31:0] p1_smul_76159_comb;
  wire [31:0] p1_smul_76160_comb;
  wire [31:0] p1_smul_76161_comb;
  wire [31:0] p1_smul_76162_comb;
  wire [31:0] p1_smul_76163_comb;
  wire [31:0] p1_smul_76164_comb;
  wire [31:0] p1_smul_76165_comb;
  wire [31:0] p1_smul_76166_comb;
  wire [31:0] p1_smul_76167_comb;
  wire [31:0] p1_smul_76168_comb;
  wire [31:0] p1_smul_76169_comb;
  wire [31:0] p1_smul_76170_comb;
  wire [31:0] p1_smul_76171_comb;
  wire [31:0] p1_smul_76172_comb;
  wire [31:0] p1_smul_76173_comb;
  wire [31:0] p1_smul_76174_comb;
  wire [31:0] p1_smul_76175_comb;
  wire [31:0] p1_smul_76176_comb;
  wire [31:0] p1_smul_76177_comb;
  wire [31:0] p1_smul_76178_comb;
  wire [31:0] p1_smul_76179_comb;
  wire [31:0] p1_smul_76180_comb;
  wire [31:0] p1_smul_76181_comb;
  wire [31:0] p1_smul_76182_comb;
  wire [31:0] p1_smul_76183_comb;
  wire [31:0] p1_smul_76184_comb;
  wire [31:0] p1_smul_76185_comb;
  wire [31:0] p1_smul_76186_comb;
  wire [31:0] p1_smul_76187_comb;
  wire [31:0] p1_smul_76188_comb;
  wire [31:0] p1_smul_76189_comb;
  wire [31:0] p1_smul_76190_comb;
  wire [31:0] p1_smul_76191_comb;
  wire [31:0] p1_smul_76192_comb;
  wire [31:0] p1_smul_76193_comb;
  wire [31:0] p1_smul_76194_comb;
  wire [31:0] p1_smul_76195_comb;
  wire [31:0] p1_smul_76196_comb;
  wire [31:0] p1_smul_76197_comb;
  wire [31:0] p1_smul_76198_comb;
  wire [31:0] p1_smul_76199_comb;
  wire [31:0] p1_smul_76200_comb;
  wire [31:0] p1_smul_76201_comb;
  wire [31:0] p1_smul_76202_comb;
  wire [31:0] p1_smul_76203_comb;
  wire [31:0] p1_smul_76204_comb;
  wire [31:0] p1_smul_76205_comb;
  wire [31:0] p1_smul_76206_comb;
  wire [31:0] p1_smul_76207_comb;
  wire [31:0] p1_smul_76208_comb;
  wire [31:0] p1_smul_76209_comb;
  wire [31:0] p1_smul_76210_comb;
  wire [31:0] p1_smul_76211_comb;
  wire [31:0] p1_smul_76212_comb;
  wire [31:0] p1_smul_76213_comb;
  wire [31:0] p1_smul_76214_comb;
  wire [31:0] p1_smul_76215_comb;
  wire [31:0] p1_smul_76216_comb;
  wire [31:0] p1_smul_76217_comb;
  wire [31:0] p1_smul_76218_comb;
  wire [31:0] p1_smul_76219_comb;
  wire [31:0] p1_smul_76220_comb;
  wire [31:0] p1_smul_76221_comb;
  wire [31:0] p1_smul_76222_comb;
  wire [31:0] p1_smul_76223_comb;
  wire [31:0] p1_smul_76224_comb;
  wire [31:0] p1_smul_76225_comb;
  wire [31:0] p1_smul_76226_comb;
  wire [31:0] p1_smul_76227_comb;
  wire [31:0] p1_smul_76228_comb;
  wire [31:0] p1_smul_76229_comb;
  wire [31:0] p1_smul_76230_comb;
  wire [31:0] p1_smul_76231_comb;
  wire [31:0] p1_smul_76232_comb;
  wire [31:0] p1_smul_76233_comb;
  wire [31:0] p1_smul_76234_comb;
  wire [31:0] p1_smul_76235_comb;
  wire [31:0] p1_smul_76236_comb;
  wire [31:0] p1_smul_76237_comb;
  wire [31:0] p1_smul_76238_comb;
  wire [31:0] p1_smul_76239_comb;
  wire [31:0] p1_smul_76240_comb;
  wire [31:0] p1_smul_76241_comb;
  wire [31:0] p1_smul_76242_comb;
  wire [31:0] p1_smul_76243_comb;
  wire [31:0] p1_smul_76244_comb;
  wire [31:0] p1_smul_76245_comb;
  wire [31:0] p1_smul_76246_comb;
  wire [31:0] p1_smul_76247_comb;
  wire [31:0] p1_smul_76248_comb;
  wire [31:0] p1_smul_76249_comb;
  wire [31:0] p1_smul_76250_comb;
  wire [31:0] p1_smul_76251_comb;
  wire [31:0] p1_smul_76252_comb;
  wire [31:0] p1_smul_76253_comb;
  wire [31:0] p1_smul_76254_comb;
  wire [31:0] p1_smul_76255_comb;
  wire [31:0] p1_smul_76256_comb;
  wire [31:0] p1_smul_76257_comb;
  wire [31:0] p1_smul_76258_comb;
  wire [31:0] p1_smul_76259_comb;
  wire [31:0] p1_smul_76260_comb;
  wire [31:0] p1_smul_76261_comb;
  wire [31:0] p1_smul_76262_comb;
  wire [31:0] p1_smul_76263_comb;
  wire [31:0] p1_smul_76264_comb;
  wire [31:0] p1_smul_76265_comb;
  wire [31:0] p1_smul_76266_comb;
  wire [31:0] p1_smul_76267_comb;
  wire [31:0] p1_smul_76268_comb;
  wire [31:0] p1_smul_76269_comb;
  wire [31:0] p1_smul_76270_comb;
  wire [31:0] p1_smul_76271_comb;
  wire [31:0] p1_smul_76272_comb;
  wire [31:0] p1_smul_76273_comb;
  wire [31:0] p1_smul_76274_comb;
  wire [31:0] p1_smul_76275_comb;
  wire [31:0] p1_smul_76276_comb;
  wire [31:0] p1_smul_76277_comb;
  wire [31:0] p1_smul_76278_comb;
  wire [31:0] p1_smul_76279_comb;
  wire [31:0] p1_smul_76280_comb;
  wire [31:0] p1_smul_76281_comb;
  wire [31:0] p1_smul_76282_comb;
  wire [31:0] p1_smul_76283_comb;
  wire [31:0] p1_smul_76284_comb;
  wire [31:0] p1_smul_76285_comb;
  wire [31:0] p1_smul_76286_comb;
  wire [31:0] p1_smul_76287_comb;
  wire [31:0] p1_smul_76288_comb;
  wire [31:0] p1_smul_76289_comb;
  wire [31:0] p1_smul_76290_comb;
  wire [31:0] p1_smul_76291_comb;
  wire [31:0] p1_smul_76292_comb;
  wire [31:0] p1_smul_76293_comb;
  wire [31:0] p1_smul_76294_comb;
  wire [31:0] p1_smul_76295_comb;
  wire [31:0] p1_smul_76296_comb;
  wire [31:0] p1_smul_76297_comb;
  wire [31:0] p1_smul_76298_comb;
  wire [31:0] p1_smul_76299_comb;
  wire [31:0] p1_smul_76300_comb;
  wire [31:0] p1_smul_76301_comb;
  wire [31:0] p1_smul_76302_comb;
  wire [31:0] p1_smul_76303_comb;
  wire [31:0] p1_smul_76304_comb;
  wire [31:0] p1_smul_76305_comb;
  wire [31:0] p1_smul_76306_comb;
  wire [31:0] p1_smul_76307_comb;
  wire [31:0] p1_smul_76308_comb;
  wire [31:0] p1_smul_76309_comb;
  wire [31:0] p1_smul_76310_comb;
  wire [31:0] p1_smul_76311_comb;
  wire [31:0] p1_smul_76312_comb;
  wire [31:0] p1_smul_76313_comb;
  wire [31:0] p1_smul_76314_comb;
  wire [31:0] p1_smul_76315_comb;
  wire [31:0] p1_smul_76316_comb;
  wire [31:0] p1_smul_76317_comb;
  wire [31:0] p1_smul_76318_comb;
  wire [31:0] p1_smul_76319_comb;
  wire [31:0] p1_smul_76320_comb;
  wire [31:0] p1_smul_76321_comb;
  wire [31:0] p1_smul_76322_comb;
  wire [31:0] p1_smul_76323_comb;
  wire [31:0] p1_smul_76324_comb;
  wire [31:0] p1_smul_76325_comb;
  wire [31:0] p1_smul_76326_comb;
  wire [31:0] p1_smul_76327_comb;
  wire [31:0] p1_smul_76328_comb;
  wire [31:0] p1_smul_76329_comb;
  wire [31:0] p1_smul_76330_comb;
  wire [31:0] p1_smul_76331_comb;
  wire [31:0] p1_smul_76332_comb;
  wire [31:0] p1_smul_76333_comb;
  wire [31:0] p1_smul_76334_comb;
  wire [31:0] p1_smul_76335_comb;
  wire [31:0] p1_smul_76336_comb;
  wire [31:0] p1_smul_76337_comb;
  wire [31:0] p1_smul_76338_comb;
  wire [31:0] p1_smul_76339_comb;
  wire [31:0] p1_smul_76340_comb;
  wire [31:0] p1_smul_76341_comb;
  wire [31:0] p1_smul_76342_comb;
  wire [31:0] p1_smul_76343_comb;
  wire [31:0] p1_smul_76344_comb;
  wire [31:0] p1_smul_76345_comb;
  wire [31:0] p1_smul_76346_comb;
  wire [31:0] p1_smul_76347_comb;
  wire [31:0] p1_smul_76348_comb;
  wire [31:0] p1_smul_76349_comb;
  wire [31:0] p1_smul_76350_comb;
  wire [31:0] p1_smul_76351_comb;
  wire [31:0] p1_smul_76352_comb;
  wire [31:0] p1_smul_76353_comb;
  wire [31:0] p1_smul_76354_comb;
  wire [31:0] p1_smul_76355_comb;
  wire [31:0] p1_smul_76356_comb;
  wire [31:0] p1_smul_76357_comb;
  wire [31:0] p1_smul_76358_comb;
  wire [31:0] p1_smul_76359_comb;
  wire [31:0] p1_smul_76360_comb;
  wire [31:0] p1_smul_76361_comb;
  wire [31:0] p1_smul_76362_comb;
  wire [31:0] p1_smul_76363_comb;
  wire [31:0] p1_smul_76364_comb;
  wire [31:0] p1_smul_76365_comb;
  wire [31:0] p1_smul_76366_comb;
  wire [31:0] p1_smul_76367_comb;
  wire [31:0] p1_smul_76368_comb;
  wire [31:0] p1_smul_76369_comb;
  wire [31:0] p1_smul_76370_comb;
  wire [31:0] p1_smul_76371_comb;
  wire [31:0] p1_smul_76372_comb;
  wire [31:0] p1_smul_76373_comb;
  wire [31:0] p1_smul_76374_comb;
  wire [31:0] p1_smul_76375_comb;
  wire [31:0] p1_smul_76376_comb;
  wire [31:0] p1_smul_76377_comb;
  wire [31:0] p1_smul_76378_comb;
  wire [31:0] p1_smul_76379_comb;
  wire [31:0] p1_smul_76380_comb;
  wire [31:0] p1_smul_76381_comb;
  wire [31:0] p1_smul_76382_comb;
  wire [31:0] p1_smul_76383_comb;
  wire [31:0] p1_smul_76384_comb;
  wire [31:0] p1_smul_76385_comb;
  wire [31:0] p1_smul_76386_comb;
  wire [31:0] p1_smul_76387_comb;
  wire [31:0] p1_smul_76388_comb;
  wire [31:0] p1_smul_76389_comb;
  wire [31:0] p1_smul_76390_comb;
  wire [31:0] p1_smul_76391_comb;
  wire [31:0] p1_smul_76392_comb;
  wire [31:0] p1_smul_76393_comb;
  wire [31:0] p1_smul_76394_comb;
  wire [31:0] p1_smul_76395_comb;
  wire [31:0] p1_smul_76396_comb;
  wire [31:0] p1_smul_76397_comb;
  wire [31:0] p1_smul_76398_comb;
  wire [31:0] p1_smul_76399_comb;
  wire [31:0] p1_smul_76400_comb;
  wire [31:0] p1_smul_76401_comb;
  wire [31:0] p1_smul_76402_comb;
  wire [31:0] p1_smul_76403_comb;
  wire [31:0] p1_smul_76404_comb;
  wire [31:0] p1_smul_76405_comb;
  wire [31:0] p1_smul_76406_comb;
  wire [31:0] p1_smul_76407_comb;
  wire [31:0] p1_smul_76408_comb;
  wire [31:0] p1_smul_76409_comb;
  wire [31:0] p1_smul_76410_comb;
  wire [31:0] p1_smul_76411_comb;
  wire [31:0] p1_smul_76412_comb;
  wire [31:0] p1_smul_76413_comb;
  wire [31:0] p1_smul_76414_comb;
  wire [31:0] p1_smul_76415_comb;
  wire [31:0] p1_smul_76416_comb;
  wire [31:0] p1_smul_76417_comb;
  wire [31:0] p1_smul_76418_comb;
  wire [31:0] p1_smul_76419_comb;
  wire [31:0] p1_smul_76420_comb;
  wire [31:0] p1_smul_76421_comb;
  wire [31:0] p1_smul_76422_comb;
  wire [31:0] p1_smul_76423_comb;
  wire [31:0] p1_smul_76424_comb;
  wire [31:0] p1_smul_76425_comb;
  wire [31:0] p1_smul_76426_comb;
  wire [31:0] p1_smul_76427_comb;
  wire [31:0] p1_smul_76428_comb;
  wire [31:0] p1_smul_76429_comb;
  wire [31:0] p1_smul_76430_comb;
  wire [31:0] p1_smul_76431_comb;
  wire [31:0] p1_smul_76432_comb;
  wire [31:0] p1_smul_76433_comb;
  wire [31:0] p1_smul_76434_comb;
  wire [31:0] p1_smul_76435_comb;
  wire [31:0] p1_smul_76436_comb;
  wire [31:0] p1_smul_76437_comb;
  wire [31:0] p1_smul_76438_comb;
  wire [31:0] p1_smul_76439_comb;
  wire [31:0] p1_smul_76440_comb;
  wire [31:0] p1_smul_76441_comb;
  wire [31:0] p1_smul_76442_comb;
  wire [31:0] p1_smul_76443_comb;
  wire [31:0] p1_smul_76444_comb;
  wire [31:0] p1_smul_76445_comb;
  wire [31:0] p1_smul_76446_comb;
  wire [31:0] p1_smul_76447_comb;
  wire [31:0] p1_smul_76448_comb;
  wire [31:0] p1_smul_76449_comb;
  wire [31:0] p1_smul_76450_comb;
  wire [31:0] p1_smul_76451_comb;
  wire [31:0] p1_smul_76452_comb;
  wire [31:0] p1_smul_76453_comb;
  wire [31:0] p1_smul_76454_comb;
  wire [31:0] p1_smul_76455_comb;
  wire [31:0] p1_smul_76456_comb;
  wire [31:0] p1_smul_76457_comb;
  wire [31:0] p1_smul_76458_comb;
  wire [31:0] p1_smul_76459_comb;
  wire [31:0] p1_smul_76460_comb;
  wire [31:0] p1_smul_76461_comb;
  wire [31:0] p1_smul_76462_comb;
  wire [31:0] p1_smul_76463_comb;
  wire [31:0] p1_smul_76464_comb;
  wire [31:0] p1_smul_76465_comb;
  wire [31:0] p1_smul_76466_comb;
  wire [31:0] p1_smul_76467_comb;
  wire [31:0] p1_smul_76468_comb;
  wire [31:0] p1_smul_76469_comb;
  wire [31:0] p1_smul_76470_comb;
  wire [31:0] p1_smul_76471_comb;
  wire [31:0] p1_smul_76472_comb;
  wire [31:0] p1_smul_76473_comb;
  wire [31:0] p1_smul_76474_comb;
  wire [31:0] p1_smul_76475_comb;
  wire [31:0] p1_smul_76476_comb;
  wire [31:0] p1_smul_76477_comb;
  wire [31:0] p1_smul_76478_comb;
  wire [31:0] p1_smul_76479_comb;
  wire [31:0] p1_smul_76480_comb;
  wire [31:0] p1_smul_76481_comb;
  wire [31:0] p1_smul_76482_comb;
  wire [31:0] p1_smul_76483_comb;
  wire [31:0] p1_smul_76484_comb;
  wire [31:0] p1_smul_76485_comb;
  wire [31:0] p1_smul_76486_comb;
  wire [31:0] p1_smul_76487_comb;
  wire [31:0] p1_smul_76488_comb;
  wire [31:0] p1_smul_76489_comb;
  wire [31:0] p1_smul_76490_comb;
  wire [31:0] p1_smul_76491_comb;
  wire [31:0] p1_smul_76492_comb;
  wire [31:0] p1_smul_76493_comb;
  wire [31:0] p1_smul_76494_comb;
  wire [31:0] p1_smul_76495_comb;
  wire [31:0] p1_smul_76496_comb;
  wire [31:0] p1_smul_76497_comb;
  wire [31:0] p1_smul_76498_comb;
  wire [31:0] p1_smul_76499_comb;
  wire [31:0] p1_smul_76500_comb;
  wire [31:0] p1_smul_76501_comb;
  wire [31:0] p1_smul_76502_comb;
  wire [31:0] p1_smul_76503_comb;
  wire [31:0] p1_smul_76504_comb;
  wire [31:0] p1_smul_76505_comb;
  wire [31:0] p1_smul_76506_comb;
  wire [31:0] p1_smul_76507_comb;
  wire [31:0] p1_smul_76508_comb;
  wire [31:0] p1_smul_76509_comb;
  wire [31:0] p1_smul_76510_comb;
  wire [31:0] p1_smul_76511_comb;
  wire [31:0] p1_smul_76512_comb;
  wire [31:0] p1_smul_76513_comb;
  wire [31:0] p1_smul_76514_comb;
  wire [31:0] p1_smul_76515_comb;
  wire [31:0] p1_smul_76516_comb;
  wire [31:0] p1_smul_76517_comb;
  wire [31:0] p1_smul_76518_comb;
  wire [31:0] p1_smul_76519_comb;
  wire [31:0] p1_smul_76520_comb;
  wire [31:0] p1_smul_76521_comb;
  wire [31:0] p1_smul_76522_comb;
  wire [31:0] p1_smul_76523_comb;
  wire [31:0] p1_smul_76524_comb;
  wire [31:0] p1_smul_76525_comb;
  wire [31:0] p1_smul_76526_comb;
  wire [31:0] p1_smul_76527_comb;
  wire [31:0] p1_smul_76528_comb;
  wire [31:0] p1_smul_76529_comb;
  wire [31:0] p1_smul_76530_comb;
  wire [31:0] p1_smul_76531_comb;
  wire [31:0] p1_smul_76532_comb;
  wire [31:0] p1_smul_76533_comb;
  wire [31:0] p1_smul_76534_comb;
  wire [31:0] p1_smul_76535_comb;
  wire [31:0] p1_smul_76536_comb;
  wire [31:0] p1_smul_76537_comb;
  wire [31:0] p1_smul_76538_comb;
  wire [31:0] p1_smul_76539_comb;
  wire [31:0] p1_smul_76540_comb;
  wire [31:0] p1_smul_76541_comb;
  wire [31:0] p1_smul_76542_comb;
  wire [31:0] p1_smul_76543_comb;
  wire [31:0] p1_smul_76544_comb;
  wire [31:0] p1_smul_76545_comb;
  wire [31:0] p1_smul_76546_comb;
  wire [31:0] p1_smul_76547_comb;
  wire [31:0] p1_smul_76548_comb;
  wire [31:0] p1_smul_76549_comb;
  wire [31:0] p1_smul_76550_comb;
  wire [31:0] p1_smul_76551_comb;
  wire [31:0] p1_smul_76552_comb;
  wire [31:0] p1_smul_76553_comb;
  wire [31:0] p1_smul_76554_comb;
  wire [31:0] p1_smul_76555_comb;
  wire [31:0] p1_smul_76556_comb;
  wire [31:0] p1_smul_76557_comb;
  wire [31:0] p1_smul_76558_comb;
  wire [31:0] p1_smul_76559_comb;
  wire [31:0] p1_smul_76560_comb;
  wire [31:0] p1_smul_76561_comb;
  wire [31:0] p1_smul_76562_comb;
  wire [31:0] p1_smul_76563_comb;
  wire [31:0] p1_smul_76564_comb;
  wire [31:0] p1_smul_76565_comb;
  wire [31:0] p1_smul_76566_comb;
  wire [31:0] p1_smul_76567_comb;
  wire [31:0] p1_smul_76568_comb;
  wire [31:0] p1_smul_76569_comb;
  wire [31:0] p1_smul_76570_comb;
  wire [31:0] p1_smul_76571_comb;
  wire [31:0] p1_smul_76572_comb;
  wire [31:0] p1_smul_76573_comb;
  wire [31:0] p1_smul_76574_comb;
  wire [31:0] p1_smul_76575_comb;
  wire [31:0] p1_smul_76576_comb;
  wire [31:0] p1_smul_76577_comb;
  wire [31:0] p1_smul_76578_comb;
  wire [31:0] p1_smul_76579_comb;
  wire [31:0] p1_smul_76580_comb;
  wire [31:0] p1_smul_76581_comb;
  wire [31:0] p1_smul_76582_comb;
  wire [31:0] p1_smul_76583_comb;
  wire [31:0] p1_smul_76584_comb;
  wire [31:0] p1_smul_76585_comb;
  wire [31:0] p1_smul_76586_comb;
  wire [31:0] p1_smul_76587_comb;
  wire [31:0] p1_smul_76588_comb;
  wire [31:0] p1_smul_76589_comb;
  wire [31:0] p1_smul_76590_comb;
  wire [31:0] p1_smul_76591_comb;
  wire [31:0] p1_smul_76592_comb;
  wire [31:0] p1_smul_76593_comb;
  wire [31:0] p1_smul_76594_comb;
  wire [31:0] p1_smul_76595_comb;
  wire [31:0] p1_smul_76596_comb;
  wire [31:0] p1_smul_76597_comb;
  wire [31:0] p1_smul_76598_comb;
  wire [31:0] p1_smul_76599_comb;
  wire [31:0] p1_smul_76600_comb;
  wire [31:0] p1_smul_76601_comb;
  wire [31:0] p1_smul_76602_comb;
  wire [31:0] p1_smul_76603_comb;
  wire [31:0] p1_smul_76604_comb;
  wire [31:0] p1_smul_76605_comb;
  wire [31:0] p1_smul_76606_comb;
  wire [31:0] p1_smul_76607_comb;
  wire [31:0] p1_smul_76608_comb;
  wire [31:0] p1_smul_76609_comb;
  wire [31:0] p1_smul_76610_comb;
  wire [31:0] p1_smul_76611_comb;
  wire [31:0] p1_smul_76612_comb;
  wire [31:0] p1_smul_76613_comb;
  wire [31:0] p1_smul_76614_comb;
  wire [31:0] p1_smul_76615_comb;
  wire [31:0] p1_smul_76616_comb;
  wire [31:0] p1_smul_76617_comb;
  wire [31:0] p1_smul_76618_comb;
  wire [31:0] p1_smul_76619_comb;
  wire [31:0] p1_smul_76620_comb;
  wire [31:0] p1_smul_76621_comb;
  wire [31:0] p1_smul_76622_comb;
  wire [31:0] p1_smul_76623_comb;
  wire [31:0] p1_smul_76624_comb;
  wire [31:0] p1_smul_76625_comb;
  wire [31:0] p1_smul_76626_comb;
  wire [31:0] p1_smul_76627_comb;
  wire [31:0] p1_smul_76628_comb;
  wire [31:0] p1_smul_76629_comb;
  wire [31:0] p1_smul_76630_comb;
  wire [31:0] p1_smul_76631_comb;
  wire [31:0] p1_smul_76632_comb;
  wire [31:0] p1_smul_76633_comb;
  wire [31:0] p1_smul_76634_comb;
  wire [31:0] p1_smul_76635_comb;
  wire [31:0] p1_smul_76636_comb;
  wire [31:0] p1_smul_76637_comb;
  wire [31:0] p1_smul_76638_comb;
  wire [31:0] p1_smul_76639_comb;
  wire [31:0] p1_smul_76640_comb;
  wire [31:0] p1_smul_76641_comb;
  wire [31:0] p1_smul_76642_comb;
  wire [31:0] p1_smul_76643_comb;
  wire [31:0] p1_smul_76644_comb;
  wire [31:0] p1_smul_76645_comb;
  wire [31:0] p1_smul_76646_comb;
  wire [31:0] p1_smul_76647_comb;
  wire [31:0] p1_smul_76648_comb;
  wire [31:0] p1_smul_76649_comb;
  wire [31:0] p1_smul_76650_comb;
  wire [31:0] p1_smul_76651_comb;
  wire [31:0] p1_smul_76652_comb;
  wire [31:0] p1_smul_76653_comb;
  wire [31:0] p1_smul_76654_comb;
  wire [31:0] p1_smul_76655_comb;
  wire [31:0] p1_smul_76656_comb;
  wire [31:0] p1_smul_76657_comb;
  wire [31:0] p1_smul_76658_comb;
  wire [31:0] p1_smul_76659_comb;
  wire [31:0] p1_smul_76660_comb;
  wire [31:0] p1_smul_76661_comb;
  wire [31:0] p1_smul_76662_comb;
  wire [31:0] p1_smul_76663_comb;
  wire [31:0] p1_smul_76664_comb;
  wire [31:0] p1_smul_76665_comb;
  wire [31:0] p1_smul_76666_comb;
  wire [31:0] p1_smul_76667_comb;
  wire [31:0] p1_smul_76668_comb;
  wire [31:0] p1_smul_76669_comb;
  wire [31:0] p1_smul_76670_comb;
  wire [31:0] p1_smul_76671_comb;
  wire [31:0] p1_smul_76672_comb;
  wire [31:0] p1_smul_76673_comb;
  wire [31:0] p1_smul_76674_comb;
  wire [31:0] p1_smul_76675_comb;
  wire [31:0] p1_smul_76676_comb;
  wire [31:0] p1_smul_76677_comb;
  wire [31:0] p1_smul_76678_comb;
  wire [31:0] p1_smul_76679_comb;
  wire [31:0] p1_smul_76680_comb;
  wire [31:0] p1_smul_76681_comb;
  wire [31:0] p1_smul_76682_comb;
  wire [31:0] p1_smul_76683_comb;
  wire [31:0] p1_smul_76684_comb;
  wire [31:0] p1_smul_76685_comb;
  wire [31:0] p1_smul_76686_comb;
  wire [31:0] p1_smul_76687_comb;
  wire [31:0] p1_smul_76688_comb;
  wire [31:0] p1_smul_76689_comb;
  wire [31:0] p1_smul_76690_comb;
  wire [31:0] p1_smul_76691_comb;
  wire [31:0] p1_smul_76692_comb;
  wire [31:0] p1_smul_76693_comb;
  wire [31:0] p1_smul_76694_comb;
  wire [31:0] p1_smul_76695_comb;
  wire [31:0] p1_smul_76696_comb;
  wire [31:0] p1_smul_76697_comb;
  wire [31:0] p1_smul_76698_comb;
  wire [31:0] p1_smul_76699_comb;
  wire [31:0] p1_smul_76700_comb;
  wire [31:0] p1_smul_76701_comb;
  wire [31:0] p1_smul_76702_comb;
  wire [31:0] p1_smul_76703_comb;
  wire [31:0] p1_smul_76704_comb;
  wire [31:0] p1_smul_76705_comb;
  wire [31:0] p1_smul_76706_comb;
  wire [31:0] p1_smul_76707_comb;
  wire [31:0] p1_smul_76708_comb;
  wire [31:0] p1_smul_76709_comb;
  wire [31:0] p1_smul_76710_comb;
  wire [31:0] p1_smul_76711_comb;
  wire [31:0] p1_smul_76712_comb;
  wire [31:0] p1_smul_76713_comb;
  wire [31:0] p1_smul_76714_comb;
  wire [31:0] p1_smul_76715_comb;
  wire [31:0] p1_smul_76716_comb;
  wire [31:0] p1_smul_76717_comb;
  wire [31:0] p1_smul_76718_comb;
  wire [31:0] p1_smul_76719_comb;
  wire [31:0] p1_smul_76720_comb;
  wire [31:0] p1_smul_76721_comb;
  wire [31:0] p1_smul_76722_comb;
  wire [31:0] p1_smul_76723_comb;
  wire [31:0] p1_smul_76724_comb;
  wire [31:0] p1_smul_76725_comb;
  wire [31:0] p1_smul_76726_comb;
  wire [31:0] p1_smul_76727_comb;
  wire [31:0] p1_smul_76728_comb;
  wire [31:0] p1_smul_76729_comb;
  wire [31:0] p1_smul_76730_comb;
  wire [31:0] p1_smul_76731_comb;
  wire [31:0] p1_smul_76732_comb;
  wire [31:0] p1_smul_76733_comb;
  wire [31:0] p1_smul_76734_comb;
  wire [31:0] p1_smul_76735_comb;
  wire [31:0] p1_smul_76736_comb;
  wire [31:0] p1_smul_76737_comb;
  wire [31:0] p1_smul_76738_comb;
  wire [31:0] p1_smul_76739_comb;
  wire [31:0] p1_smul_76740_comb;
  wire [31:0] p1_smul_76741_comb;
  wire [31:0] p1_smul_76742_comb;
  wire [31:0] p1_smul_76743_comb;
  wire [31:0] p1_smul_76744_comb;
  wire [31:0] p1_smul_76745_comb;
  wire [31:0] p1_smul_76746_comb;
  wire [31:0] p1_smul_76747_comb;
  wire [31:0] p1_smul_76748_comb;
  wire [31:0] p1_smul_76749_comb;
  wire [31:0] p1_smul_76750_comb;
  wire [31:0] p1_smul_76751_comb;
  wire [31:0] p1_smul_76752_comb;
  wire [31:0] p1_smul_76753_comb;
  wire [31:0] p1_smul_76754_comb;
  wire [31:0] p1_smul_76755_comb;
  wire [31:0] p1_smul_76756_comb;
  wire [31:0] p1_smul_76757_comb;
  wire [31:0] p1_smul_76758_comb;
  wire [31:0] p1_smul_76759_comb;
  wire [31:0] p1_smul_76760_comb;
  wire [31:0] p1_smul_76761_comb;
  wire [31:0] p1_smul_76762_comb;
  wire [31:0] p1_smul_76763_comb;
  wire [31:0] p1_smul_76764_comb;
  wire [31:0] p1_smul_76765_comb;
  wire [31:0] p1_smul_76766_comb;
  wire [31:0] p1_smul_76767_comb;
  wire [31:0] p1_smul_76768_comb;
  wire [31:0] p1_smul_76769_comb;
  wire [31:0] p1_smul_76770_comb;
  wire [31:0] p1_smul_76771_comb;
  wire [31:0] p1_smul_76772_comb;
  wire [31:0] p1_smul_76773_comb;
  wire [31:0] p1_smul_76774_comb;
  wire [31:0] p1_smul_76775_comb;
  wire [31:0] p1_smul_76776_comb;
  wire [31:0] p1_smul_76777_comb;
  wire [31:0] p1_smul_76778_comb;
  wire [31:0] p1_smul_76779_comb;
  wire [31:0] p1_smul_76780_comb;
  wire [31:0] p1_smul_76781_comb;
  wire [31:0] p1_smul_76782_comb;
  wire [31:0] p1_smul_76783_comb;
  wire [31:0] p1_smul_76784_comb;
  wire [31:0] p1_smul_76785_comb;
  wire [31:0] p1_smul_76786_comb;
  wire [31:0] p1_smul_76787_comb;
  wire [31:0] p1_smul_76788_comb;
  wire [31:0] p1_smul_76789_comb;
  wire [31:0] p1_smul_76790_comb;
  wire [31:0] p1_smul_76791_comb;
  wire [31:0] p1_smul_76792_comb;
  wire [31:0] p1_smul_76793_comb;
  wire [31:0] p1_smul_76794_comb;
  wire [31:0] p1_smul_76795_comb;
  wire [31:0] p1_smul_76796_comb;
  wire [31:0] p1_smul_76797_comb;
  wire [31:0] p1_smul_76798_comb;
  wire [31:0] p1_smul_76799_comb;
  wire [31:0] p1_smul_76800_comb;
  wire [31:0] p1_smul_76801_comb;
  wire [31:0] p1_smul_76802_comb;
  wire [31:0] p1_smul_76803_comb;
  wire [31:0] p1_smul_76804_comb;
  wire [31:0] p1_smul_76805_comb;
  wire [31:0] p1_smul_76806_comb;
  wire [31:0] p1_smul_76807_comb;
  wire [31:0] p1_smul_76808_comb;
  wire [31:0] p1_smul_76809_comb;
  wire [31:0] p1_smul_76810_comb;
  wire [31:0] p1_smul_76811_comb;
  wire [31:0] p1_smul_76812_comb;
  wire [31:0] p1_smul_76813_comb;
  wire [31:0] p1_smul_76814_comb;
  wire [31:0] p1_smul_76815_comb;
  wire [31:0] p1_smul_76816_comb;
  wire [31:0] p1_smul_76817_comb;
  wire [31:0] p1_smul_76818_comb;
  wire [31:0] p1_smul_76819_comb;
  wire [31:0] p1_smul_76820_comb;
  wire [31:0] p1_smul_76821_comb;
  wire [31:0] p1_smul_76822_comb;
  wire [31:0] p1_smul_76823_comb;
  wire [31:0] p1_smul_76824_comb;
  wire [31:0] p1_smul_76825_comb;
  wire [31:0] p1_smul_76826_comb;
  wire [31:0] p1_smul_76827_comb;
  wire [31:0] p1_smul_76828_comb;
  wire [31:0] p1_smul_76829_comb;
  wire [31:0] p1_smul_76830_comb;
  wire [31:0] p1_smul_76831_comb;
  wire [31:0] p1_smul_76832_comb;
  wire [31:0] p1_smul_76833_comb;
  wire [31:0] p1_smul_76834_comb;
  wire [31:0] p1_smul_76835_comb;
  wire [31:0] p1_smul_76836_comb;
  wire [31:0] p1_smul_76837_comb;
  wire [31:0] p1_smul_76838_comb;
  wire [31:0] p1_smul_76839_comb;
  wire [31:0] p1_smul_76840_comb;
  wire [31:0] p1_smul_76841_comb;
  wire [31:0] p1_smul_76842_comb;
  wire [31:0] p1_smul_76843_comb;
  wire [31:0] p1_smul_76844_comb;
  wire [31:0] p1_smul_76845_comb;
  wire [31:0] p1_smul_76846_comb;
  wire [31:0] p1_smul_76847_comb;
  wire [31:0] p1_smul_76848_comb;
  wire [31:0] p1_smul_76849_comb;
  wire [31:0] p1_smul_76850_comb;
  wire [31:0] p1_smul_76851_comb;
  wire [31:0] p1_smul_76852_comb;
  wire [31:0] p1_smul_76853_comb;
  wire [31:0] p1_smul_76854_comb;
  wire [31:0] p1_smul_76855_comb;
  wire [31:0] p1_smul_76856_comb;
  wire [31:0] p1_smul_76857_comb;
  wire [31:0] p1_smul_76858_comb;
  wire [31:0] p1_smul_76859_comb;
  wire [31:0] p1_smul_76860_comb;
  wire [31:0] p1_smul_76861_comb;
  wire [31:0] p1_smul_76862_comb;
  wire [31:0] p1_smul_76863_comb;
  wire [31:0] p1_smul_76864_comb;
  wire [31:0] p1_smul_76865_comb;
  wire [31:0] p1_smul_76866_comb;
  wire [31:0] p1_smul_76867_comb;
  wire [31:0] p1_smul_76868_comb;
  wire [31:0] p1_smul_76869_comb;
  wire [31:0] p1_smul_76870_comb;
  wire [31:0] p1_smul_76871_comb;
  wire [31:0] p1_smul_76872_comb;
  wire [31:0] p1_smul_76873_comb;
  wire [31:0] p1_smul_76874_comb;
  wire [31:0] p1_smul_76875_comb;
  wire [31:0] p1_smul_76876_comb;
  wire [31:0] p1_smul_76877_comb;
  wire [31:0] p1_smul_76878_comb;
  wire [31:0] p1_smul_76879_comb;
  wire [31:0] p1_smul_76880_comb;
  wire [31:0] p1_smul_76881_comb;
  wire [31:0] p1_smul_76882_comb;
  wire [31:0] p1_smul_76883_comb;
  wire [31:0] p1_smul_76884_comb;
  wire [31:0] p1_smul_76885_comb;
  wire [31:0] p1_smul_76886_comb;
  wire [31:0] p1_smul_76887_comb;
  wire [31:0] p1_smul_76888_comb;
  wire [31:0] p1_smul_76889_comb;
  wire [31:0] p1_smul_76890_comb;
  wire [31:0] p1_smul_76891_comb;
  wire [31:0] p1_smul_76892_comb;
  wire [31:0] p1_smul_76893_comb;
  wire [31:0] p1_smul_76894_comb;
  wire [31:0] p1_smul_76895_comb;
  wire [31:0] p1_smul_76896_comb;
  wire [31:0] p1_smul_76897_comb;
  wire [31:0] p1_smul_76898_comb;
  wire [31:0] p1_smul_76899_comb;
  wire [31:0] p1_smul_76900_comb;
  wire [31:0] p1_smul_76901_comb;
  wire [31:0] p1_smul_76902_comb;
  wire [31:0] p1_smul_76903_comb;
  wire [31:0] p1_smul_76904_comb;
  wire [31:0] p1_smul_76905_comb;
  wire [31:0] p1_smul_76906_comb;
  wire [31:0] p1_smul_76907_comb;
  wire [31:0] p1_smul_76908_comb;
  wire [31:0] p1_smul_76909_comb;
  wire [31:0] p1_smul_76910_comb;
  wire [31:0] p1_smul_76911_comb;
  wire [31:0] p1_smul_76912_comb;
  wire [31:0] p1_smul_76913_comb;
  wire [31:0] p1_smul_76914_comb;
  wire [31:0] p1_smul_76915_comb;
  wire [31:0] p1_smul_76916_comb;
  wire [31:0] p1_smul_76917_comb;
  wire [31:0] p1_smul_76918_comb;
  wire [31:0] p1_smul_76919_comb;
  wire [31:0] p1_smul_76920_comb;
  wire [31:0] p1_smul_76921_comb;
  wire [31:0] p1_smul_76922_comb;
  wire [31:0] p1_smul_76923_comb;
  wire [31:0] p1_smul_76924_comb;
  wire [31:0] p1_smul_76925_comb;
  wire [31:0] p1_smul_76926_comb;
  wire [31:0] p1_smul_76927_comb;
  wire [31:0] p1_smul_76928_comb;
  wire [31:0] p1_smul_76929_comb;
  wire [31:0] p1_smul_76930_comb;
  wire [31:0] p1_smul_76931_comb;
  wire [31:0] p1_smul_76932_comb;
  wire [31:0] p1_smul_76933_comb;
  wire [31:0] p1_smul_76934_comb;
  wire [31:0] p1_smul_76935_comb;
  wire [31:0] p1_smul_76936_comb;
  wire [31:0] p1_smul_76937_comb;
  wire [31:0] p1_smul_76938_comb;
  wire [31:0] p1_smul_76939_comb;
  wire [31:0] p1_smul_76940_comb;
  wire [31:0] p1_smul_76941_comb;
  wire [31:0] p1_smul_76942_comb;
  wire [31:0] p1_smul_76943_comb;
  wire [31:0] p1_smul_76944_comb;
  wire [31:0] p1_smul_76945_comb;
  wire [31:0] p1_smul_76946_comb;
  wire [31:0] p1_smul_76947_comb;
  wire [31:0] p1_smul_76948_comb;
  wire [31:0] p1_smul_76949_comb;
  wire [31:0] p1_smul_76950_comb;
  wire [31:0] p1_smul_76951_comb;
  wire [31:0] p1_smul_76952_comb;
  wire [31:0] p1_smul_76953_comb;
  wire [31:0] p1_smul_76954_comb;
  wire [31:0] p1_smul_76955_comb;
  wire [31:0] p1_smul_76956_comb;
  wire [31:0] p1_smul_76957_comb;
  wire [31:0] p1_smul_76958_comb;
  wire [31:0] p1_smul_76959_comb;
  wire [31:0] p1_smul_76960_comb;
  wire [31:0] p1_smul_76961_comb;
  wire [31:0] p1_smul_76962_comb;
  wire [31:0] p1_smul_76963_comb;
  wire [31:0] p1_smul_76964_comb;
  wire [31:0] p1_smul_76965_comb;
  wire [31:0] p1_smul_76966_comb;
  wire [31:0] p1_smul_76967_comb;
  wire [31:0] p1_smul_76968_comb;
  wire [31:0] p1_smul_76969_comb;
  wire [31:0] p1_smul_76970_comb;
  wire [31:0] p1_smul_76971_comb;
  assign p1_smul_75972_comb = smul32b_32b_x_32b(p0_TestBlock__A_op0, p0_TestBlock__B_op0);
  assign p1_smul_75973_comb = smul32b_32b_x_32b(p0_TestBlock__A_op1, p0_TestBlock__B_op10);
  assign p1_smul_75974_comb = smul32b_32b_x_32b(p0_TestBlock__A_op2, p0_TestBlock__B_op20);
  assign p1_smul_75975_comb = smul32b_32b_x_32b(p0_TestBlock__A_op3, p0_TestBlock__B_op30);
  assign p1_smul_75976_comb = smul32b_32b_x_32b(p0_TestBlock__A_op0, p0_TestBlock__B_op1);
  assign p1_smul_75977_comb = smul32b_32b_x_32b(p0_TestBlock__A_op1, p0_TestBlock__B_op11);
  assign p1_smul_75978_comb = smul32b_32b_x_32b(p0_TestBlock__A_op2, p0_TestBlock__B_op21);
  assign p1_smul_75979_comb = smul32b_32b_x_32b(p0_TestBlock__A_op3, p0_TestBlock__B_op31);
  assign p1_smul_75980_comb = smul32b_32b_x_32b(p0_TestBlock__A_op0, p0_TestBlock__B_op2);
  assign p1_smul_75981_comb = smul32b_32b_x_32b(p0_TestBlock__A_op1, p0_TestBlock__B_op12);
  assign p1_smul_75982_comb = smul32b_32b_x_32b(p0_TestBlock__A_op2, p0_TestBlock__B_op22);
  assign p1_smul_75983_comb = smul32b_32b_x_32b(p0_TestBlock__A_op3, p0_TestBlock__B_op32);
  assign p1_smul_75984_comb = smul32b_32b_x_32b(p0_TestBlock__A_op0, p0_TestBlock__B_op3);
  assign p1_smul_75985_comb = smul32b_32b_x_32b(p0_TestBlock__A_op1, p0_TestBlock__B_op13);
  assign p1_smul_75986_comb = smul32b_32b_x_32b(p0_TestBlock__A_op2, p0_TestBlock__B_op23);
  assign p1_smul_75987_comb = smul32b_32b_x_32b(p0_TestBlock__A_op3, p0_TestBlock__B_op33);
  assign p1_smul_75988_comb = smul32b_32b_x_32b(p0_TestBlock__A_op0, p0_TestBlock__B_op4);
  assign p1_smul_75989_comb = smul32b_32b_x_32b(p0_TestBlock__A_op1, p0_TestBlock__B_op14);
  assign p1_smul_75990_comb = smul32b_32b_x_32b(p0_TestBlock__A_op2, p0_TestBlock__B_op24);
  assign p1_smul_75991_comb = smul32b_32b_x_32b(p0_TestBlock__A_op3, p0_TestBlock__B_op34);
  assign p1_smul_75992_comb = smul32b_32b_x_32b(p0_TestBlock__A_op0, p0_TestBlock__B_op5);
  assign p1_smul_75993_comb = smul32b_32b_x_32b(p0_TestBlock__A_op1, p0_TestBlock__B_op15);
  assign p1_smul_75994_comb = smul32b_32b_x_32b(p0_TestBlock__A_op2, p0_TestBlock__B_op25);
  assign p1_smul_75995_comb = smul32b_32b_x_32b(p0_TestBlock__A_op3, p0_TestBlock__B_op35);
  assign p1_smul_75996_comb = smul32b_32b_x_32b(p0_TestBlock__A_op0, p0_TestBlock__B_op6);
  assign p1_smul_75997_comb = smul32b_32b_x_32b(p0_TestBlock__A_op1, p0_TestBlock__B_op16);
  assign p1_smul_75998_comb = smul32b_32b_x_32b(p0_TestBlock__A_op2, p0_TestBlock__B_op26);
  assign p1_smul_75999_comb = smul32b_32b_x_32b(p0_TestBlock__A_op3, p0_TestBlock__B_op36);
  assign p1_smul_76000_comb = smul32b_32b_x_32b(p0_TestBlock__A_op0, p0_TestBlock__B_op7);
  assign p1_smul_76001_comb = smul32b_32b_x_32b(p0_TestBlock__A_op1, p0_TestBlock__B_op17);
  assign p1_smul_76002_comb = smul32b_32b_x_32b(p0_TestBlock__A_op2, p0_TestBlock__B_op27);
  assign p1_smul_76003_comb = smul32b_32b_x_32b(p0_TestBlock__A_op3, p0_TestBlock__B_op37);
  assign p1_smul_76004_comb = smul32b_32b_x_32b(p0_TestBlock__A_op0, p0_TestBlock__B_op8);
  assign p1_smul_76005_comb = smul32b_32b_x_32b(p0_TestBlock__A_op1, p0_TestBlock__B_op18);
  assign p1_smul_76006_comb = smul32b_32b_x_32b(p0_TestBlock__A_op2, p0_TestBlock__B_op28);
  assign p1_smul_76007_comb = smul32b_32b_x_32b(p0_TestBlock__A_op3, p0_TestBlock__B_op38);
  assign p1_smul_76008_comb = smul32b_32b_x_32b(p0_TestBlock__A_op0, p0_TestBlock__B_op9);
  assign p1_smul_76009_comb = smul32b_32b_x_32b(p0_TestBlock__A_op1, p0_TestBlock__B_op19);
  assign p1_smul_76010_comb = smul32b_32b_x_32b(p0_TestBlock__A_op2, p0_TestBlock__B_op29);
  assign p1_smul_76011_comb = smul32b_32b_x_32b(p0_TestBlock__A_op3, p0_TestBlock__B_op39);
  assign p1_smul_76012_comb = smul32b_32b_x_32b(p0_TestBlock__A_op10, p0_TestBlock__B_op0);
  assign p1_smul_76013_comb = smul32b_32b_x_32b(p0_TestBlock__A_op11, p0_TestBlock__B_op10);
  assign p1_smul_76014_comb = smul32b_32b_x_32b(p0_TestBlock__A_op12, p0_TestBlock__B_op20);
  assign p1_smul_76015_comb = smul32b_32b_x_32b(p0_TestBlock__A_op13, p0_TestBlock__B_op30);
  assign p1_smul_76016_comb = smul32b_32b_x_32b(p0_TestBlock__A_op10, p0_TestBlock__B_op1);
  assign p1_smul_76017_comb = smul32b_32b_x_32b(p0_TestBlock__A_op11, p0_TestBlock__B_op11);
  assign p1_smul_76018_comb = smul32b_32b_x_32b(p0_TestBlock__A_op12, p0_TestBlock__B_op21);
  assign p1_smul_76019_comb = smul32b_32b_x_32b(p0_TestBlock__A_op13, p0_TestBlock__B_op31);
  assign p1_smul_76020_comb = smul32b_32b_x_32b(p0_TestBlock__A_op10, p0_TestBlock__B_op2);
  assign p1_smul_76021_comb = smul32b_32b_x_32b(p0_TestBlock__A_op11, p0_TestBlock__B_op12);
  assign p1_smul_76022_comb = smul32b_32b_x_32b(p0_TestBlock__A_op12, p0_TestBlock__B_op22);
  assign p1_smul_76023_comb = smul32b_32b_x_32b(p0_TestBlock__A_op13, p0_TestBlock__B_op32);
  assign p1_smul_76024_comb = smul32b_32b_x_32b(p0_TestBlock__A_op10, p0_TestBlock__B_op3);
  assign p1_smul_76025_comb = smul32b_32b_x_32b(p0_TestBlock__A_op11, p0_TestBlock__B_op13);
  assign p1_smul_76026_comb = smul32b_32b_x_32b(p0_TestBlock__A_op12, p0_TestBlock__B_op23);
  assign p1_smul_76027_comb = smul32b_32b_x_32b(p0_TestBlock__A_op13, p0_TestBlock__B_op33);
  assign p1_smul_76028_comb = smul32b_32b_x_32b(p0_TestBlock__A_op10, p0_TestBlock__B_op4);
  assign p1_smul_76029_comb = smul32b_32b_x_32b(p0_TestBlock__A_op11, p0_TestBlock__B_op14);
  assign p1_smul_76030_comb = smul32b_32b_x_32b(p0_TestBlock__A_op12, p0_TestBlock__B_op24);
  assign p1_smul_76031_comb = smul32b_32b_x_32b(p0_TestBlock__A_op13, p0_TestBlock__B_op34);
  assign p1_smul_76032_comb = smul32b_32b_x_32b(p0_TestBlock__A_op10, p0_TestBlock__B_op5);
  assign p1_smul_76033_comb = smul32b_32b_x_32b(p0_TestBlock__A_op11, p0_TestBlock__B_op15);
  assign p1_smul_76034_comb = smul32b_32b_x_32b(p0_TestBlock__A_op12, p0_TestBlock__B_op25);
  assign p1_smul_76035_comb = smul32b_32b_x_32b(p0_TestBlock__A_op13, p0_TestBlock__B_op35);
  assign p1_smul_76036_comb = smul32b_32b_x_32b(p0_TestBlock__A_op10, p0_TestBlock__B_op6);
  assign p1_smul_76037_comb = smul32b_32b_x_32b(p0_TestBlock__A_op11, p0_TestBlock__B_op16);
  assign p1_smul_76038_comb = smul32b_32b_x_32b(p0_TestBlock__A_op12, p0_TestBlock__B_op26);
  assign p1_smul_76039_comb = smul32b_32b_x_32b(p0_TestBlock__A_op13, p0_TestBlock__B_op36);
  assign p1_smul_76040_comb = smul32b_32b_x_32b(p0_TestBlock__A_op10, p0_TestBlock__B_op7);
  assign p1_smul_76041_comb = smul32b_32b_x_32b(p0_TestBlock__A_op11, p0_TestBlock__B_op17);
  assign p1_smul_76042_comb = smul32b_32b_x_32b(p0_TestBlock__A_op12, p0_TestBlock__B_op27);
  assign p1_smul_76043_comb = smul32b_32b_x_32b(p0_TestBlock__A_op13, p0_TestBlock__B_op37);
  assign p1_smul_76044_comb = smul32b_32b_x_32b(p0_TestBlock__A_op10, p0_TestBlock__B_op8);
  assign p1_smul_76045_comb = smul32b_32b_x_32b(p0_TestBlock__A_op11, p0_TestBlock__B_op18);
  assign p1_smul_76046_comb = smul32b_32b_x_32b(p0_TestBlock__A_op12, p0_TestBlock__B_op28);
  assign p1_smul_76047_comb = smul32b_32b_x_32b(p0_TestBlock__A_op13, p0_TestBlock__B_op38);
  assign p1_smul_76048_comb = smul32b_32b_x_32b(p0_TestBlock__A_op10, p0_TestBlock__B_op9);
  assign p1_smul_76049_comb = smul32b_32b_x_32b(p0_TestBlock__A_op11, p0_TestBlock__B_op19);
  assign p1_smul_76050_comb = smul32b_32b_x_32b(p0_TestBlock__A_op12, p0_TestBlock__B_op29);
  assign p1_smul_76051_comb = smul32b_32b_x_32b(p0_TestBlock__A_op13, p0_TestBlock__B_op39);
  assign p1_smul_76052_comb = smul32b_32b_x_32b(p0_TestBlock__A_op20, p0_TestBlock__B_op0);
  assign p1_smul_76053_comb = smul32b_32b_x_32b(p0_TestBlock__A_op21, p0_TestBlock__B_op10);
  assign p1_smul_76054_comb = smul32b_32b_x_32b(p0_TestBlock__A_op22, p0_TestBlock__B_op20);
  assign p1_smul_76055_comb = smul32b_32b_x_32b(p0_TestBlock__A_op23, p0_TestBlock__B_op30);
  assign p1_smul_76056_comb = smul32b_32b_x_32b(p0_TestBlock__A_op20, p0_TestBlock__B_op1);
  assign p1_smul_76057_comb = smul32b_32b_x_32b(p0_TestBlock__A_op21, p0_TestBlock__B_op11);
  assign p1_smul_76058_comb = smul32b_32b_x_32b(p0_TestBlock__A_op22, p0_TestBlock__B_op21);
  assign p1_smul_76059_comb = smul32b_32b_x_32b(p0_TestBlock__A_op23, p0_TestBlock__B_op31);
  assign p1_smul_76060_comb = smul32b_32b_x_32b(p0_TestBlock__A_op20, p0_TestBlock__B_op2);
  assign p1_smul_76061_comb = smul32b_32b_x_32b(p0_TestBlock__A_op21, p0_TestBlock__B_op12);
  assign p1_smul_76062_comb = smul32b_32b_x_32b(p0_TestBlock__A_op22, p0_TestBlock__B_op22);
  assign p1_smul_76063_comb = smul32b_32b_x_32b(p0_TestBlock__A_op23, p0_TestBlock__B_op32);
  assign p1_smul_76064_comb = smul32b_32b_x_32b(p0_TestBlock__A_op20, p0_TestBlock__B_op3);
  assign p1_smul_76065_comb = smul32b_32b_x_32b(p0_TestBlock__A_op21, p0_TestBlock__B_op13);
  assign p1_smul_76066_comb = smul32b_32b_x_32b(p0_TestBlock__A_op22, p0_TestBlock__B_op23);
  assign p1_smul_76067_comb = smul32b_32b_x_32b(p0_TestBlock__A_op23, p0_TestBlock__B_op33);
  assign p1_smul_76068_comb = smul32b_32b_x_32b(p0_TestBlock__A_op20, p0_TestBlock__B_op4);
  assign p1_smul_76069_comb = smul32b_32b_x_32b(p0_TestBlock__A_op21, p0_TestBlock__B_op14);
  assign p1_smul_76070_comb = smul32b_32b_x_32b(p0_TestBlock__A_op22, p0_TestBlock__B_op24);
  assign p1_smul_76071_comb = smul32b_32b_x_32b(p0_TestBlock__A_op23, p0_TestBlock__B_op34);
  assign p1_smul_76072_comb = smul32b_32b_x_32b(p0_TestBlock__A_op20, p0_TestBlock__B_op5);
  assign p1_smul_76073_comb = smul32b_32b_x_32b(p0_TestBlock__A_op21, p0_TestBlock__B_op15);
  assign p1_smul_76074_comb = smul32b_32b_x_32b(p0_TestBlock__A_op22, p0_TestBlock__B_op25);
  assign p1_smul_76075_comb = smul32b_32b_x_32b(p0_TestBlock__A_op23, p0_TestBlock__B_op35);
  assign p1_smul_76076_comb = smul32b_32b_x_32b(p0_TestBlock__A_op20, p0_TestBlock__B_op6);
  assign p1_smul_76077_comb = smul32b_32b_x_32b(p0_TestBlock__A_op21, p0_TestBlock__B_op16);
  assign p1_smul_76078_comb = smul32b_32b_x_32b(p0_TestBlock__A_op22, p0_TestBlock__B_op26);
  assign p1_smul_76079_comb = smul32b_32b_x_32b(p0_TestBlock__A_op23, p0_TestBlock__B_op36);
  assign p1_smul_76080_comb = smul32b_32b_x_32b(p0_TestBlock__A_op20, p0_TestBlock__B_op7);
  assign p1_smul_76081_comb = smul32b_32b_x_32b(p0_TestBlock__A_op21, p0_TestBlock__B_op17);
  assign p1_smul_76082_comb = smul32b_32b_x_32b(p0_TestBlock__A_op22, p0_TestBlock__B_op27);
  assign p1_smul_76083_comb = smul32b_32b_x_32b(p0_TestBlock__A_op23, p0_TestBlock__B_op37);
  assign p1_smul_76084_comb = smul32b_32b_x_32b(p0_TestBlock__A_op20, p0_TestBlock__B_op8);
  assign p1_smul_76085_comb = smul32b_32b_x_32b(p0_TestBlock__A_op21, p0_TestBlock__B_op18);
  assign p1_smul_76086_comb = smul32b_32b_x_32b(p0_TestBlock__A_op22, p0_TestBlock__B_op28);
  assign p1_smul_76087_comb = smul32b_32b_x_32b(p0_TestBlock__A_op23, p0_TestBlock__B_op38);
  assign p1_smul_76088_comb = smul32b_32b_x_32b(p0_TestBlock__A_op20, p0_TestBlock__B_op9);
  assign p1_smul_76089_comb = smul32b_32b_x_32b(p0_TestBlock__A_op21, p0_TestBlock__B_op19);
  assign p1_smul_76090_comb = smul32b_32b_x_32b(p0_TestBlock__A_op22, p0_TestBlock__B_op29);
  assign p1_smul_76091_comb = smul32b_32b_x_32b(p0_TestBlock__A_op23, p0_TestBlock__B_op39);
  assign p1_smul_76092_comb = smul32b_32b_x_32b(p0_TestBlock__A_op30, p0_TestBlock__B_op0);
  assign p1_smul_76093_comb = smul32b_32b_x_32b(p0_TestBlock__A_op31, p0_TestBlock__B_op10);
  assign p1_smul_76094_comb = smul32b_32b_x_32b(p0_TestBlock__A_op32, p0_TestBlock__B_op20);
  assign p1_smul_76095_comb = smul32b_32b_x_32b(p0_TestBlock__A_op33, p0_TestBlock__B_op30);
  assign p1_smul_76096_comb = smul32b_32b_x_32b(p0_TestBlock__A_op30, p0_TestBlock__B_op1);
  assign p1_smul_76097_comb = smul32b_32b_x_32b(p0_TestBlock__A_op31, p0_TestBlock__B_op11);
  assign p1_smul_76098_comb = smul32b_32b_x_32b(p0_TestBlock__A_op32, p0_TestBlock__B_op21);
  assign p1_smul_76099_comb = smul32b_32b_x_32b(p0_TestBlock__A_op33, p0_TestBlock__B_op31);
  assign p1_smul_76100_comb = smul32b_32b_x_32b(p0_TestBlock__A_op30, p0_TestBlock__B_op2);
  assign p1_smul_76101_comb = smul32b_32b_x_32b(p0_TestBlock__A_op31, p0_TestBlock__B_op12);
  assign p1_smul_76102_comb = smul32b_32b_x_32b(p0_TestBlock__A_op32, p0_TestBlock__B_op22);
  assign p1_smul_76103_comb = smul32b_32b_x_32b(p0_TestBlock__A_op33, p0_TestBlock__B_op32);
  assign p1_smul_76104_comb = smul32b_32b_x_32b(p0_TestBlock__A_op30, p0_TestBlock__B_op3);
  assign p1_smul_76105_comb = smul32b_32b_x_32b(p0_TestBlock__A_op31, p0_TestBlock__B_op13);
  assign p1_smul_76106_comb = smul32b_32b_x_32b(p0_TestBlock__A_op32, p0_TestBlock__B_op23);
  assign p1_smul_76107_comb = smul32b_32b_x_32b(p0_TestBlock__A_op33, p0_TestBlock__B_op33);
  assign p1_smul_76108_comb = smul32b_32b_x_32b(p0_TestBlock__A_op30, p0_TestBlock__B_op4);
  assign p1_smul_76109_comb = smul32b_32b_x_32b(p0_TestBlock__A_op31, p0_TestBlock__B_op14);
  assign p1_smul_76110_comb = smul32b_32b_x_32b(p0_TestBlock__A_op32, p0_TestBlock__B_op24);
  assign p1_smul_76111_comb = smul32b_32b_x_32b(p0_TestBlock__A_op33, p0_TestBlock__B_op34);
  assign p1_smul_76112_comb = smul32b_32b_x_32b(p0_TestBlock__A_op30, p0_TestBlock__B_op5);
  assign p1_smul_76113_comb = smul32b_32b_x_32b(p0_TestBlock__A_op31, p0_TestBlock__B_op15);
  assign p1_smul_76114_comb = smul32b_32b_x_32b(p0_TestBlock__A_op32, p0_TestBlock__B_op25);
  assign p1_smul_76115_comb = smul32b_32b_x_32b(p0_TestBlock__A_op33, p0_TestBlock__B_op35);
  assign p1_smul_76116_comb = smul32b_32b_x_32b(p0_TestBlock__A_op30, p0_TestBlock__B_op6);
  assign p1_smul_76117_comb = smul32b_32b_x_32b(p0_TestBlock__A_op31, p0_TestBlock__B_op16);
  assign p1_smul_76118_comb = smul32b_32b_x_32b(p0_TestBlock__A_op32, p0_TestBlock__B_op26);
  assign p1_smul_76119_comb = smul32b_32b_x_32b(p0_TestBlock__A_op33, p0_TestBlock__B_op36);
  assign p1_smul_76120_comb = smul32b_32b_x_32b(p0_TestBlock__A_op30, p0_TestBlock__B_op7);
  assign p1_smul_76121_comb = smul32b_32b_x_32b(p0_TestBlock__A_op31, p0_TestBlock__B_op17);
  assign p1_smul_76122_comb = smul32b_32b_x_32b(p0_TestBlock__A_op32, p0_TestBlock__B_op27);
  assign p1_smul_76123_comb = smul32b_32b_x_32b(p0_TestBlock__A_op33, p0_TestBlock__B_op37);
  assign p1_smul_76124_comb = smul32b_32b_x_32b(p0_TestBlock__A_op30, p0_TestBlock__B_op8);
  assign p1_smul_76125_comb = smul32b_32b_x_32b(p0_TestBlock__A_op31, p0_TestBlock__B_op18);
  assign p1_smul_76126_comb = smul32b_32b_x_32b(p0_TestBlock__A_op32, p0_TestBlock__B_op28);
  assign p1_smul_76127_comb = smul32b_32b_x_32b(p0_TestBlock__A_op33, p0_TestBlock__B_op38);
  assign p1_smul_76128_comb = smul32b_32b_x_32b(p0_TestBlock__A_op30, p0_TestBlock__B_op9);
  assign p1_smul_76129_comb = smul32b_32b_x_32b(p0_TestBlock__A_op31, p0_TestBlock__B_op19);
  assign p1_smul_76130_comb = smul32b_32b_x_32b(p0_TestBlock__A_op32, p0_TestBlock__B_op29);
  assign p1_smul_76131_comb = smul32b_32b_x_32b(p0_TestBlock__A_op33, p0_TestBlock__B_op39);
  assign p1_smul_76132_comb = smul32b_32b_x_32b(p0_TestBlock__A_op40, p0_TestBlock__B_op0);
  assign p1_smul_76133_comb = smul32b_32b_x_32b(p0_TestBlock__A_op41, p0_TestBlock__B_op10);
  assign p1_smul_76134_comb = smul32b_32b_x_32b(p0_TestBlock__A_op42, p0_TestBlock__B_op20);
  assign p1_smul_76135_comb = smul32b_32b_x_32b(p0_TestBlock__A_op43, p0_TestBlock__B_op30);
  assign p1_smul_76136_comb = smul32b_32b_x_32b(p0_TestBlock__A_op40, p0_TestBlock__B_op1);
  assign p1_smul_76137_comb = smul32b_32b_x_32b(p0_TestBlock__A_op41, p0_TestBlock__B_op11);
  assign p1_smul_76138_comb = smul32b_32b_x_32b(p0_TestBlock__A_op42, p0_TestBlock__B_op21);
  assign p1_smul_76139_comb = smul32b_32b_x_32b(p0_TestBlock__A_op43, p0_TestBlock__B_op31);
  assign p1_smul_76140_comb = smul32b_32b_x_32b(p0_TestBlock__A_op40, p0_TestBlock__B_op2);
  assign p1_smul_76141_comb = smul32b_32b_x_32b(p0_TestBlock__A_op41, p0_TestBlock__B_op12);
  assign p1_smul_76142_comb = smul32b_32b_x_32b(p0_TestBlock__A_op42, p0_TestBlock__B_op22);
  assign p1_smul_76143_comb = smul32b_32b_x_32b(p0_TestBlock__A_op43, p0_TestBlock__B_op32);
  assign p1_smul_76144_comb = smul32b_32b_x_32b(p0_TestBlock__A_op40, p0_TestBlock__B_op3);
  assign p1_smul_76145_comb = smul32b_32b_x_32b(p0_TestBlock__A_op41, p0_TestBlock__B_op13);
  assign p1_smul_76146_comb = smul32b_32b_x_32b(p0_TestBlock__A_op42, p0_TestBlock__B_op23);
  assign p1_smul_76147_comb = smul32b_32b_x_32b(p0_TestBlock__A_op43, p0_TestBlock__B_op33);
  assign p1_smul_76148_comb = smul32b_32b_x_32b(p0_TestBlock__A_op40, p0_TestBlock__B_op4);
  assign p1_smul_76149_comb = smul32b_32b_x_32b(p0_TestBlock__A_op41, p0_TestBlock__B_op14);
  assign p1_smul_76150_comb = smul32b_32b_x_32b(p0_TestBlock__A_op42, p0_TestBlock__B_op24);
  assign p1_smul_76151_comb = smul32b_32b_x_32b(p0_TestBlock__A_op43, p0_TestBlock__B_op34);
  assign p1_smul_76152_comb = smul32b_32b_x_32b(p0_TestBlock__A_op40, p0_TestBlock__B_op5);
  assign p1_smul_76153_comb = smul32b_32b_x_32b(p0_TestBlock__A_op41, p0_TestBlock__B_op15);
  assign p1_smul_76154_comb = smul32b_32b_x_32b(p0_TestBlock__A_op42, p0_TestBlock__B_op25);
  assign p1_smul_76155_comb = smul32b_32b_x_32b(p0_TestBlock__A_op43, p0_TestBlock__B_op35);
  assign p1_smul_76156_comb = smul32b_32b_x_32b(p0_TestBlock__A_op40, p0_TestBlock__B_op6);
  assign p1_smul_76157_comb = smul32b_32b_x_32b(p0_TestBlock__A_op41, p0_TestBlock__B_op16);
  assign p1_smul_76158_comb = smul32b_32b_x_32b(p0_TestBlock__A_op42, p0_TestBlock__B_op26);
  assign p1_smul_76159_comb = smul32b_32b_x_32b(p0_TestBlock__A_op43, p0_TestBlock__B_op36);
  assign p1_smul_76160_comb = smul32b_32b_x_32b(p0_TestBlock__A_op40, p0_TestBlock__B_op7);
  assign p1_smul_76161_comb = smul32b_32b_x_32b(p0_TestBlock__A_op41, p0_TestBlock__B_op17);
  assign p1_smul_76162_comb = smul32b_32b_x_32b(p0_TestBlock__A_op42, p0_TestBlock__B_op27);
  assign p1_smul_76163_comb = smul32b_32b_x_32b(p0_TestBlock__A_op43, p0_TestBlock__B_op37);
  assign p1_smul_76164_comb = smul32b_32b_x_32b(p0_TestBlock__A_op40, p0_TestBlock__B_op8);
  assign p1_smul_76165_comb = smul32b_32b_x_32b(p0_TestBlock__A_op41, p0_TestBlock__B_op18);
  assign p1_smul_76166_comb = smul32b_32b_x_32b(p0_TestBlock__A_op42, p0_TestBlock__B_op28);
  assign p1_smul_76167_comb = smul32b_32b_x_32b(p0_TestBlock__A_op43, p0_TestBlock__B_op38);
  assign p1_smul_76168_comb = smul32b_32b_x_32b(p0_TestBlock__A_op40, p0_TestBlock__B_op9);
  assign p1_smul_76169_comb = smul32b_32b_x_32b(p0_TestBlock__A_op41, p0_TestBlock__B_op19);
  assign p1_smul_76170_comb = smul32b_32b_x_32b(p0_TestBlock__A_op42, p0_TestBlock__B_op29);
  assign p1_smul_76171_comb = smul32b_32b_x_32b(p0_TestBlock__A_op43, p0_TestBlock__B_op39);
  assign p1_smul_76172_comb = smul32b_32b_x_32b(p0_TestBlock__A_op50, p0_TestBlock__B_op0);
  assign p1_smul_76173_comb = smul32b_32b_x_32b(p0_TestBlock__A_op51, p0_TestBlock__B_op10);
  assign p1_smul_76174_comb = smul32b_32b_x_32b(p0_TestBlock__A_op52, p0_TestBlock__B_op20);
  assign p1_smul_76175_comb = smul32b_32b_x_32b(p0_TestBlock__A_op53, p0_TestBlock__B_op30);
  assign p1_smul_76176_comb = smul32b_32b_x_32b(p0_TestBlock__A_op50, p0_TestBlock__B_op1);
  assign p1_smul_76177_comb = smul32b_32b_x_32b(p0_TestBlock__A_op51, p0_TestBlock__B_op11);
  assign p1_smul_76178_comb = smul32b_32b_x_32b(p0_TestBlock__A_op52, p0_TestBlock__B_op21);
  assign p1_smul_76179_comb = smul32b_32b_x_32b(p0_TestBlock__A_op53, p0_TestBlock__B_op31);
  assign p1_smul_76180_comb = smul32b_32b_x_32b(p0_TestBlock__A_op50, p0_TestBlock__B_op2);
  assign p1_smul_76181_comb = smul32b_32b_x_32b(p0_TestBlock__A_op51, p0_TestBlock__B_op12);
  assign p1_smul_76182_comb = smul32b_32b_x_32b(p0_TestBlock__A_op52, p0_TestBlock__B_op22);
  assign p1_smul_76183_comb = smul32b_32b_x_32b(p0_TestBlock__A_op53, p0_TestBlock__B_op32);
  assign p1_smul_76184_comb = smul32b_32b_x_32b(p0_TestBlock__A_op50, p0_TestBlock__B_op3);
  assign p1_smul_76185_comb = smul32b_32b_x_32b(p0_TestBlock__A_op51, p0_TestBlock__B_op13);
  assign p1_smul_76186_comb = smul32b_32b_x_32b(p0_TestBlock__A_op52, p0_TestBlock__B_op23);
  assign p1_smul_76187_comb = smul32b_32b_x_32b(p0_TestBlock__A_op53, p0_TestBlock__B_op33);
  assign p1_smul_76188_comb = smul32b_32b_x_32b(p0_TestBlock__A_op50, p0_TestBlock__B_op4);
  assign p1_smul_76189_comb = smul32b_32b_x_32b(p0_TestBlock__A_op51, p0_TestBlock__B_op14);
  assign p1_smul_76190_comb = smul32b_32b_x_32b(p0_TestBlock__A_op52, p0_TestBlock__B_op24);
  assign p1_smul_76191_comb = smul32b_32b_x_32b(p0_TestBlock__A_op53, p0_TestBlock__B_op34);
  assign p1_smul_76192_comb = smul32b_32b_x_32b(p0_TestBlock__A_op50, p0_TestBlock__B_op5);
  assign p1_smul_76193_comb = smul32b_32b_x_32b(p0_TestBlock__A_op51, p0_TestBlock__B_op15);
  assign p1_smul_76194_comb = smul32b_32b_x_32b(p0_TestBlock__A_op52, p0_TestBlock__B_op25);
  assign p1_smul_76195_comb = smul32b_32b_x_32b(p0_TestBlock__A_op53, p0_TestBlock__B_op35);
  assign p1_smul_76196_comb = smul32b_32b_x_32b(p0_TestBlock__A_op50, p0_TestBlock__B_op6);
  assign p1_smul_76197_comb = smul32b_32b_x_32b(p0_TestBlock__A_op51, p0_TestBlock__B_op16);
  assign p1_smul_76198_comb = smul32b_32b_x_32b(p0_TestBlock__A_op52, p0_TestBlock__B_op26);
  assign p1_smul_76199_comb = smul32b_32b_x_32b(p0_TestBlock__A_op53, p0_TestBlock__B_op36);
  assign p1_smul_76200_comb = smul32b_32b_x_32b(p0_TestBlock__A_op50, p0_TestBlock__B_op7);
  assign p1_smul_76201_comb = smul32b_32b_x_32b(p0_TestBlock__A_op51, p0_TestBlock__B_op17);
  assign p1_smul_76202_comb = smul32b_32b_x_32b(p0_TestBlock__A_op52, p0_TestBlock__B_op27);
  assign p1_smul_76203_comb = smul32b_32b_x_32b(p0_TestBlock__A_op53, p0_TestBlock__B_op37);
  assign p1_smul_76204_comb = smul32b_32b_x_32b(p0_TestBlock__A_op50, p0_TestBlock__B_op8);
  assign p1_smul_76205_comb = smul32b_32b_x_32b(p0_TestBlock__A_op51, p0_TestBlock__B_op18);
  assign p1_smul_76206_comb = smul32b_32b_x_32b(p0_TestBlock__A_op52, p0_TestBlock__B_op28);
  assign p1_smul_76207_comb = smul32b_32b_x_32b(p0_TestBlock__A_op53, p0_TestBlock__B_op38);
  assign p1_smul_76208_comb = smul32b_32b_x_32b(p0_TestBlock__A_op50, p0_TestBlock__B_op9);
  assign p1_smul_76209_comb = smul32b_32b_x_32b(p0_TestBlock__A_op51, p0_TestBlock__B_op19);
  assign p1_smul_76210_comb = smul32b_32b_x_32b(p0_TestBlock__A_op52, p0_TestBlock__B_op29);
  assign p1_smul_76211_comb = smul32b_32b_x_32b(p0_TestBlock__A_op53, p0_TestBlock__B_op39);
  assign p1_smul_76212_comb = smul32b_32b_x_32b(p0_TestBlock__A_op60, p0_TestBlock__B_op0);
  assign p1_smul_76213_comb = smul32b_32b_x_32b(p0_TestBlock__A_op61, p0_TestBlock__B_op10);
  assign p1_smul_76214_comb = smul32b_32b_x_32b(p0_TestBlock__A_op62, p0_TestBlock__B_op20);
  assign p1_smul_76215_comb = smul32b_32b_x_32b(p0_TestBlock__A_op63, p0_TestBlock__B_op30);
  assign p1_smul_76216_comb = smul32b_32b_x_32b(p0_TestBlock__A_op60, p0_TestBlock__B_op1);
  assign p1_smul_76217_comb = smul32b_32b_x_32b(p0_TestBlock__A_op61, p0_TestBlock__B_op11);
  assign p1_smul_76218_comb = smul32b_32b_x_32b(p0_TestBlock__A_op62, p0_TestBlock__B_op21);
  assign p1_smul_76219_comb = smul32b_32b_x_32b(p0_TestBlock__A_op63, p0_TestBlock__B_op31);
  assign p1_smul_76220_comb = smul32b_32b_x_32b(p0_TestBlock__A_op60, p0_TestBlock__B_op2);
  assign p1_smul_76221_comb = smul32b_32b_x_32b(p0_TestBlock__A_op61, p0_TestBlock__B_op12);
  assign p1_smul_76222_comb = smul32b_32b_x_32b(p0_TestBlock__A_op62, p0_TestBlock__B_op22);
  assign p1_smul_76223_comb = smul32b_32b_x_32b(p0_TestBlock__A_op63, p0_TestBlock__B_op32);
  assign p1_smul_76224_comb = smul32b_32b_x_32b(p0_TestBlock__A_op60, p0_TestBlock__B_op3);
  assign p1_smul_76225_comb = smul32b_32b_x_32b(p0_TestBlock__A_op61, p0_TestBlock__B_op13);
  assign p1_smul_76226_comb = smul32b_32b_x_32b(p0_TestBlock__A_op62, p0_TestBlock__B_op23);
  assign p1_smul_76227_comb = smul32b_32b_x_32b(p0_TestBlock__A_op63, p0_TestBlock__B_op33);
  assign p1_smul_76228_comb = smul32b_32b_x_32b(p0_TestBlock__A_op60, p0_TestBlock__B_op4);
  assign p1_smul_76229_comb = smul32b_32b_x_32b(p0_TestBlock__A_op61, p0_TestBlock__B_op14);
  assign p1_smul_76230_comb = smul32b_32b_x_32b(p0_TestBlock__A_op62, p0_TestBlock__B_op24);
  assign p1_smul_76231_comb = smul32b_32b_x_32b(p0_TestBlock__A_op63, p0_TestBlock__B_op34);
  assign p1_smul_76232_comb = smul32b_32b_x_32b(p0_TestBlock__A_op60, p0_TestBlock__B_op5);
  assign p1_smul_76233_comb = smul32b_32b_x_32b(p0_TestBlock__A_op61, p0_TestBlock__B_op15);
  assign p1_smul_76234_comb = smul32b_32b_x_32b(p0_TestBlock__A_op62, p0_TestBlock__B_op25);
  assign p1_smul_76235_comb = smul32b_32b_x_32b(p0_TestBlock__A_op63, p0_TestBlock__B_op35);
  assign p1_smul_76236_comb = smul32b_32b_x_32b(p0_TestBlock__A_op60, p0_TestBlock__B_op6);
  assign p1_smul_76237_comb = smul32b_32b_x_32b(p0_TestBlock__A_op61, p0_TestBlock__B_op16);
  assign p1_smul_76238_comb = smul32b_32b_x_32b(p0_TestBlock__A_op62, p0_TestBlock__B_op26);
  assign p1_smul_76239_comb = smul32b_32b_x_32b(p0_TestBlock__A_op63, p0_TestBlock__B_op36);
  assign p1_smul_76240_comb = smul32b_32b_x_32b(p0_TestBlock__A_op60, p0_TestBlock__B_op7);
  assign p1_smul_76241_comb = smul32b_32b_x_32b(p0_TestBlock__A_op61, p0_TestBlock__B_op17);
  assign p1_smul_76242_comb = smul32b_32b_x_32b(p0_TestBlock__A_op62, p0_TestBlock__B_op27);
  assign p1_smul_76243_comb = smul32b_32b_x_32b(p0_TestBlock__A_op63, p0_TestBlock__B_op37);
  assign p1_smul_76244_comb = smul32b_32b_x_32b(p0_TestBlock__A_op60, p0_TestBlock__B_op8);
  assign p1_smul_76245_comb = smul32b_32b_x_32b(p0_TestBlock__A_op61, p0_TestBlock__B_op18);
  assign p1_smul_76246_comb = smul32b_32b_x_32b(p0_TestBlock__A_op62, p0_TestBlock__B_op28);
  assign p1_smul_76247_comb = smul32b_32b_x_32b(p0_TestBlock__A_op63, p0_TestBlock__B_op38);
  assign p1_smul_76248_comb = smul32b_32b_x_32b(p0_TestBlock__A_op60, p0_TestBlock__B_op9);
  assign p1_smul_76249_comb = smul32b_32b_x_32b(p0_TestBlock__A_op61, p0_TestBlock__B_op19);
  assign p1_smul_76250_comb = smul32b_32b_x_32b(p0_TestBlock__A_op62, p0_TestBlock__B_op29);
  assign p1_smul_76251_comb = smul32b_32b_x_32b(p0_TestBlock__A_op63, p0_TestBlock__B_op39);
  assign p1_smul_76252_comb = smul32b_32b_x_32b(p0_TestBlock__A_op70, p0_TestBlock__B_op0);
  assign p1_smul_76253_comb = smul32b_32b_x_32b(p0_TestBlock__A_op71, p0_TestBlock__B_op10);
  assign p1_smul_76254_comb = smul32b_32b_x_32b(p0_TestBlock__A_op72, p0_TestBlock__B_op20);
  assign p1_smul_76255_comb = smul32b_32b_x_32b(p0_TestBlock__A_op73, p0_TestBlock__B_op30);
  assign p1_smul_76256_comb = smul32b_32b_x_32b(p0_TestBlock__A_op70, p0_TestBlock__B_op1);
  assign p1_smul_76257_comb = smul32b_32b_x_32b(p0_TestBlock__A_op71, p0_TestBlock__B_op11);
  assign p1_smul_76258_comb = smul32b_32b_x_32b(p0_TestBlock__A_op72, p0_TestBlock__B_op21);
  assign p1_smul_76259_comb = smul32b_32b_x_32b(p0_TestBlock__A_op73, p0_TestBlock__B_op31);
  assign p1_smul_76260_comb = smul32b_32b_x_32b(p0_TestBlock__A_op70, p0_TestBlock__B_op2);
  assign p1_smul_76261_comb = smul32b_32b_x_32b(p0_TestBlock__A_op71, p0_TestBlock__B_op12);
  assign p1_smul_76262_comb = smul32b_32b_x_32b(p0_TestBlock__A_op72, p0_TestBlock__B_op22);
  assign p1_smul_76263_comb = smul32b_32b_x_32b(p0_TestBlock__A_op73, p0_TestBlock__B_op32);
  assign p1_smul_76264_comb = smul32b_32b_x_32b(p0_TestBlock__A_op70, p0_TestBlock__B_op3);
  assign p1_smul_76265_comb = smul32b_32b_x_32b(p0_TestBlock__A_op71, p0_TestBlock__B_op13);
  assign p1_smul_76266_comb = smul32b_32b_x_32b(p0_TestBlock__A_op72, p0_TestBlock__B_op23);
  assign p1_smul_76267_comb = smul32b_32b_x_32b(p0_TestBlock__A_op73, p0_TestBlock__B_op33);
  assign p1_smul_76268_comb = smul32b_32b_x_32b(p0_TestBlock__A_op70, p0_TestBlock__B_op4);
  assign p1_smul_76269_comb = smul32b_32b_x_32b(p0_TestBlock__A_op71, p0_TestBlock__B_op14);
  assign p1_smul_76270_comb = smul32b_32b_x_32b(p0_TestBlock__A_op72, p0_TestBlock__B_op24);
  assign p1_smul_76271_comb = smul32b_32b_x_32b(p0_TestBlock__A_op73, p0_TestBlock__B_op34);
  assign p1_smul_76272_comb = smul32b_32b_x_32b(p0_TestBlock__A_op70, p0_TestBlock__B_op5);
  assign p1_smul_76273_comb = smul32b_32b_x_32b(p0_TestBlock__A_op71, p0_TestBlock__B_op15);
  assign p1_smul_76274_comb = smul32b_32b_x_32b(p0_TestBlock__A_op72, p0_TestBlock__B_op25);
  assign p1_smul_76275_comb = smul32b_32b_x_32b(p0_TestBlock__A_op73, p0_TestBlock__B_op35);
  assign p1_smul_76276_comb = smul32b_32b_x_32b(p0_TestBlock__A_op70, p0_TestBlock__B_op6);
  assign p1_smul_76277_comb = smul32b_32b_x_32b(p0_TestBlock__A_op71, p0_TestBlock__B_op16);
  assign p1_smul_76278_comb = smul32b_32b_x_32b(p0_TestBlock__A_op72, p0_TestBlock__B_op26);
  assign p1_smul_76279_comb = smul32b_32b_x_32b(p0_TestBlock__A_op73, p0_TestBlock__B_op36);
  assign p1_smul_76280_comb = smul32b_32b_x_32b(p0_TestBlock__A_op70, p0_TestBlock__B_op7);
  assign p1_smul_76281_comb = smul32b_32b_x_32b(p0_TestBlock__A_op71, p0_TestBlock__B_op17);
  assign p1_smul_76282_comb = smul32b_32b_x_32b(p0_TestBlock__A_op72, p0_TestBlock__B_op27);
  assign p1_smul_76283_comb = smul32b_32b_x_32b(p0_TestBlock__A_op73, p0_TestBlock__B_op37);
  assign p1_smul_76284_comb = smul32b_32b_x_32b(p0_TestBlock__A_op70, p0_TestBlock__B_op8);
  assign p1_smul_76285_comb = smul32b_32b_x_32b(p0_TestBlock__A_op71, p0_TestBlock__B_op18);
  assign p1_smul_76286_comb = smul32b_32b_x_32b(p0_TestBlock__A_op72, p0_TestBlock__B_op28);
  assign p1_smul_76287_comb = smul32b_32b_x_32b(p0_TestBlock__A_op73, p0_TestBlock__B_op38);
  assign p1_smul_76288_comb = smul32b_32b_x_32b(p0_TestBlock__A_op70, p0_TestBlock__B_op9);
  assign p1_smul_76289_comb = smul32b_32b_x_32b(p0_TestBlock__A_op71, p0_TestBlock__B_op19);
  assign p1_smul_76290_comb = smul32b_32b_x_32b(p0_TestBlock__A_op72, p0_TestBlock__B_op29);
  assign p1_smul_76291_comb = smul32b_32b_x_32b(p0_TestBlock__A_op73, p0_TestBlock__B_op39);
  assign p1_smul_76292_comb = smul32b_32b_x_32b(p0_TestBlock__A_op80, p0_TestBlock__B_op0);
  assign p1_smul_76293_comb = smul32b_32b_x_32b(p0_TestBlock__A_op81, p0_TestBlock__B_op10);
  assign p1_smul_76294_comb = smul32b_32b_x_32b(p0_TestBlock__A_op82, p0_TestBlock__B_op20);
  assign p1_smul_76295_comb = smul32b_32b_x_32b(p0_TestBlock__A_op83, p0_TestBlock__B_op30);
  assign p1_smul_76296_comb = smul32b_32b_x_32b(p0_TestBlock__A_op80, p0_TestBlock__B_op1);
  assign p1_smul_76297_comb = smul32b_32b_x_32b(p0_TestBlock__A_op81, p0_TestBlock__B_op11);
  assign p1_smul_76298_comb = smul32b_32b_x_32b(p0_TestBlock__A_op82, p0_TestBlock__B_op21);
  assign p1_smul_76299_comb = smul32b_32b_x_32b(p0_TestBlock__A_op83, p0_TestBlock__B_op31);
  assign p1_smul_76300_comb = smul32b_32b_x_32b(p0_TestBlock__A_op80, p0_TestBlock__B_op2);
  assign p1_smul_76301_comb = smul32b_32b_x_32b(p0_TestBlock__A_op81, p0_TestBlock__B_op12);
  assign p1_smul_76302_comb = smul32b_32b_x_32b(p0_TestBlock__A_op82, p0_TestBlock__B_op22);
  assign p1_smul_76303_comb = smul32b_32b_x_32b(p0_TestBlock__A_op83, p0_TestBlock__B_op32);
  assign p1_smul_76304_comb = smul32b_32b_x_32b(p0_TestBlock__A_op80, p0_TestBlock__B_op3);
  assign p1_smul_76305_comb = smul32b_32b_x_32b(p0_TestBlock__A_op81, p0_TestBlock__B_op13);
  assign p1_smul_76306_comb = smul32b_32b_x_32b(p0_TestBlock__A_op82, p0_TestBlock__B_op23);
  assign p1_smul_76307_comb = smul32b_32b_x_32b(p0_TestBlock__A_op83, p0_TestBlock__B_op33);
  assign p1_smul_76308_comb = smul32b_32b_x_32b(p0_TestBlock__A_op80, p0_TestBlock__B_op4);
  assign p1_smul_76309_comb = smul32b_32b_x_32b(p0_TestBlock__A_op81, p0_TestBlock__B_op14);
  assign p1_smul_76310_comb = smul32b_32b_x_32b(p0_TestBlock__A_op82, p0_TestBlock__B_op24);
  assign p1_smul_76311_comb = smul32b_32b_x_32b(p0_TestBlock__A_op83, p0_TestBlock__B_op34);
  assign p1_smul_76312_comb = smul32b_32b_x_32b(p0_TestBlock__A_op80, p0_TestBlock__B_op5);
  assign p1_smul_76313_comb = smul32b_32b_x_32b(p0_TestBlock__A_op81, p0_TestBlock__B_op15);
  assign p1_smul_76314_comb = smul32b_32b_x_32b(p0_TestBlock__A_op82, p0_TestBlock__B_op25);
  assign p1_smul_76315_comb = smul32b_32b_x_32b(p0_TestBlock__A_op83, p0_TestBlock__B_op35);
  assign p1_smul_76316_comb = smul32b_32b_x_32b(p0_TestBlock__A_op80, p0_TestBlock__B_op6);
  assign p1_smul_76317_comb = smul32b_32b_x_32b(p0_TestBlock__A_op81, p0_TestBlock__B_op16);
  assign p1_smul_76318_comb = smul32b_32b_x_32b(p0_TestBlock__A_op82, p0_TestBlock__B_op26);
  assign p1_smul_76319_comb = smul32b_32b_x_32b(p0_TestBlock__A_op83, p0_TestBlock__B_op36);
  assign p1_smul_76320_comb = smul32b_32b_x_32b(p0_TestBlock__A_op80, p0_TestBlock__B_op7);
  assign p1_smul_76321_comb = smul32b_32b_x_32b(p0_TestBlock__A_op81, p0_TestBlock__B_op17);
  assign p1_smul_76322_comb = smul32b_32b_x_32b(p0_TestBlock__A_op82, p0_TestBlock__B_op27);
  assign p1_smul_76323_comb = smul32b_32b_x_32b(p0_TestBlock__A_op83, p0_TestBlock__B_op37);
  assign p1_smul_76324_comb = smul32b_32b_x_32b(p0_TestBlock__A_op80, p0_TestBlock__B_op8);
  assign p1_smul_76325_comb = smul32b_32b_x_32b(p0_TestBlock__A_op81, p0_TestBlock__B_op18);
  assign p1_smul_76326_comb = smul32b_32b_x_32b(p0_TestBlock__A_op82, p0_TestBlock__B_op28);
  assign p1_smul_76327_comb = smul32b_32b_x_32b(p0_TestBlock__A_op83, p0_TestBlock__B_op38);
  assign p1_smul_76328_comb = smul32b_32b_x_32b(p0_TestBlock__A_op80, p0_TestBlock__B_op9);
  assign p1_smul_76329_comb = smul32b_32b_x_32b(p0_TestBlock__A_op81, p0_TestBlock__B_op19);
  assign p1_smul_76330_comb = smul32b_32b_x_32b(p0_TestBlock__A_op82, p0_TestBlock__B_op29);
  assign p1_smul_76331_comb = smul32b_32b_x_32b(p0_TestBlock__A_op83, p0_TestBlock__B_op39);
  assign p1_smul_76332_comb = smul32b_32b_x_32b(p0_TestBlock__A_op90, p0_TestBlock__B_op0);
  assign p1_smul_76333_comb = smul32b_32b_x_32b(p0_TestBlock__A_op91, p0_TestBlock__B_op10);
  assign p1_smul_76334_comb = smul32b_32b_x_32b(p0_TestBlock__A_op92, p0_TestBlock__B_op20);
  assign p1_smul_76335_comb = smul32b_32b_x_32b(p0_TestBlock__A_op93, p0_TestBlock__B_op30);
  assign p1_smul_76336_comb = smul32b_32b_x_32b(p0_TestBlock__A_op90, p0_TestBlock__B_op1);
  assign p1_smul_76337_comb = smul32b_32b_x_32b(p0_TestBlock__A_op91, p0_TestBlock__B_op11);
  assign p1_smul_76338_comb = smul32b_32b_x_32b(p0_TestBlock__A_op92, p0_TestBlock__B_op21);
  assign p1_smul_76339_comb = smul32b_32b_x_32b(p0_TestBlock__A_op93, p0_TestBlock__B_op31);
  assign p1_smul_76340_comb = smul32b_32b_x_32b(p0_TestBlock__A_op90, p0_TestBlock__B_op2);
  assign p1_smul_76341_comb = smul32b_32b_x_32b(p0_TestBlock__A_op91, p0_TestBlock__B_op12);
  assign p1_smul_76342_comb = smul32b_32b_x_32b(p0_TestBlock__A_op92, p0_TestBlock__B_op22);
  assign p1_smul_76343_comb = smul32b_32b_x_32b(p0_TestBlock__A_op93, p0_TestBlock__B_op32);
  assign p1_smul_76344_comb = smul32b_32b_x_32b(p0_TestBlock__A_op90, p0_TestBlock__B_op3);
  assign p1_smul_76345_comb = smul32b_32b_x_32b(p0_TestBlock__A_op91, p0_TestBlock__B_op13);
  assign p1_smul_76346_comb = smul32b_32b_x_32b(p0_TestBlock__A_op92, p0_TestBlock__B_op23);
  assign p1_smul_76347_comb = smul32b_32b_x_32b(p0_TestBlock__A_op93, p0_TestBlock__B_op33);
  assign p1_smul_76348_comb = smul32b_32b_x_32b(p0_TestBlock__A_op90, p0_TestBlock__B_op4);
  assign p1_smul_76349_comb = smul32b_32b_x_32b(p0_TestBlock__A_op91, p0_TestBlock__B_op14);
  assign p1_smul_76350_comb = smul32b_32b_x_32b(p0_TestBlock__A_op92, p0_TestBlock__B_op24);
  assign p1_smul_76351_comb = smul32b_32b_x_32b(p0_TestBlock__A_op93, p0_TestBlock__B_op34);
  assign p1_smul_76352_comb = smul32b_32b_x_32b(p0_TestBlock__A_op90, p0_TestBlock__B_op5);
  assign p1_smul_76353_comb = smul32b_32b_x_32b(p0_TestBlock__A_op91, p0_TestBlock__B_op15);
  assign p1_smul_76354_comb = smul32b_32b_x_32b(p0_TestBlock__A_op92, p0_TestBlock__B_op25);
  assign p1_smul_76355_comb = smul32b_32b_x_32b(p0_TestBlock__A_op93, p0_TestBlock__B_op35);
  assign p1_smul_76356_comb = smul32b_32b_x_32b(p0_TestBlock__A_op90, p0_TestBlock__B_op6);
  assign p1_smul_76357_comb = smul32b_32b_x_32b(p0_TestBlock__A_op91, p0_TestBlock__B_op16);
  assign p1_smul_76358_comb = smul32b_32b_x_32b(p0_TestBlock__A_op92, p0_TestBlock__B_op26);
  assign p1_smul_76359_comb = smul32b_32b_x_32b(p0_TestBlock__A_op93, p0_TestBlock__B_op36);
  assign p1_smul_76360_comb = smul32b_32b_x_32b(p0_TestBlock__A_op90, p0_TestBlock__B_op7);
  assign p1_smul_76361_comb = smul32b_32b_x_32b(p0_TestBlock__A_op91, p0_TestBlock__B_op17);
  assign p1_smul_76362_comb = smul32b_32b_x_32b(p0_TestBlock__A_op92, p0_TestBlock__B_op27);
  assign p1_smul_76363_comb = smul32b_32b_x_32b(p0_TestBlock__A_op93, p0_TestBlock__B_op37);
  assign p1_smul_76364_comb = smul32b_32b_x_32b(p0_TestBlock__A_op90, p0_TestBlock__B_op8);
  assign p1_smul_76365_comb = smul32b_32b_x_32b(p0_TestBlock__A_op91, p0_TestBlock__B_op18);
  assign p1_smul_76366_comb = smul32b_32b_x_32b(p0_TestBlock__A_op92, p0_TestBlock__B_op28);
  assign p1_smul_76367_comb = smul32b_32b_x_32b(p0_TestBlock__A_op93, p0_TestBlock__B_op38);
  assign p1_smul_76368_comb = smul32b_32b_x_32b(p0_TestBlock__A_op90, p0_TestBlock__B_op9);
  assign p1_smul_76369_comb = smul32b_32b_x_32b(p0_TestBlock__A_op91, p0_TestBlock__B_op19);
  assign p1_smul_76370_comb = smul32b_32b_x_32b(p0_TestBlock__A_op92, p0_TestBlock__B_op29);
  assign p1_smul_76371_comb = smul32b_32b_x_32b(p0_TestBlock__A_op93, p0_TestBlock__B_op39);
  assign p1_smul_76372_comb = smul32b_32b_x_32b(p0_TestBlock__A_op4, p0_TestBlock__B_op40);
  assign p1_smul_76373_comb = smul32b_32b_x_32b(p0_TestBlock__A_op5, p0_TestBlock__B_op50);
  assign p1_smul_76374_comb = smul32b_32b_x_32b(p0_TestBlock__A_op6, p0_TestBlock__B_op60);
  assign p1_smul_76375_comb = smul32b_32b_x_32b(p0_TestBlock__A_op7, p0_TestBlock__B_op70);
  assign p1_smul_76376_comb = smul32b_32b_x_32b(p0_TestBlock__A_op8, p0_TestBlock__B_op80);
  assign p1_smul_76377_comb = smul32b_32b_x_32b(p0_TestBlock__A_op9, p0_TestBlock__B_op90);
  assign p1_smul_76378_comb = smul32b_32b_x_32b(p0_TestBlock__A_op4, p0_TestBlock__B_op41);
  assign p1_smul_76379_comb = smul32b_32b_x_32b(p0_TestBlock__A_op5, p0_TestBlock__B_op51);
  assign p1_smul_76380_comb = smul32b_32b_x_32b(p0_TestBlock__A_op6, p0_TestBlock__B_op61);
  assign p1_smul_76381_comb = smul32b_32b_x_32b(p0_TestBlock__A_op7, p0_TestBlock__B_op71);
  assign p1_smul_76382_comb = smul32b_32b_x_32b(p0_TestBlock__A_op8, p0_TestBlock__B_op81);
  assign p1_smul_76383_comb = smul32b_32b_x_32b(p0_TestBlock__A_op9, p0_TestBlock__B_op91);
  assign p1_smul_76384_comb = smul32b_32b_x_32b(p0_TestBlock__A_op4, p0_TestBlock__B_op42);
  assign p1_smul_76385_comb = smul32b_32b_x_32b(p0_TestBlock__A_op5, p0_TestBlock__B_op52);
  assign p1_smul_76386_comb = smul32b_32b_x_32b(p0_TestBlock__A_op6, p0_TestBlock__B_op62);
  assign p1_smul_76387_comb = smul32b_32b_x_32b(p0_TestBlock__A_op7, p0_TestBlock__B_op72);
  assign p1_smul_76388_comb = smul32b_32b_x_32b(p0_TestBlock__A_op8, p0_TestBlock__B_op82);
  assign p1_smul_76389_comb = smul32b_32b_x_32b(p0_TestBlock__A_op9, p0_TestBlock__B_op92);
  assign p1_smul_76390_comb = smul32b_32b_x_32b(p0_TestBlock__A_op4, p0_TestBlock__B_op43);
  assign p1_smul_76391_comb = smul32b_32b_x_32b(p0_TestBlock__A_op5, p0_TestBlock__B_op53);
  assign p1_smul_76392_comb = smul32b_32b_x_32b(p0_TestBlock__A_op6, p0_TestBlock__B_op63);
  assign p1_smul_76393_comb = smul32b_32b_x_32b(p0_TestBlock__A_op7, p0_TestBlock__B_op73);
  assign p1_smul_76394_comb = smul32b_32b_x_32b(p0_TestBlock__A_op8, p0_TestBlock__B_op83);
  assign p1_smul_76395_comb = smul32b_32b_x_32b(p0_TestBlock__A_op9, p0_TestBlock__B_op93);
  assign p1_smul_76396_comb = smul32b_32b_x_32b(p0_TestBlock__A_op4, p0_TestBlock__B_op44);
  assign p1_smul_76397_comb = smul32b_32b_x_32b(p0_TestBlock__A_op5, p0_TestBlock__B_op54);
  assign p1_smul_76398_comb = smul32b_32b_x_32b(p0_TestBlock__A_op6, p0_TestBlock__B_op64);
  assign p1_smul_76399_comb = smul32b_32b_x_32b(p0_TestBlock__A_op7, p0_TestBlock__B_op74);
  assign p1_smul_76400_comb = smul32b_32b_x_32b(p0_TestBlock__A_op8, p0_TestBlock__B_op84);
  assign p1_smul_76401_comb = smul32b_32b_x_32b(p0_TestBlock__A_op9, p0_TestBlock__B_op94);
  assign p1_smul_76402_comb = smul32b_32b_x_32b(p0_TestBlock__A_op4, p0_TestBlock__B_op45);
  assign p1_smul_76403_comb = smul32b_32b_x_32b(p0_TestBlock__A_op5, p0_TestBlock__B_op55);
  assign p1_smul_76404_comb = smul32b_32b_x_32b(p0_TestBlock__A_op6, p0_TestBlock__B_op65);
  assign p1_smul_76405_comb = smul32b_32b_x_32b(p0_TestBlock__A_op7, p0_TestBlock__B_op75);
  assign p1_smul_76406_comb = smul32b_32b_x_32b(p0_TestBlock__A_op8, p0_TestBlock__B_op85);
  assign p1_smul_76407_comb = smul32b_32b_x_32b(p0_TestBlock__A_op9, p0_TestBlock__B_op95);
  assign p1_smul_76408_comb = smul32b_32b_x_32b(p0_TestBlock__A_op4, p0_TestBlock__B_op46);
  assign p1_smul_76409_comb = smul32b_32b_x_32b(p0_TestBlock__A_op5, p0_TestBlock__B_op56);
  assign p1_smul_76410_comb = smul32b_32b_x_32b(p0_TestBlock__A_op6, p0_TestBlock__B_op66);
  assign p1_smul_76411_comb = smul32b_32b_x_32b(p0_TestBlock__A_op7, p0_TestBlock__B_op76);
  assign p1_smul_76412_comb = smul32b_32b_x_32b(p0_TestBlock__A_op8, p0_TestBlock__B_op86);
  assign p1_smul_76413_comb = smul32b_32b_x_32b(p0_TestBlock__A_op9, p0_TestBlock__B_op96);
  assign p1_smul_76414_comb = smul32b_32b_x_32b(p0_TestBlock__A_op4, p0_TestBlock__B_op47);
  assign p1_smul_76415_comb = smul32b_32b_x_32b(p0_TestBlock__A_op5, p0_TestBlock__B_op57);
  assign p1_smul_76416_comb = smul32b_32b_x_32b(p0_TestBlock__A_op6, p0_TestBlock__B_op67);
  assign p1_smul_76417_comb = smul32b_32b_x_32b(p0_TestBlock__A_op7, p0_TestBlock__B_op77);
  assign p1_smul_76418_comb = smul32b_32b_x_32b(p0_TestBlock__A_op8, p0_TestBlock__B_op87);
  assign p1_smul_76419_comb = smul32b_32b_x_32b(p0_TestBlock__A_op9, p0_TestBlock__B_op97);
  assign p1_smul_76420_comb = smul32b_32b_x_32b(p0_TestBlock__A_op4, p0_TestBlock__B_op48);
  assign p1_smul_76421_comb = smul32b_32b_x_32b(p0_TestBlock__A_op5, p0_TestBlock__B_op58);
  assign p1_smul_76422_comb = smul32b_32b_x_32b(p0_TestBlock__A_op6, p0_TestBlock__B_op68);
  assign p1_smul_76423_comb = smul32b_32b_x_32b(p0_TestBlock__A_op7, p0_TestBlock__B_op78);
  assign p1_smul_76424_comb = smul32b_32b_x_32b(p0_TestBlock__A_op8, p0_TestBlock__B_op88);
  assign p1_smul_76425_comb = smul32b_32b_x_32b(p0_TestBlock__A_op9, p0_TestBlock__B_op98);
  assign p1_smul_76426_comb = smul32b_32b_x_32b(p0_TestBlock__A_op4, p0_TestBlock__B_op49);
  assign p1_smul_76427_comb = smul32b_32b_x_32b(p0_TestBlock__A_op5, p0_TestBlock__B_op59);
  assign p1_smul_76428_comb = smul32b_32b_x_32b(p0_TestBlock__A_op6, p0_TestBlock__B_op69);
  assign p1_smul_76429_comb = smul32b_32b_x_32b(p0_TestBlock__A_op7, p0_TestBlock__B_op79);
  assign p1_smul_76430_comb = smul32b_32b_x_32b(p0_TestBlock__A_op8, p0_TestBlock__B_op89);
  assign p1_smul_76431_comb = smul32b_32b_x_32b(p0_TestBlock__A_op9, p0_TestBlock__B_op99);
  assign p1_smul_76432_comb = smul32b_32b_x_32b(p0_TestBlock__A_op14, p0_TestBlock__B_op40);
  assign p1_smul_76433_comb = smul32b_32b_x_32b(p0_TestBlock__A_op15, p0_TestBlock__B_op50);
  assign p1_smul_76434_comb = smul32b_32b_x_32b(p0_TestBlock__A_op16, p0_TestBlock__B_op60);
  assign p1_smul_76435_comb = smul32b_32b_x_32b(p0_TestBlock__A_op17, p0_TestBlock__B_op70);
  assign p1_smul_76436_comb = smul32b_32b_x_32b(p0_TestBlock__A_op18, p0_TestBlock__B_op80);
  assign p1_smul_76437_comb = smul32b_32b_x_32b(p0_TestBlock__A_op19, p0_TestBlock__B_op90);
  assign p1_smul_76438_comb = smul32b_32b_x_32b(p0_TestBlock__A_op14, p0_TestBlock__B_op41);
  assign p1_smul_76439_comb = smul32b_32b_x_32b(p0_TestBlock__A_op15, p0_TestBlock__B_op51);
  assign p1_smul_76440_comb = smul32b_32b_x_32b(p0_TestBlock__A_op16, p0_TestBlock__B_op61);
  assign p1_smul_76441_comb = smul32b_32b_x_32b(p0_TestBlock__A_op17, p0_TestBlock__B_op71);
  assign p1_smul_76442_comb = smul32b_32b_x_32b(p0_TestBlock__A_op18, p0_TestBlock__B_op81);
  assign p1_smul_76443_comb = smul32b_32b_x_32b(p0_TestBlock__A_op19, p0_TestBlock__B_op91);
  assign p1_smul_76444_comb = smul32b_32b_x_32b(p0_TestBlock__A_op14, p0_TestBlock__B_op42);
  assign p1_smul_76445_comb = smul32b_32b_x_32b(p0_TestBlock__A_op15, p0_TestBlock__B_op52);
  assign p1_smul_76446_comb = smul32b_32b_x_32b(p0_TestBlock__A_op16, p0_TestBlock__B_op62);
  assign p1_smul_76447_comb = smul32b_32b_x_32b(p0_TestBlock__A_op17, p0_TestBlock__B_op72);
  assign p1_smul_76448_comb = smul32b_32b_x_32b(p0_TestBlock__A_op18, p0_TestBlock__B_op82);
  assign p1_smul_76449_comb = smul32b_32b_x_32b(p0_TestBlock__A_op19, p0_TestBlock__B_op92);
  assign p1_smul_76450_comb = smul32b_32b_x_32b(p0_TestBlock__A_op14, p0_TestBlock__B_op43);
  assign p1_smul_76451_comb = smul32b_32b_x_32b(p0_TestBlock__A_op15, p0_TestBlock__B_op53);
  assign p1_smul_76452_comb = smul32b_32b_x_32b(p0_TestBlock__A_op16, p0_TestBlock__B_op63);
  assign p1_smul_76453_comb = smul32b_32b_x_32b(p0_TestBlock__A_op17, p0_TestBlock__B_op73);
  assign p1_smul_76454_comb = smul32b_32b_x_32b(p0_TestBlock__A_op18, p0_TestBlock__B_op83);
  assign p1_smul_76455_comb = smul32b_32b_x_32b(p0_TestBlock__A_op19, p0_TestBlock__B_op93);
  assign p1_smul_76456_comb = smul32b_32b_x_32b(p0_TestBlock__A_op14, p0_TestBlock__B_op44);
  assign p1_smul_76457_comb = smul32b_32b_x_32b(p0_TestBlock__A_op15, p0_TestBlock__B_op54);
  assign p1_smul_76458_comb = smul32b_32b_x_32b(p0_TestBlock__A_op16, p0_TestBlock__B_op64);
  assign p1_smul_76459_comb = smul32b_32b_x_32b(p0_TestBlock__A_op17, p0_TestBlock__B_op74);
  assign p1_smul_76460_comb = smul32b_32b_x_32b(p0_TestBlock__A_op18, p0_TestBlock__B_op84);
  assign p1_smul_76461_comb = smul32b_32b_x_32b(p0_TestBlock__A_op19, p0_TestBlock__B_op94);
  assign p1_smul_76462_comb = smul32b_32b_x_32b(p0_TestBlock__A_op14, p0_TestBlock__B_op45);
  assign p1_smul_76463_comb = smul32b_32b_x_32b(p0_TestBlock__A_op15, p0_TestBlock__B_op55);
  assign p1_smul_76464_comb = smul32b_32b_x_32b(p0_TestBlock__A_op16, p0_TestBlock__B_op65);
  assign p1_smul_76465_comb = smul32b_32b_x_32b(p0_TestBlock__A_op17, p0_TestBlock__B_op75);
  assign p1_smul_76466_comb = smul32b_32b_x_32b(p0_TestBlock__A_op18, p0_TestBlock__B_op85);
  assign p1_smul_76467_comb = smul32b_32b_x_32b(p0_TestBlock__A_op19, p0_TestBlock__B_op95);
  assign p1_smul_76468_comb = smul32b_32b_x_32b(p0_TestBlock__A_op14, p0_TestBlock__B_op46);
  assign p1_smul_76469_comb = smul32b_32b_x_32b(p0_TestBlock__A_op15, p0_TestBlock__B_op56);
  assign p1_smul_76470_comb = smul32b_32b_x_32b(p0_TestBlock__A_op16, p0_TestBlock__B_op66);
  assign p1_smul_76471_comb = smul32b_32b_x_32b(p0_TestBlock__A_op17, p0_TestBlock__B_op76);
  assign p1_smul_76472_comb = smul32b_32b_x_32b(p0_TestBlock__A_op18, p0_TestBlock__B_op86);
  assign p1_smul_76473_comb = smul32b_32b_x_32b(p0_TestBlock__A_op19, p0_TestBlock__B_op96);
  assign p1_smul_76474_comb = smul32b_32b_x_32b(p0_TestBlock__A_op14, p0_TestBlock__B_op47);
  assign p1_smul_76475_comb = smul32b_32b_x_32b(p0_TestBlock__A_op15, p0_TestBlock__B_op57);
  assign p1_smul_76476_comb = smul32b_32b_x_32b(p0_TestBlock__A_op16, p0_TestBlock__B_op67);
  assign p1_smul_76477_comb = smul32b_32b_x_32b(p0_TestBlock__A_op17, p0_TestBlock__B_op77);
  assign p1_smul_76478_comb = smul32b_32b_x_32b(p0_TestBlock__A_op18, p0_TestBlock__B_op87);
  assign p1_smul_76479_comb = smul32b_32b_x_32b(p0_TestBlock__A_op19, p0_TestBlock__B_op97);
  assign p1_smul_76480_comb = smul32b_32b_x_32b(p0_TestBlock__A_op14, p0_TestBlock__B_op48);
  assign p1_smul_76481_comb = smul32b_32b_x_32b(p0_TestBlock__A_op15, p0_TestBlock__B_op58);
  assign p1_smul_76482_comb = smul32b_32b_x_32b(p0_TestBlock__A_op16, p0_TestBlock__B_op68);
  assign p1_smul_76483_comb = smul32b_32b_x_32b(p0_TestBlock__A_op17, p0_TestBlock__B_op78);
  assign p1_smul_76484_comb = smul32b_32b_x_32b(p0_TestBlock__A_op18, p0_TestBlock__B_op88);
  assign p1_smul_76485_comb = smul32b_32b_x_32b(p0_TestBlock__A_op19, p0_TestBlock__B_op98);
  assign p1_smul_76486_comb = smul32b_32b_x_32b(p0_TestBlock__A_op14, p0_TestBlock__B_op49);
  assign p1_smul_76487_comb = smul32b_32b_x_32b(p0_TestBlock__A_op15, p0_TestBlock__B_op59);
  assign p1_smul_76488_comb = smul32b_32b_x_32b(p0_TestBlock__A_op16, p0_TestBlock__B_op69);
  assign p1_smul_76489_comb = smul32b_32b_x_32b(p0_TestBlock__A_op17, p0_TestBlock__B_op79);
  assign p1_smul_76490_comb = smul32b_32b_x_32b(p0_TestBlock__A_op18, p0_TestBlock__B_op89);
  assign p1_smul_76491_comb = smul32b_32b_x_32b(p0_TestBlock__A_op19, p0_TestBlock__B_op99);
  assign p1_smul_76492_comb = smul32b_32b_x_32b(p0_TestBlock__A_op24, p0_TestBlock__B_op40);
  assign p1_smul_76493_comb = smul32b_32b_x_32b(p0_TestBlock__A_op25, p0_TestBlock__B_op50);
  assign p1_smul_76494_comb = smul32b_32b_x_32b(p0_TestBlock__A_op26, p0_TestBlock__B_op60);
  assign p1_smul_76495_comb = smul32b_32b_x_32b(p0_TestBlock__A_op27, p0_TestBlock__B_op70);
  assign p1_smul_76496_comb = smul32b_32b_x_32b(p0_TestBlock__A_op28, p0_TestBlock__B_op80);
  assign p1_smul_76497_comb = smul32b_32b_x_32b(p0_TestBlock__A_op29, p0_TestBlock__B_op90);
  assign p1_smul_76498_comb = smul32b_32b_x_32b(p0_TestBlock__A_op24, p0_TestBlock__B_op41);
  assign p1_smul_76499_comb = smul32b_32b_x_32b(p0_TestBlock__A_op25, p0_TestBlock__B_op51);
  assign p1_smul_76500_comb = smul32b_32b_x_32b(p0_TestBlock__A_op26, p0_TestBlock__B_op61);
  assign p1_smul_76501_comb = smul32b_32b_x_32b(p0_TestBlock__A_op27, p0_TestBlock__B_op71);
  assign p1_smul_76502_comb = smul32b_32b_x_32b(p0_TestBlock__A_op28, p0_TestBlock__B_op81);
  assign p1_smul_76503_comb = smul32b_32b_x_32b(p0_TestBlock__A_op29, p0_TestBlock__B_op91);
  assign p1_smul_76504_comb = smul32b_32b_x_32b(p0_TestBlock__A_op24, p0_TestBlock__B_op42);
  assign p1_smul_76505_comb = smul32b_32b_x_32b(p0_TestBlock__A_op25, p0_TestBlock__B_op52);
  assign p1_smul_76506_comb = smul32b_32b_x_32b(p0_TestBlock__A_op26, p0_TestBlock__B_op62);
  assign p1_smul_76507_comb = smul32b_32b_x_32b(p0_TestBlock__A_op27, p0_TestBlock__B_op72);
  assign p1_smul_76508_comb = smul32b_32b_x_32b(p0_TestBlock__A_op28, p0_TestBlock__B_op82);
  assign p1_smul_76509_comb = smul32b_32b_x_32b(p0_TestBlock__A_op29, p0_TestBlock__B_op92);
  assign p1_smul_76510_comb = smul32b_32b_x_32b(p0_TestBlock__A_op24, p0_TestBlock__B_op43);
  assign p1_smul_76511_comb = smul32b_32b_x_32b(p0_TestBlock__A_op25, p0_TestBlock__B_op53);
  assign p1_smul_76512_comb = smul32b_32b_x_32b(p0_TestBlock__A_op26, p0_TestBlock__B_op63);
  assign p1_smul_76513_comb = smul32b_32b_x_32b(p0_TestBlock__A_op27, p0_TestBlock__B_op73);
  assign p1_smul_76514_comb = smul32b_32b_x_32b(p0_TestBlock__A_op28, p0_TestBlock__B_op83);
  assign p1_smul_76515_comb = smul32b_32b_x_32b(p0_TestBlock__A_op29, p0_TestBlock__B_op93);
  assign p1_smul_76516_comb = smul32b_32b_x_32b(p0_TestBlock__A_op24, p0_TestBlock__B_op44);
  assign p1_smul_76517_comb = smul32b_32b_x_32b(p0_TestBlock__A_op25, p0_TestBlock__B_op54);
  assign p1_smul_76518_comb = smul32b_32b_x_32b(p0_TestBlock__A_op26, p0_TestBlock__B_op64);
  assign p1_smul_76519_comb = smul32b_32b_x_32b(p0_TestBlock__A_op27, p0_TestBlock__B_op74);
  assign p1_smul_76520_comb = smul32b_32b_x_32b(p0_TestBlock__A_op28, p0_TestBlock__B_op84);
  assign p1_smul_76521_comb = smul32b_32b_x_32b(p0_TestBlock__A_op29, p0_TestBlock__B_op94);
  assign p1_smul_76522_comb = smul32b_32b_x_32b(p0_TestBlock__A_op24, p0_TestBlock__B_op45);
  assign p1_smul_76523_comb = smul32b_32b_x_32b(p0_TestBlock__A_op25, p0_TestBlock__B_op55);
  assign p1_smul_76524_comb = smul32b_32b_x_32b(p0_TestBlock__A_op26, p0_TestBlock__B_op65);
  assign p1_smul_76525_comb = smul32b_32b_x_32b(p0_TestBlock__A_op27, p0_TestBlock__B_op75);
  assign p1_smul_76526_comb = smul32b_32b_x_32b(p0_TestBlock__A_op28, p0_TestBlock__B_op85);
  assign p1_smul_76527_comb = smul32b_32b_x_32b(p0_TestBlock__A_op29, p0_TestBlock__B_op95);
  assign p1_smul_76528_comb = smul32b_32b_x_32b(p0_TestBlock__A_op24, p0_TestBlock__B_op46);
  assign p1_smul_76529_comb = smul32b_32b_x_32b(p0_TestBlock__A_op25, p0_TestBlock__B_op56);
  assign p1_smul_76530_comb = smul32b_32b_x_32b(p0_TestBlock__A_op26, p0_TestBlock__B_op66);
  assign p1_smul_76531_comb = smul32b_32b_x_32b(p0_TestBlock__A_op27, p0_TestBlock__B_op76);
  assign p1_smul_76532_comb = smul32b_32b_x_32b(p0_TestBlock__A_op28, p0_TestBlock__B_op86);
  assign p1_smul_76533_comb = smul32b_32b_x_32b(p0_TestBlock__A_op29, p0_TestBlock__B_op96);
  assign p1_smul_76534_comb = smul32b_32b_x_32b(p0_TestBlock__A_op24, p0_TestBlock__B_op47);
  assign p1_smul_76535_comb = smul32b_32b_x_32b(p0_TestBlock__A_op25, p0_TestBlock__B_op57);
  assign p1_smul_76536_comb = smul32b_32b_x_32b(p0_TestBlock__A_op26, p0_TestBlock__B_op67);
  assign p1_smul_76537_comb = smul32b_32b_x_32b(p0_TestBlock__A_op27, p0_TestBlock__B_op77);
  assign p1_smul_76538_comb = smul32b_32b_x_32b(p0_TestBlock__A_op28, p0_TestBlock__B_op87);
  assign p1_smul_76539_comb = smul32b_32b_x_32b(p0_TestBlock__A_op29, p0_TestBlock__B_op97);
  assign p1_smul_76540_comb = smul32b_32b_x_32b(p0_TestBlock__A_op24, p0_TestBlock__B_op48);
  assign p1_smul_76541_comb = smul32b_32b_x_32b(p0_TestBlock__A_op25, p0_TestBlock__B_op58);
  assign p1_smul_76542_comb = smul32b_32b_x_32b(p0_TestBlock__A_op26, p0_TestBlock__B_op68);
  assign p1_smul_76543_comb = smul32b_32b_x_32b(p0_TestBlock__A_op27, p0_TestBlock__B_op78);
  assign p1_smul_76544_comb = smul32b_32b_x_32b(p0_TestBlock__A_op28, p0_TestBlock__B_op88);
  assign p1_smul_76545_comb = smul32b_32b_x_32b(p0_TestBlock__A_op29, p0_TestBlock__B_op98);
  assign p1_smul_76546_comb = smul32b_32b_x_32b(p0_TestBlock__A_op24, p0_TestBlock__B_op49);
  assign p1_smul_76547_comb = smul32b_32b_x_32b(p0_TestBlock__A_op25, p0_TestBlock__B_op59);
  assign p1_smul_76548_comb = smul32b_32b_x_32b(p0_TestBlock__A_op26, p0_TestBlock__B_op69);
  assign p1_smul_76549_comb = smul32b_32b_x_32b(p0_TestBlock__A_op27, p0_TestBlock__B_op79);
  assign p1_smul_76550_comb = smul32b_32b_x_32b(p0_TestBlock__A_op28, p0_TestBlock__B_op89);
  assign p1_smul_76551_comb = smul32b_32b_x_32b(p0_TestBlock__A_op29, p0_TestBlock__B_op99);
  assign p1_smul_76552_comb = smul32b_32b_x_32b(p0_TestBlock__A_op34, p0_TestBlock__B_op40);
  assign p1_smul_76553_comb = smul32b_32b_x_32b(p0_TestBlock__A_op35, p0_TestBlock__B_op50);
  assign p1_smul_76554_comb = smul32b_32b_x_32b(p0_TestBlock__A_op36, p0_TestBlock__B_op60);
  assign p1_smul_76555_comb = smul32b_32b_x_32b(p0_TestBlock__A_op37, p0_TestBlock__B_op70);
  assign p1_smul_76556_comb = smul32b_32b_x_32b(p0_TestBlock__A_op38, p0_TestBlock__B_op80);
  assign p1_smul_76557_comb = smul32b_32b_x_32b(p0_TestBlock__A_op39, p0_TestBlock__B_op90);
  assign p1_smul_76558_comb = smul32b_32b_x_32b(p0_TestBlock__A_op34, p0_TestBlock__B_op41);
  assign p1_smul_76559_comb = smul32b_32b_x_32b(p0_TestBlock__A_op35, p0_TestBlock__B_op51);
  assign p1_smul_76560_comb = smul32b_32b_x_32b(p0_TestBlock__A_op36, p0_TestBlock__B_op61);
  assign p1_smul_76561_comb = smul32b_32b_x_32b(p0_TestBlock__A_op37, p0_TestBlock__B_op71);
  assign p1_smul_76562_comb = smul32b_32b_x_32b(p0_TestBlock__A_op38, p0_TestBlock__B_op81);
  assign p1_smul_76563_comb = smul32b_32b_x_32b(p0_TestBlock__A_op39, p0_TestBlock__B_op91);
  assign p1_smul_76564_comb = smul32b_32b_x_32b(p0_TestBlock__A_op34, p0_TestBlock__B_op42);
  assign p1_smul_76565_comb = smul32b_32b_x_32b(p0_TestBlock__A_op35, p0_TestBlock__B_op52);
  assign p1_smul_76566_comb = smul32b_32b_x_32b(p0_TestBlock__A_op36, p0_TestBlock__B_op62);
  assign p1_smul_76567_comb = smul32b_32b_x_32b(p0_TestBlock__A_op37, p0_TestBlock__B_op72);
  assign p1_smul_76568_comb = smul32b_32b_x_32b(p0_TestBlock__A_op38, p0_TestBlock__B_op82);
  assign p1_smul_76569_comb = smul32b_32b_x_32b(p0_TestBlock__A_op39, p0_TestBlock__B_op92);
  assign p1_smul_76570_comb = smul32b_32b_x_32b(p0_TestBlock__A_op34, p0_TestBlock__B_op43);
  assign p1_smul_76571_comb = smul32b_32b_x_32b(p0_TestBlock__A_op35, p0_TestBlock__B_op53);
  assign p1_smul_76572_comb = smul32b_32b_x_32b(p0_TestBlock__A_op36, p0_TestBlock__B_op63);
  assign p1_smul_76573_comb = smul32b_32b_x_32b(p0_TestBlock__A_op37, p0_TestBlock__B_op73);
  assign p1_smul_76574_comb = smul32b_32b_x_32b(p0_TestBlock__A_op38, p0_TestBlock__B_op83);
  assign p1_smul_76575_comb = smul32b_32b_x_32b(p0_TestBlock__A_op39, p0_TestBlock__B_op93);
  assign p1_smul_76576_comb = smul32b_32b_x_32b(p0_TestBlock__A_op34, p0_TestBlock__B_op44);
  assign p1_smul_76577_comb = smul32b_32b_x_32b(p0_TestBlock__A_op35, p0_TestBlock__B_op54);
  assign p1_smul_76578_comb = smul32b_32b_x_32b(p0_TestBlock__A_op36, p0_TestBlock__B_op64);
  assign p1_smul_76579_comb = smul32b_32b_x_32b(p0_TestBlock__A_op37, p0_TestBlock__B_op74);
  assign p1_smul_76580_comb = smul32b_32b_x_32b(p0_TestBlock__A_op38, p0_TestBlock__B_op84);
  assign p1_smul_76581_comb = smul32b_32b_x_32b(p0_TestBlock__A_op39, p0_TestBlock__B_op94);
  assign p1_smul_76582_comb = smul32b_32b_x_32b(p0_TestBlock__A_op34, p0_TestBlock__B_op45);
  assign p1_smul_76583_comb = smul32b_32b_x_32b(p0_TestBlock__A_op35, p0_TestBlock__B_op55);
  assign p1_smul_76584_comb = smul32b_32b_x_32b(p0_TestBlock__A_op36, p0_TestBlock__B_op65);
  assign p1_smul_76585_comb = smul32b_32b_x_32b(p0_TestBlock__A_op37, p0_TestBlock__B_op75);
  assign p1_smul_76586_comb = smul32b_32b_x_32b(p0_TestBlock__A_op38, p0_TestBlock__B_op85);
  assign p1_smul_76587_comb = smul32b_32b_x_32b(p0_TestBlock__A_op39, p0_TestBlock__B_op95);
  assign p1_smul_76588_comb = smul32b_32b_x_32b(p0_TestBlock__A_op34, p0_TestBlock__B_op46);
  assign p1_smul_76589_comb = smul32b_32b_x_32b(p0_TestBlock__A_op35, p0_TestBlock__B_op56);
  assign p1_smul_76590_comb = smul32b_32b_x_32b(p0_TestBlock__A_op36, p0_TestBlock__B_op66);
  assign p1_smul_76591_comb = smul32b_32b_x_32b(p0_TestBlock__A_op37, p0_TestBlock__B_op76);
  assign p1_smul_76592_comb = smul32b_32b_x_32b(p0_TestBlock__A_op38, p0_TestBlock__B_op86);
  assign p1_smul_76593_comb = smul32b_32b_x_32b(p0_TestBlock__A_op39, p0_TestBlock__B_op96);
  assign p1_smul_76594_comb = smul32b_32b_x_32b(p0_TestBlock__A_op34, p0_TestBlock__B_op47);
  assign p1_smul_76595_comb = smul32b_32b_x_32b(p0_TestBlock__A_op35, p0_TestBlock__B_op57);
  assign p1_smul_76596_comb = smul32b_32b_x_32b(p0_TestBlock__A_op36, p0_TestBlock__B_op67);
  assign p1_smul_76597_comb = smul32b_32b_x_32b(p0_TestBlock__A_op37, p0_TestBlock__B_op77);
  assign p1_smul_76598_comb = smul32b_32b_x_32b(p0_TestBlock__A_op38, p0_TestBlock__B_op87);
  assign p1_smul_76599_comb = smul32b_32b_x_32b(p0_TestBlock__A_op39, p0_TestBlock__B_op97);
  assign p1_smul_76600_comb = smul32b_32b_x_32b(p0_TestBlock__A_op34, p0_TestBlock__B_op48);
  assign p1_smul_76601_comb = smul32b_32b_x_32b(p0_TestBlock__A_op35, p0_TestBlock__B_op58);
  assign p1_smul_76602_comb = smul32b_32b_x_32b(p0_TestBlock__A_op36, p0_TestBlock__B_op68);
  assign p1_smul_76603_comb = smul32b_32b_x_32b(p0_TestBlock__A_op37, p0_TestBlock__B_op78);
  assign p1_smul_76604_comb = smul32b_32b_x_32b(p0_TestBlock__A_op38, p0_TestBlock__B_op88);
  assign p1_smul_76605_comb = smul32b_32b_x_32b(p0_TestBlock__A_op39, p0_TestBlock__B_op98);
  assign p1_smul_76606_comb = smul32b_32b_x_32b(p0_TestBlock__A_op34, p0_TestBlock__B_op49);
  assign p1_smul_76607_comb = smul32b_32b_x_32b(p0_TestBlock__A_op35, p0_TestBlock__B_op59);
  assign p1_smul_76608_comb = smul32b_32b_x_32b(p0_TestBlock__A_op36, p0_TestBlock__B_op69);
  assign p1_smul_76609_comb = smul32b_32b_x_32b(p0_TestBlock__A_op37, p0_TestBlock__B_op79);
  assign p1_smul_76610_comb = smul32b_32b_x_32b(p0_TestBlock__A_op38, p0_TestBlock__B_op89);
  assign p1_smul_76611_comb = smul32b_32b_x_32b(p0_TestBlock__A_op39, p0_TestBlock__B_op99);
  assign p1_smul_76612_comb = smul32b_32b_x_32b(p0_TestBlock__A_op44, p0_TestBlock__B_op40);
  assign p1_smul_76613_comb = smul32b_32b_x_32b(p0_TestBlock__A_op45, p0_TestBlock__B_op50);
  assign p1_smul_76614_comb = smul32b_32b_x_32b(p0_TestBlock__A_op46, p0_TestBlock__B_op60);
  assign p1_smul_76615_comb = smul32b_32b_x_32b(p0_TestBlock__A_op47, p0_TestBlock__B_op70);
  assign p1_smul_76616_comb = smul32b_32b_x_32b(p0_TestBlock__A_op48, p0_TestBlock__B_op80);
  assign p1_smul_76617_comb = smul32b_32b_x_32b(p0_TestBlock__A_op49, p0_TestBlock__B_op90);
  assign p1_smul_76618_comb = smul32b_32b_x_32b(p0_TestBlock__A_op44, p0_TestBlock__B_op41);
  assign p1_smul_76619_comb = smul32b_32b_x_32b(p0_TestBlock__A_op45, p0_TestBlock__B_op51);
  assign p1_smul_76620_comb = smul32b_32b_x_32b(p0_TestBlock__A_op46, p0_TestBlock__B_op61);
  assign p1_smul_76621_comb = smul32b_32b_x_32b(p0_TestBlock__A_op47, p0_TestBlock__B_op71);
  assign p1_smul_76622_comb = smul32b_32b_x_32b(p0_TestBlock__A_op48, p0_TestBlock__B_op81);
  assign p1_smul_76623_comb = smul32b_32b_x_32b(p0_TestBlock__A_op49, p0_TestBlock__B_op91);
  assign p1_smul_76624_comb = smul32b_32b_x_32b(p0_TestBlock__A_op44, p0_TestBlock__B_op42);
  assign p1_smul_76625_comb = smul32b_32b_x_32b(p0_TestBlock__A_op45, p0_TestBlock__B_op52);
  assign p1_smul_76626_comb = smul32b_32b_x_32b(p0_TestBlock__A_op46, p0_TestBlock__B_op62);
  assign p1_smul_76627_comb = smul32b_32b_x_32b(p0_TestBlock__A_op47, p0_TestBlock__B_op72);
  assign p1_smul_76628_comb = smul32b_32b_x_32b(p0_TestBlock__A_op48, p0_TestBlock__B_op82);
  assign p1_smul_76629_comb = smul32b_32b_x_32b(p0_TestBlock__A_op49, p0_TestBlock__B_op92);
  assign p1_smul_76630_comb = smul32b_32b_x_32b(p0_TestBlock__A_op44, p0_TestBlock__B_op43);
  assign p1_smul_76631_comb = smul32b_32b_x_32b(p0_TestBlock__A_op45, p0_TestBlock__B_op53);
  assign p1_smul_76632_comb = smul32b_32b_x_32b(p0_TestBlock__A_op46, p0_TestBlock__B_op63);
  assign p1_smul_76633_comb = smul32b_32b_x_32b(p0_TestBlock__A_op47, p0_TestBlock__B_op73);
  assign p1_smul_76634_comb = smul32b_32b_x_32b(p0_TestBlock__A_op48, p0_TestBlock__B_op83);
  assign p1_smul_76635_comb = smul32b_32b_x_32b(p0_TestBlock__A_op49, p0_TestBlock__B_op93);
  assign p1_smul_76636_comb = smul32b_32b_x_32b(p0_TestBlock__A_op44, p0_TestBlock__B_op44);
  assign p1_smul_76637_comb = smul32b_32b_x_32b(p0_TestBlock__A_op45, p0_TestBlock__B_op54);
  assign p1_smul_76638_comb = smul32b_32b_x_32b(p0_TestBlock__A_op46, p0_TestBlock__B_op64);
  assign p1_smul_76639_comb = smul32b_32b_x_32b(p0_TestBlock__A_op47, p0_TestBlock__B_op74);
  assign p1_smul_76640_comb = smul32b_32b_x_32b(p0_TestBlock__A_op48, p0_TestBlock__B_op84);
  assign p1_smul_76641_comb = smul32b_32b_x_32b(p0_TestBlock__A_op49, p0_TestBlock__B_op94);
  assign p1_smul_76642_comb = smul32b_32b_x_32b(p0_TestBlock__A_op44, p0_TestBlock__B_op45);
  assign p1_smul_76643_comb = smul32b_32b_x_32b(p0_TestBlock__A_op45, p0_TestBlock__B_op55);
  assign p1_smul_76644_comb = smul32b_32b_x_32b(p0_TestBlock__A_op46, p0_TestBlock__B_op65);
  assign p1_smul_76645_comb = smul32b_32b_x_32b(p0_TestBlock__A_op47, p0_TestBlock__B_op75);
  assign p1_smul_76646_comb = smul32b_32b_x_32b(p0_TestBlock__A_op48, p0_TestBlock__B_op85);
  assign p1_smul_76647_comb = smul32b_32b_x_32b(p0_TestBlock__A_op49, p0_TestBlock__B_op95);
  assign p1_smul_76648_comb = smul32b_32b_x_32b(p0_TestBlock__A_op44, p0_TestBlock__B_op46);
  assign p1_smul_76649_comb = smul32b_32b_x_32b(p0_TestBlock__A_op45, p0_TestBlock__B_op56);
  assign p1_smul_76650_comb = smul32b_32b_x_32b(p0_TestBlock__A_op46, p0_TestBlock__B_op66);
  assign p1_smul_76651_comb = smul32b_32b_x_32b(p0_TestBlock__A_op47, p0_TestBlock__B_op76);
  assign p1_smul_76652_comb = smul32b_32b_x_32b(p0_TestBlock__A_op48, p0_TestBlock__B_op86);
  assign p1_smul_76653_comb = smul32b_32b_x_32b(p0_TestBlock__A_op49, p0_TestBlock__B_op96);
  assign p1_smul_76654_comb = smul32b_32b_x_32b(p0_TestBlock__A_op44, p0_TestBlock__B_op47);
  assign p1_smul_76655_comb = smul32b_32b_x_32b(p0_TestBlock__A_op45, p0_TestBlock__B_op57);
  assign p1_smul_76656_comb = smul32b_32b_x_32b(p0_TestBlock__A_op46, p0_TestBlock__B_op67);
  assign p1_smul_76657_comb = smul32b_32b_x_32b(p0_TestBlock__A_op47, p0_TestBlock__B_op77);
  assign p1_smul_76658_comb = smul32b_32b_x_32b(p0_TestBlock__A_op48, p0_TestBlock__B_op87);
  assign p1_smul_76659_comb = smul32b_32b_x_32b(p0_TestBlock__A_op49, p0_TestBlock__B_op97);
  assign p1_smul_76660_comb = smul32b_32b_x_32b(p0_TestBlock__A_op44, p0_TestBlock__B_op48);
  assign p1_smul_76661_comb = smul32b_32b_x_32b(p0_TestBlock__A_op45, p0_TestBlock__B_op58);
  assign p1_smul_76662_comb = smul32b_32b_x_32b(p0_TestBlock__A_op46, p0_TestBlock__B_op68);
  assign p1_smul_76663_comb = smul32b_32b_x_32b(p0_TestBlock__A_op47, p0_TestBlock__B_op78);
  assign p1_smul_76664_comb = smul32b_32b_x_32b(p0_TestBlock__A_op48, p0_TestBlock__B_op88);
  assign p1_smul_76665_comb = smul32b_32b_x_32b(p0_TestBlock__A_op49, p0_TestBlock__B_op98);
  assign p1_smul_76666_comb = smul32b_32b_x_32b(p0_TestBlock__A_op44, p0_TestBlock__B_op49);
  assign p1_smul_76667_comb = smul32b_32b_x_32b(p0_TestBlock__A_op45, p0_TestBlock__B_op59);
  assign p1_smul_76668_comb = smul32b_32b_x_32b(p0_TestBlock__A_op46, p0_TestBlock__B_op69);
  assign p1_smul_76669_comb = smul32b_32b_x_32b(p0_TestBlock__A_op47, p0_TestBlock__B_op79);
  assign p1_smul_76670_comb = smul32b_32b_x_32b(p0_TestBlock__A_op48, p0_TestBlock__B_op89);
  assign p1_smul_76671_comb = smul32b_32b_x_32b(p0_TestBlock__A_op49, p0_TestBlock__B_op99);
  assign p1_smul_76672_comb = smul32b_32b_x_32b(p0_TestBlock__A_op54, p0_TestBlock__B_op40);
  assign p1_smul_76673_comb = smul32b_32b_x_32b(p0_TestBlock__A_op55, p0_TestBlock__B_op50);
  assign p1_smul_76674_comb = smul32b_32b_x_32b(p0_TestBlock__A_op56, p0_TestBlock__B_op60);
  assign p1_smul_76675_comb = smul32b_32b_x_32b(p0_TestBlock__A_op57, p0_TestBlock__B_op70);
  assign p1_smul_76676_comb = smul32b_32b_x_32b(p0_TestBlock__A_op58, p0_TestBlock__B_op80);
  assign p1_smul_76677_comb = smul32b_32b_x_32b(p0_TestBlock__A_op59, p0_TestBlock__B_op90);
  assign p1_smul_76678_comb = smul32b_32b_x_32b(p0_TestBlock__A_op54, p0_TestBlock__B_op41);
  assign p1_smul_76679_comb = smul32b_32b_x_32b(p0_TestBlock__A_op55, p0_TestBlock__B_op51);
  assign p1_smul_76680_comb = smul32b_32b_x_32b(p0_TestBlock__A_op56, p0_TestBlock__B_op61);
  assign p1_smul_76681_comb = smul32b_32b_x_32b(p0_TestBlock__A_op57, p0_TestBlock__B_op71);
  assign p1_smul_76682_comb = smul32b_32b_x_32b(p0_TestBlock__A_op58, p0_TestBlock__B_op81);
  assign p1_smul_76683_comb = smul32b_32b_x_32b(p0_TestBlock__A_op59, p0_TestBlock__B_op91);
  assign p1_smul_76684_comb = smul32b_32b_x_32b(p0_TestBlock__A_op54, p0_TestBlock__B_op42);
  assign p1_smul_76685_comb = smul32b_32b_x_32b(p0_TestBlock__A_op55, p0_TestBlock__B_op52);
  assign p1_smul_76686_comb = smul32b_32b_x_32b(p0_TestBlock__A_op56, p0_TestBlock__B_op62);
  assign p1_smul_76687_comb = smul32b_32b_x_32b(p0_TestBlock__A_op57, p0_TestBlock__B_op72);
  assign p1_smul_76688_comb = smul32b_32b_x_32b(p0_TestBlock__A_op58, p0_TestBlock__B_op82);
  assign p1_smul_76689_comb = smul32b_32b_x_32b(p0_TestBlock__A_op59, p0_TestBlock__B_op92);
  assign p1_smul_76690_comb = smul32b_32b_x_32b(p0_TestBlock__A_op54, p0_TestBlock__B_op43);
  assign p1_smul_76691_comb = smul32b_32b_x_32b(p0_TestBlock__A_op55, p0_TestBlock__B_op53);
  assign p1_smul_76692_comb = smul32b_32b_x_32b(p0_TestBlock__A_op56, p0_TestBlock__B_op63);
  assign p1_smul_76693_comb = smul32b_32b_x_32b(p0_TestBlock__A_op57, p0_TestBlock__B_op73);
  assign p1_smul_76694_comb = smul32b_32b_x_32b(p0_TestBlock__A_op58, p0_TestBlock__B_op83);
  assign p1_smul_76695_comb = smul32b_32b_x_32b(p0_TestBlock__A_op59, p0_TestBlock__B_op93);
  assign p1_smul_76696_comb = smul32b_32b_x_32b(p0_TestBlock__A_op54, p0_TestBlock__B_op44);
  assign p1_smul_76697_comb = smul32b_32b_x_32b(p0_TestBlock__A_op55, p0_TestBlock__B_op54);
  assign p1_smul_76698_comb = smul32b_32b_x_32b(p0_TestBlock__A_op56, p0_TestBlock__B_op64);
  assign p1_smul_76699_comb = smul32b_32b_x_32b(p0_TestBlock__A_op57, p0_TestBlock__B_op74);
  assign p1_smul_76700_comb = smul32b_32b_x_32b(p0_TestBlock__A_op58, p0_TestBlock__B_op84);
  assign p1_smul_76701_comb = smul32b_32b_x_32b(p0_TestBlock__A_op59, p0_TestBlock__B_op94);
  assign p1_smul_76702_comb = smul32b_32b_x_32b(p0_TestBlock__A_op54, p0_TestBlock__B_op45);
  assign p1_smul_76703_comb = smul32b_32b_x_32b(p0_TestBlock__A_op55, p0_TestBlock__B_op55);
  assign p1_smul_76704_comb = smul32b_32b_x_32b(p0_TestBlock__A_op56, p0_TestBlock__B_op65);
  assign p1_smul_76705_comb = smul32b_32b_x_32b(p0_TestBlock__A_op57, p0_TestBlock__B_op75);
  assign p1_smul_76706_comb = smul32b_32b_x_32b(p0_TestBlock__A_op58, p0_TestBlock__B_op85);
  assign p1_smul_76707_comb = smul32b_32b_x_32b(p0_TestBlock__A_op59, p0_TestBlock__B_op95);
  assign p1_smul_76708_comb = smul32b_32b_x_32b(p0_TestBlock__A_op54, p0_TestBlock__B_op46);
  assign p1_smul_76709_comb = smul32b_32b_x_32b(p0_TestBlock__A_op55, p0_TestBlock__B_op56);
  assign p1_smul_76710_comb = smul32b_32b_x_32b(p0_TestBlock__A_op56, p0_TestBlock__B_op66);
  assign p1_smul_76711_comb = smul32b_32b_x_32b(p0_TestBlock__A_op57, p0_TestBlock__B_op76);
  assign p1_smul_76712_comb = smul32b_32b_x_32b(p0_TestBlock__A_op58, p0_TestBlock__B_op86);
  assign p1_smul_76713_comb = smul32b_32b_x_32b(p0_TestBlock__A_op59, p0_TestBlock__B_op96);
  assign p1_smul_76714_comb = smul32b_32b_x_32b(p0_TestBlock__A_op54, p0_TestBlock__B_op47);
  assign p1_smul_76715_comb = smul32b_32b_x_32b(p0_TestBlock__A_op55, p0_TestBlock__B_op57);
  assign p1_smul_76716_comb = smul32b_32b_x_32b(p0_TestBlock__A_op56, p0_TestBlock__B_op67);
  assign p1_smul_76717_comb = smul32b_32b_x_32b(p0_TestBlock__A_op57, p0_TestBlock__B_op77);
  assign p1_smul_76718_comb = smul32b_32b_x_32b(p0_TestBlock__A_op58, p0_TestBlock__B_op87);
  assign p1_smul_76719_comb = smul32b_32b_x_32b(p0_TestBlock__A_op59, p0_TestBlock__B_op97);
  assign p1_smul_76720_comb = smul32b_32b_x_32b(p0_TestBlock__A_op54, p0_TestBlock__B_op48);
  assign p1_smul_76721_comb = smul32b_32b_x_32b(p0_TestBlock__A_op55, p0_TestBlock__B_op58);
  assign p1_smul_76722_comb = smul32b_32b_x_32b(p0_TestBlock__A_op56, p0_TestBlock__B_op68);
  assign p1_smul_76723_comb = smul32b_32b_x_32b(p0_TestBlock__A_op57, p0_TestBlock__B_op78);
  assign p1_smul_76724_comb = smul32b_32b_x_32b(p0_TestBlock__A_op58, p0_TestBlock__B_op88);
  assign p1_smul_76725_comb = smul32b_32b_x_32b(p0_TestBlock__A_op59, p0_TestBlock__B_op98);
  assign p1_smul_76726_comb = smul32b_32b_x_32b(p0_TestBlock__A_op54, p0_TestBlock__B_op49);
  assign p1_smul_76727_comb = smul32b_32b_x_32b(p0_TestBlock__A_op55, p0_TestBlock__B_op59);
  assign p1_smul_76728_comb = smul32b_32b_x_32b(p0_TestBlock__A_op56, p0_TestBlock__B_op69);
  assign p1_smul_76729_comb = smul32b_32b_x_32b(p0_TestBlock__A_op57, p0_TestBlock__B_op79);
  assign p1_smul_76730_comb = smul32b_32b_x_32b(p0_TestBlock__A_op58, p0_TestBlock__B_op89);
  assign p1_smul_76731_comb = smul32b_32b_x_32b(p0_TestBlock__A_op59, p0_TestBlock__B_op99);
  assign p1_smul_76732_comb = smul32b_32b_x_32b(p0_TestBlock__A_op64, p0_TestBlock__B_op40);
  assign p1_smul_76733_comb = smul32b_32b_x_32b(p0_TestBlock__A_op65, p0_TestBlock__B_op50);
  assign p1_smul_76734_comb = smul32b_32b_x_32b(p0_TestBlock__A_op66, p0_TestBlock__B_op60);
  assign p1_smul_76735_comb = smul32b_32b_x_32b(p0_TestBlock__A_op67, p0_TestBlock__B_op70);
  assign p1_smul_76736_comb = smul32b_32b_x_32b(p0_TestBlock__A_op68, p0_TestBlock__B_op80);
  assign p1_smul_76737_comb = smul32b_32b_x_32b(p0_TestBlock__A_op69, p0_TestBlock__B_op90);
  assign p1_smul_76738_comb = smul32b_32b_x_32b(p0_TestBlock__A_op64, p0_TestBlock__B_op41);
  assign p1_smul_76739_comb = smul32b_32b_x_32b(p0_TestBlock__A_op65, p0_TestBlock__B_op51);
  assign p1_smul_76740_comb = smul32b_32b_x_32b(p0_TestBlock__A_op66, p0_TestBlock__B_op61);
  assign p1_smul_76741_comb = smul32b_32b_x_32b(p0_TestBlock__A_op67, p0_TestBlock__B_op71);
  assign p1_smul_76742_comb = smul32b_32b_x_32b(p0_TestBlock__A_op68, p0_TestBlock__B_op81);
  assign p1_smul_76743_comb = smul32b_32b_x_32b(p0_TestBlock__A_op69, p0_TestBlock__B_op91);
  assign p1_smul_76744_comb = smul32b_32b_x_32b(p0_TestBlock__A_op64, p0_TestBlock__B_op42);
  assign p1_smul_76745_comb = smul32b_32b_x_32b(p0_TestBlock__A_op65, p0_TestBlock__B_op52);
  assign p1_smul_76746_comb = smul32b_32b_x_32b(p0_TestBlock__A_op66, p0_TestBlock__B_op62);
  assign p1_smul_76747_comb = smul32b_32b_x_32b(p0_TestBlock__A_op67, p0_TestBlock__B_op72);
  assign p1_smul_76748_comb = smul32b_32b_x_32b(p0_TestBlock__A_op68, p0_TestBlock__B_op82);
  assign p1_smul_76749_comb = smul32b_32b_x_32b(p0_TestBlock__A_op69, p0_TestBlock__B_op92);
  assign p1_smul_76750_comb = smul32b_32b_x_32b(p0_TestBlock__A_op64, p0_TestBlock__B_op43);
  assign p1_smul_76751_comb = smul32b_32b_x_32b(p0_TestBlock__A_op65, p0_TestBlock__B_op53);
  assign p1_smul_76752_comb = smul32b_32b_x_32b(p0_TestBlock__A_op66, p0_TestBlock__B_op63);
  assign p1_smul_76753_comb = smul32b_32b_x_32b(p0_TestBlock__A_op67, p0_TestBlock__B_op73);
  assign p1_smul_76754_comb = smul32b_32b_x_32b(p0_TestBlock__A_op68, p0_TestBlock__B_op83);
  assign p1_smul_76755_comb = smul32b_32b_x_32b(p0_TestBlock__A_op69, p0_TestBlock__B_op93);
  assign p1_smul_76756_comb = smul32b_32b_x_32b(p0_TestBlock__A_op64, p0_TestBlock__B_op44);
  assign p1_smul_76757_comb = smul32b_32b_x_32b(p0_TestBlock__A_op65, p0_TestBlock__B_op54);
  assign p1_smul_76758_comb = smul32b_32b_x_32b(p0_TestBlock__A_op66, p0_TestBlock__B_op64);
  assign p1_smul_76759_comb = smul32b_32b_x_32b(p0_TestBlock__A_op67, p0_TestBlock__B_op74);
  assign p1_smul_76760_comb = smul32b_32b_x_32b(p0_TestBlock__A_op68, p0_TestBlock__B_op84);
  assign p1_smul_76761_comb = smul32b_32b_x_32b(p0_TestBlock__A_op69, p0_TestBlock__B_op94);
  assign p1_smul_76762_comb = smul32b_32b_x_32b(p0_TestBlock__A_op64, p0_TestBlock__B_op45);
  assign p1_smul_76763_comb = smul32b_32b_x_32b(p0_TestBlock__A_op65, p0_TestBlock__B_op55);
  assign p1_smul_76764_comb = smul32b_32b_x_32b(p0_TestBlock__A_op66, p0_TestBlock__B_op65);
  assign p1_smul_76765_comb = smul32b_32b_x_32b(p0_TestBlock__A_op67, p0_TestBlock__B_op75);
  assign p1_smul_76766_comb = smul32b_32b_x_32b(p0_TestBlock__A_op68, p0_TestBlock__B_op85);
  assign p1_smul_76767_comb = smul32b_32b_x_32b(p0_TestBlock__A_op69, p0_TestBlock__B_op95);
  assign p1_smul_76768_comb = smul32b_32b_x_32b(p0_TestBlock__A_op64, p0_TestBlock__B_op46);
  assign p1_smul_76769_comb = smul32b_32b_x_32b(p0_TestBlock__A_op65, p0_TestBlock__B_op56);
  assign p1_smul_76770_comb = smul32b_32b_x_32b(p0_TestBlock__A_op66, p0_TestBlock__B_op66);
  assign p1_smul_76771_comb = smul32b_32b_x_32b(p0_TestBlock__A_op67, p0_TestBlock__B_op76);
  assign p1_smul_76772_comb = smul32b_32b_x_32b(p0_TestBlock__A_op68, p0_TestBlock__B_op86);
  assign p1_smul_76773_comb = smul32b_32b_x_32b(p0_TestBlock__A_op69, p0_TestBlock__B_op96);
  assign p1_smul_76774_comb = smul32b_32b_x_32b(p0_TestBlock__A_op64, p0_TestBlock__B_op47);
  assign p1_smul_76775_comb = smul32b_32b_x_32b(p0_TestBlock__A_op65, p0_TestBlock__B_op57);
  assign p1_smul_76776_comb = smul32b_32b_x_32b(p0_TestBlock__A_op66, p0_TestBlock__B_op67);
  assign p1_smul_76777_comb = smul32b_32b_x_32b(p0_TestBlock__A_op67, p0_TestBlock__B_op77);
  assign p1_smul_76778_comb = smul32b_32b_x_32b(p0_TestBlock__A_op68, p0_TestBlock__B_op87);
  assign p1_smul_76779_comb = smul32b_32b_x_32b(p0_TestBlock__A_op69, p0_TestBlock__B_op97);
  assign p1_smul_76780_comb = smul32b_32b_x_32b(p0_TestBlock__A_op64, p0_TestBlock__B_op48);
  assign p1_smul_76781_comb = smul32b_32b_x_32b(p0_TestBlock__A_op65, p0_TestBlock__B_op58);
  assign p1_smul_76782_comb = smul32b_32b_x_32b(p0_TestBlock__A_op66, p0_TestBlock__B_op68);
  assign p1_smul_76783_comb = smul32b_32b_x_32b(p0_TestBlock__A_op67, p0_TestBlock__B_op78);
  assign p1_smul_76784_comb = smul32b_32b_x_32b(p0_TestBlock__A_op68, p0_TestBlock__B_op88);
  assign p1_smul_76785_comb = smul32b_32b_x_32b(p0_TestBlock__A_op69, p0_TestBlock__B_op98);
  assign p1_smul_76786_comb = smul32b_32b_x_32b(p0_TestBlock__A_op64, p0_TestBlock__B_op49);
  assign p1_smul_76787_comb = smul32b_32b_x_32b(p0_TestBlock__A_op65, p0_TestBlock__B_op59);
  assign p1_smul_76788_comb = smul32b_32b_x_32b(p0_TestBlock__A_op66, p0_TestBlock__B_op69);
  assign p1_smul_76789_comb = smul32b_32b_x_32b(p0_TestBlock__A_op67, p0_TestBlock__B_op79);
  assign p1_smul_76790_comb = smul32b_32b_x_32b(p0_TestBlock__A_op68, p0_TestBlock__B_op89);
  assign p1_smul_76791_comb = smul32b_32b_x_32b(p0_TestBlock__A_op69, p0_TestBlock__B_op99);
  assign p1_smul_76792_comb = smul32b_32b_x_32b(p0_TestBlock__A_op74, p0_TestBlock__B_op40);
  assign p1_smul_76793_comb = smul32b_32b_x_32b(p0_TestBlock__A_op75, p0_TestBlock__B_op50);
  assign p1_smul_76794_comb = smul32b_32b_x_32b(p0_TestBlock__A_op76, p0_TestBlock__B_op60);
  assign p1_smul_76795_comb = smul32b_32b_x_32b(p0_TestBlock__A_op77, p0_TestBlock__B_op70);
  assign p1_smul_76796_comb = smul32b_32b_x_32b(p0_TestBlock__A_op78, p0_TestBlock__B_op80);
  assign p1_smul_76797_comb = smul32b_32b_x_32b(p0_TestBlock__A_op79, p0_TestBlock__B_op90);
  assign p1_smul_76798_comb = smul32b_32b_x_32b(p0_TestBlock__A_op74, p0_TestBlock__B_op41);
  assign p1_smul_76799_comb = smul32b_32b_x_32b(p0_TestBlock__A_op75, p0_TestBlock__B_op51);
  assign p1_smul_76800_comb = smul32b_32b_x_32b(p0_TestBlock__A_op76, p0_TestBlock__B_op61);
  assign p1_smul_76801_comb = smul32b_32b_x_32b(p0_TestBlock__A_op77, p0_TestBlock__B_op71);
  assign p1_smul_76802_comb = smul32b_32b_x_32b(p0_TestBlock__A_op78, p0_TestBlock__B_op81);
  assign p1_smul_76803_comb = smul32b_32b_x_32b(p0_TestBlock__A_op79, p0_TestBlock__B_op91);
  assign p1_smul_76804_comb = smul32b_32b_x_32b(p0_TestBlock__A_op74, p0_TestBlock__B_op42);
  assign p1_smul_76805_comb = smul32b_32b_x_32b(p0_TestBlock__A_op75, p0_TestBlock__B_op52);
  assign p1_smul_76806_comb = smul32b_32b_x_32b(p0_TestBlock__A_op76, p0_TestBlock__B_op62);
  assign p1_smul_76807_comb = smul32b_32b_x_32b(p0_TestBlock__A_op77, p0_TestBlock__B_op72);
  assign p1_smul_76808_comb = smul32b_32b_x_32b(p0_TestBlock__A_op78, p0_TestBlock__B_op82);
  assign p1_smul_76809_comb = smul32b_32b_x_32b(p0_TestBlock__A_op79, p0_TestBlock__B_op92);
  assign p1_smul_76810_comb = smul32b_32b_x_32b(p0_TestBlock__A_op74, p0_TestBlock__B_op43);
  assign p1_smul_76811_comb = smul32b_32b_x_32b(p0_TestBlock__A_op75, p0_TestBlock__B_op53);
  assign p1_smul_76812_comb = smul32b_32b_x_32b(p0_TestBlock__A_op76, p0_TestBlock__B_op63);
  assign p1_smul_76813_comb = smul32b_32b_x_32b(p0_TestBlock__A_op77, p0_TestBlock__B_op73);
  assign p1_smul_76814_comb = smul32b_32b_x_32b(p0_TestBlock__A_op78, p0_TestBlock__B_op83);
  assign p1_smul_76815_comb = smul32b_32b_x_32b(p0_TestBlock__A_op79, p0_TestBlock__B_op93);
  assign p1_smul_76816_comb = smul32b_32b_x_32b(p0_TestBlock__A_op74, p0_TestBlock__B_op44);
  assign p1_smul_76817_comb = smul32b_32b_x_32b(p0_TestBlock__A_op75, p0_TestBlock__B_op54);
  assign p1_smul_76818_comb = smul32b_32b_x_32b(p0_TestBlock__A_op76, p0_TestBlock__B_op64);
  assign p1_smul_76819_comb = smul32b_32b_x_32b(p0_TestBlock__A_op77, p0_TestBlock__B_op74);
  assign p1_smul_76820_comb = smul32b_32b_x_32b(p0_TestBlock__A_op78, p0_TestBlock__B_op84);
  assign p1_smul_76821_comb = smul32b_32b_x_32b(p0_TestBlock__A_op79, p0_TestBlock__B_op94);
  assign p1_smul_76822_comb = smul32b_32b_x_32b(p0_TestBlock__A_op74, p0_TestBlock__B_op45);
  assign p1_smul_76823_comb = smul32b_32b_x_32b(p0_TestBlock__A_op75, p0_TestBlock__B_op55);
  assign p1_smul_76824_comb = smul32b_32b_x_32b(p0_TestBlock__A_op76, p0_TestBlock__B_op65);
  assign p1_smul_76825_comb = smul32b_32b_x_32b(p0_TestBlock__A_op77, p0_TestBlock__B_op75);
  assign p1_smul_76826_comb = smul32b_32b_x_32b(p0_TestBlock__A_op78, p0_TestBlock__B_op85);
  assign p1_smul_76827_comb = smul32b_32b_x_32b(p0_TestBlock__A_op79, p0_TestBlock__B_op95);
  assign p1_smul_76828_comb = smul32b_32b_x_32b(p0_TestBlock__A_op74, p0_TestBlock__B_op46);
  assign p1_smul_76829_comb = smul32b_32b_x_32b(p0_TestBlock__A_op75, p0_TestBlock__B_op56);
  assign p1_smul_76830_comb = smul32b_32b_x_32b(p0_TestBlock__A_op76, p0_TestBlock__B_op66);
  assign p1_smul_76831_comb = smul32b_32b_x_32b(p0_TestBlock__A_op77, p0_TestBlock__B_op76);
  assign p1_smul_76832_comb = smul32b_32b_x_32b(p0_TestBlock__A_op78, p0_TestBlock__B_op86);
  assign p1_smul_76833_comb = smul32b_32b_x_32b(p0_TestBlock__A_op79, p0_TestBlock__B_op96);
  assign p1_smul_76834_comb = smul32b_32b_x_32b(p0_TestBlock__A_op74, p0_TestBlock__B_op47);
  assign p1_smul_76835_comb = smul32b_32b_x_32b(p0_TestBlock__A_op75, p0_TestBlock__B_op57);
  assign p1_smul_76836_comb = smul32b_32b_x_32b(p0_TestBlock__A_op76, p0_TestBlock__B_op67);
  assign p1_smul_76837_comb = smul32b_32b_x_32b(p0_TestBlock__A_op77, p0_TestBlock__B_op77);
  assign p1_smul_76838_comb = smul32b_32b_x_32b(p0_TestBlock__A_op78, p0_TestBlock__B_op87);
  assign p1_smul_76839_comb = smul32b_32b_x_32b(p0_TestBlock__A_op79, p0_TestBlock__B_op97);
  assign p1_smul_76840_comb = smul32b_32b_x_32b(p0_TestBlock__A_op74, p0_TestBlock__B_op48);
  assign p1_smul_76841_comb = smul32b_32b_x_32b(p0_TestBlock__A_op75, p0_TestBlock__B_op58);
  assign p1_smul_76842_comb = smul32b_32b_x_32b(p0_TestBlock__A_op76, p0_TestBlock__B_op68);
  assign p1_smul_76843_comb = smul32b_32b_x_32b(p0_TestBlock__A_op77, p0_TestBlock__B_op78);
  assign p1_smul_76844_comb = smul32b_32b_x_32b(p0_TestBlock__A_op78, p0_TestBlock__B_op88);
  assign p1_smul_76845_comb = smul32b_32b_x_32b(p0_TestBlock__A_op79, p0_TestBlock__B_op98);
  assign p1_smul_76846_comb = smul32b_32b_x_32b(p0_TestBlock__A_op74, p0_TestBlock__B_op49);
  assign p1_smul_76847_comb = smul32b_32b_x_32b(p0_TestBlock__A_op75, p0_TestBlock__B_op59);
  assign p1_smul_76848_comb = smul32b_32b_x_32b(p0_TestBlock__A_op76, p0_TestBlock__B_op69);
  assign p1_smul_76849_comb = smul32b_32b_x_32b(p0_TestBlock__A_op77, p0_TestBlock__B_op79);
  assign p1_smul_76850_comb = smul32b_32b_x_32b(p0_TestBlock__A_op78, p0_TestBlock__B_op89);
  assign p1_smul_76851_comb = smul32b_32b_x_32b(p0_TestBlock__A_op79, p0_TestBlock__B_op99);
  assign p1_smul_76852_comb = smul32b_32b_x_32b(p0_TestBlock__A_op84, p0_TestBlock__B_op40);
  assign p1_smul_76853_comb = smul32b_32b_x_32b(p0_TestBlock__A_op85, p0_TestBlock__B_op50);
  assign p1_smul_76854_comb = smul32b_32b_x_32b(p0_TestBlock__A_op86, p0_TestBlock__B_op60);
  assign p1_smul_76855_comb = smul32b_32b_x_32b(p0_TestBlock__A_op87, p0_TestBlock__B_op70);
  assign p1_smul_76856_comb = smul32b_32b_x_32b(p0_TestBlock__A_op88, p0_TestBlock__B_op80);
  assign p1_smul_76857_comb = smul32b_32b_x_32b(p0_TestBlock__A_op89, p0_TestBlock__B_op90);
  assign p1_smul_76858_comb = smul32b_32b_x_32b(p0_TestBlock__A_op84, p0_TestBlock__B_op41);
  assign p1_smul_76859_comb = smul32b_32b_x_32b(p0_TestBlock__A_op85, p0_TestBlock__B_op51);
  assign p1_smul_76860_comb = smul32b_32b_x_32b(p0_TestBlock__A_op86, p0_TestBlock__B_op61);
  assign p1_smul_76861_comb = smul32b_32b_x_32b(p0_TestBlock__A_op87, p0_TestBlock__B_op71);
  assign p1_smul_76862_comb = smul32b_32b_x_32b(p0_TestBlock__A_op88, p0_TestBlock__B_op81);
  assign p1_smul_76863_comb = smul32b_32b_x_32b(p0_TestBlock__A_op89, p0_TestBlock__B_op91);
  assign p1_smul_76864_comb = smul32b_32b_x_32b(p0_TestBlock__A_op84, p0_TestBlock__B_op42);
  assign p1_smul_76865_comb = smul32b_32b_x_32b(p0_TestBlock__A_op85, p0_TestBlock__B_op52);
  assign p1_smul_76866_comb = smul32b_32b_x_32b(p0_TestBlock__A_op86, p0_TestBlock__B_op62);
  assign p1_smul_76867_comb = smul32b_32b_x_32b(p0_TestBlock__A_op87, p0_TestBlock__B_op72);
  assign p1_smul_76868_comb = smul32b_32b_x_32b(p0_TestBlock__A_op88, p0_TestBlock__B_op82);
  assign p1_smul_76869_comb = smul32b_32b_x_32b(p0_TestBlock__A_op89, p0_TestBlock__B_op92);
  assign p1_smul_76870_comb = smul32b_32b_x_32b(p0_TestBlock__A_op84, p0_TestBlock__B_op43);
  assign p1_smul_76871_comb = smul32b_32b_x_32b(p0_TestBlock__A_op85, p0_TestBlock__B_op53);
  assign p1_smul_76872_comb = smul32b_32b_x_32b(p0_TestBlock__A_op86, p0_TestBlock__B_op63);
  assign p1_smul_76873_comb = smul32b_32b_x_32b(p0_TestBlock__A_op87, p0_TestBlock__B_op73);
  assign p1_smul_76874_comb = smul32b_32b_x_32b(p0_TestBlock__A_op88, p0_TestBlock__B_op83);
  assign p1_smul_76875_comb = smul32b_32b_x_32b(p0_TestBlock__A_op89, p0_TestBlock__B_op93);
  assign p1_smul_76876_comb = smul32b_32b_x_32b(p0_TestBlock__A_op84, p0_TestBlock__B_op44);
  assign p1_smul_76877_comb = smul32b_32b_x_32b(p0_TestBlock__A_op85, p0_TestBlock__B_op54);
  assign p1_smul_76878_comb = smul32b_32b_x_32b(p0_TestBlock__A_op86, p0_TestBlock__B_op64);
  assign p1_smul_76879_comb = smul32b_32b_x_32b(p0_TestBlock__A_op87, p0_TestBlock__B_op74);
  assign p1_smul_76880_comb = smul32b_32b_x_32b(p0_TestBlock__A_op88, p0_TestBlock__B_op84);
  assign p1_smul_76881_comb = smul32b_32b_x_32b(p0_TestBlock__A_op89, p0_TestBlock__B_op94);
  assign p1_smul_76882_comb = smul32b_32b_x_32b(p0_TestBlock__A_op84, p0_TestBlock__B_op45);
  assign p1_smul_76883_comb = smul32b_32b_x_32b(p0_TestBlock__A_op85, p0_TestBlock__B_op55);
  assign p1_smul_76884_comb = smul32b_32b_x_32b(p0_TestBlock__A_op86, p0_TestBlock__B_op65);
  assign p1_smul_76885_comb = smul32b_32b_x_32b(p0_TestBlock__A_op87, p0_TestBlock__B_op75);
  assign p1_smul_76886_comb = smul32b_32b_x_32b(p0_TestBlock__A_op88, p0_TestBlock__B_op85);
  assign p1_smul_76887_comb = smul32b_32b_x_32b(p0_TestBlock__A_op89, p0_TestBlock__B_op95);
  assign p1_smul_76888_comb = smul32b_32b_x_32b(p0_TestBlock__A_op84, p0_TestBlock__B_op46);
  assign p1_smul_76889_comb = smul32b_32b_x_32b(p0_TestBlock__A_op85, p0_TestBlock__B_op56);
  assign p1_smul_76890_comb = smul32b_32b_x_32b(p0_TestBlock__A_op86, p0_TestBlock__B_op66);
  assign p1_smul_76891_comb = smul32b_32b_x_32b(p0_TestBlock__A_op87, p0_TestBlock__B_op76);
  assign p1_smul_76892_comb = smul32b_32b_x_32b(p0_TestBlock__A_op88, p0_TestBlock__B_op86);
  assign p1_smul_76893_comb = smul32b_32b_x_32b(p0_TestBlock__A_op89, p0_TestBlock__B_op96);
  assign p1_smul_76894_comb = smul32b_32b_x_32b(p0_TestBlock__A_op84, p0_TestBlock__B_op47);
  assign p1_smul_76895_comb = smul32b_32b_x_32b(p0_TestBlock__A_op85, p0_TestBlock__B_op57);
  assign p1_smul_76896_comb = smul32b_32b_x_32b(p0_TestBlock__A_op86, p0_TestBlock__B_op67);
  assign p1_smul_76897_comb = smul32b_32b_x_32b(p0_TestBlock__A_op87, p0_TestBlock__B_op77);
  assign p1_smul_76898_comb = smul32b_32b_x_32b(p0_TestBlock__A_op88, p0_TestBlock__B_op87);
  assign p1_smul_76899_comb = smul32b_32b_x_32b(p0_TestBlock__A_op89, p0_TestBlock__B_op97);
  assign p1_smul_76900_comb = smul32b_32b_x_32b(p0_TestBlock__A_op84, p0_TestBlock__B_op48);
  assign p1_smul_76901_comb = smul32b_32b_x_32b(p0_TestBlock__A_op85, p0_TestBlock__B_op58);
  assign p1_smul_76902_comb = smul32b_32b_x_32b(p0_TestBlock__A_op86, p0_TestBlock__B_op68);
  assign p1_smul_76903_comb = smul32b_32b_x_32b(p0_TestBlock__A_op87, p0_TestBlock__B_op78);
  assign p1_smul_76904_comb = smul32b_32b_x_32b(p0_TestBlock__A_op88, p0_TestBlock__B_op88);
  assign p1_smul_76905_comb = smul32b_32b_x_32b(p0_TestBlock__A_op89, p0_TestBlock__B_op98);
  assign p1_smul_76906_comb = smul32b_32b_x_32b(p0_TestBlock__A_op84, p0_TestBlock__B_op49);
  assign p1_smul_76907_comb = smul32b_32b_x_32b(p0_TestBlock__A_op85, p0_TestBlock__B_op59);
  assign p1_smul_76908_comb = smul32b_32b_x_32b(p0_TestBlock__A_op86, p0_TestBlock__B_op69);
  assign p1_smul_76909_comb = smul32b_32b_x_32b(p0_TestBlock__A_op87, p0_TestBlock__B_op79);
  assign p1_smul_76910_comb = smul32b_32b_x_32b(p0_TestBlock__A_op88, p0_TestBlock__B_op89);
  assign p1_smul_76911_comb = smul32b_32b_x_32b(p0_TestBlock__A_op89, p0_TestBlock__B_op99);
  assign p1_smul_76912_comb = smul32b_32b_x_32b(p0_TestBlock__A_op94, p0_TestBlock__B_op40);
  assign p1_smul_76913_comb = smul32b_32b_x_32b(p0_TestBlock__A_op95, p0_TestBlock__B_op50);
  assign p1_smul_76914_comb = smul32b_32b_x_32b(p0_TestBlock__A_op96, p0_TestBlock__B_op60);
  assign p1_smul_76915_comb = smul32b_32b_x_32b(p0_TestBlock__A_op97, p0_TestBlock__B_op70);
  assign p1_smul_76916_comb = smul32b_32b_x_32b(p0_TestBlock__A_op98, p0_TestBlock__B_op80);
  assign p1_smul_76917_comb = smul32b_32b_x_32b(p0_TestBlock__A_op99, p0_TestBlock__B_op90);
  assign p1_smul_76918_comb = smul32b_32b_x_32b(p0_TestBlock__A_op94, p0_TestBlock__B_op41);
  assign p1_smul_76919_comb = smul32b_32b_x_32b(p0_TestBlock__A_op95, p0_TestBlock__B_op51);
  assign p1_smul_76920_comb = smul32b_32b_x_32b(p0_TestBlock__A_op96, p0_TestBlock__B_op61);
  assign p1_smul_76921_comb = smul32b_32b_x_32b(p0_TestBlock__A_op97, p0_TestBlock__B_op71);
  assign p1_smul_76922_comb = smul32b_32b_x_32b(p0_TestBlock__A_op98, p0_TestBlock__B_op81);
  assign p1_smul_76923_comb = smul32b_32b_x_32b(p0_TestBlock__A_op99, p0_TestBlock__B_op91);
  assign p1_smul_76924_comb = smul32b_32b_x_32b(p0_TestBlock__A_op94, p0_TestBlock__B_op42);
  assign p1_smul_76925_comb = smul32b_32b_x_32b(p0_TestBlock__A_op95, p0_TestBlock__B_op52);
  assign p1_smul_76926_comb = smul32b_32b_x_32b(p0_TestBlock__A_op96, p0_TestBlock__B_op62);
  assign p1_smul_76927_comb = smul32b_32b_x_32b(p0_TestBlock__A_op97, p0_TestBlock__B_op72);
  assign p1_smul_76928_comb = smul32b_32b_x_32b(p0_TestBlock__A_op98, p0_TestBlock__B_op82);
  assign p1_smul_76929_comb = smul32b_32b_x_32b(p0_TestBlock__A_op99, p0_TestBlock__B_op92);
  assign p1_smul_76930_comb = smul32b_32b_x_32b(p0_TestBlock__A_op94, p0_TestBlock__B_op43);
  assign p1_smul_76931_comb = smul32b_32b_x_32b(p0_TestBlock__A_op95, p0_TestBlock__B_op53);
  assign p1_smul_76932_comb = smul32b_32b_x_32b(p0_TestBlock__A_op96, p0_TestBlock__B_op63);
  assign p1_smul_76933_comb = smul32b_32b_x_32b(p0_TestBlock__A_op97, p0_TestBlock__B_op73);
  assign p1_smul_76934_comb = smul32b_32b_x_32b(p0_TestBlock__A_op98, p0_TestBlock__B_op83);
  assign p1_smul_76935_comb = smul32b_32b_x_32b(p0_TestBlock__A_op99, p0_TestBlock__B_op93);
  assign p1_smul_76936_comb = smul32b_32b_x_32b(p0_TestBlock__A_op94, p0_TestBlock__B_op44);
  assign p1_smul_76937_comb = smul32b_32b_x_32b(p0_TestBlock__A_op95, p0_TestBlock__B_op54);
  assign p1_smul_76938_comb = smul32b_32b_x_32b(p0_TestBlock__A_op96, p0_TestBlock__B_op64);
  assign p1_smul_76939_comb = smul32b_32b_x_32b(p0_TestBlock__A_op97, p0_TestBlock__B_op74);
  assign p1_smul_76940_comb = smul32b_32b_x_32b(p0_TestBlock__A_op98, p0_TestBlock__B_op84);
  assign p1_smul_76941_comb = smul32b_32b_x_32b(p0_TestBlock__A_op99, p0_TestBlock__B_op94);
  assign p1_smul_76942_comb = smul32b_32b_x_32b(p0_TestBlock__A_op94, p0_TestBlock__B_op45);
  assign p1_smul_76943_comb = smul32b_32b_x_32b(p0_TestBlock__A_op95, p0_TestBlock__B_op55);
  assign p1_smul_76944_comb = smul32b_32b_x_32b(p0_TestBlock__A_op96, p0_TestBlock__B_op65);
  assign p1_smul_76945_comb = smul32b_32b_x_32b(p0_TestBlock__A_op97, p0_TestBlock__B_op75);
  assign p1_smul_76946_comb = smul32b_32b_x_32b(p0_TestBlock__A_op98, p0_TestBlock__B_op85);
  assign p1_smul_76947_comb = smul32b_32b_x_32b(p0_TestBlock__A_op99, p0_TestBlock__B_op95);
  assign p1_smul_76948_comb = smul32b_32b_x_32b(p0_TestBlock__A_op94, p0_TestBlock__B_op46);
  assign p1_smul_76949_comb = smul32b_32b_x_32b(p0_TestBlock__A_op95, p0_TestBlock__B_op56);
  assign p1_smul_76950_comb = smul32b_32b_x_32b(p0_TestBlock__A_op96, p0_TestBlock__B_op66);
  assign p1_smul_76951_comb = smul32b_32b_x_32b(p0_TestBlock__A_op97, p0_TestBlock__B_op76);
  assign p1_smul_76952_comb = smul32b_32b_x_32b(p0_TestBlock__A_op98, p0_TestBlock__B_op86);
  assign p1_smul_76953_comb = smul32b_32b_x_32b(p0_TestBlock__A_op99, p0_TestBlock__B_op96);
  assign p1_smul_76954_comb = smul32b_32b_x_32b(p0_TestBlock__A_op94, p0_TestBlock__B_op47);
  assign p1_smul_76955_comb = smul32b_32b_x_32b(p0_TestBlock__A_op95, p0_TestBlock__B_op57);
  assign p1_smul_76956_comb = smul32b_32b_x_32b(p0_TestBlock__A_op96, p0_TestBlock__B_op67);
  assign p1_smul_76957_comb = smul32b_32b_x_32b(p0_TestBlock__A_op97, p0_TestBlock__B_op77);
  assign p1_smul_76958_comb = smul32b_32b_x_32b(p0_TestBlock__A_op98, p0_TestBlock__B_op87);
  assign p1_smul_76959_comb = smul32b_32b_x_32b(p0_TestBlock__A_op99, p0_TestBlock__B_op97);
  assign p1_smul_76960_comb = smul32b_32b_x_32b(p0_TestBlock__A_op94, p0_TestBlock__B_op48);
  assign p1_smul_76961_comb = smul32b_32b_x_32b(p0_TestBlock__A_op95, p0_TestBlock__B_op58);
  assign p1_smul_76962_comb = smul32b_32b_x_32b(p0_TestBlock__A_op96, p0_TestBlock__B_op68);
  assign p1_smul_76963_comb = smul32b_32b_x_32b(p0_TestBlock__A_op97, p0_TestBlock__B_op78);
  assign p1_smul_76964_comb = smul32b_32b_x_32b(p0_TestBlock__A_op98, p0_TestBlock__B_op88);
  assign p1_smul_76965_comb = smul32b_32b_x_32b(p0_TestBlock__A_op99, p0_TestBlock__B_op98);
  assign p1_smul_76966_comb = smul32b_32b_x_32b(p0_TestBlock__A_op94, p0_TestBlock__B_op49);
  assign p1_smul_76967_comb = smul32b_32b_x_32b(p0_TestBlock__A_op95, p0_TestBlock__B_op59);
  assign p1_smul_76968_comb = smul32b_32b_x_32b(p0_TestBlock__A_op96, p0_TestBlock__B_op69);
  assign p1_smul_76969_comb = smul32b_32b_x_32b(p0_TestBlock__A_op97, p0_TestBlock__B_op79);
  assign p1_smul_76970_comb = smul32b_32b_x_32b(p0_TestBlock__A_op98, p0_TestBlock__B_op89);
  assign p1_smul_76971_comb = smul32b_32b_x_32b(p0_TestBlock__A_op99, p0_TestBlock__B_op99);

  // Registers for pipe stage 1:
  reg [31:0] p1_smul_75972;
  reg [31:0] p1_smul_75973;
  reg [31:0] p1_smul_75974;
  reg [31:0] p1_smul_75975;
  reg [31:0] p1_smul_75976;
  reg [31:0] p1_smul_75977;
  reg [31:0] p1_smul_75978;
  reg [31:0] p1_smul_75979;
  reg [31:0] p1_smul_75980;
  reg [31:0] p1_smul_75981;
  reg [31:0] p1_smul_75982;
  reg [31:0] p1_smul_75983;
  reg [31:0] p1_smul_75984;
  reg [31:0] p1_smul_75985;
  reg [31:0] p1_smul_75986;
  reg [31:0] p1_smul_75987;
  reg [31:0] p1_smul_75988;
  reg [31:0] p1_smul_75989;
  reg [31:0] p1_smul_75990;
  reg [31:0] p1_smul_75991;
  reg [31:0] p1_smul_75992;
  reg [31:0] p1_smul_75993;
  reg [31:0] p1_smul_75994;
  reg [31:0] p1_smul_75995;
  reg [31:0] p1_smul_75996;
  reg [31:0] p1_smul_75997;
  reg [31:0] p1_smul_75998;
  reg [31:0] p1_smul_75999;
  reg [31:0] p1_smul_76000;
  reg [31:0] p1_smul_76001;
  reg [31:0] p1_smul_76002;
  reg [31:0] p1_smul_76003;
  reg [31:0] p1_smul_76004;
  reg [31:0] p1_smul_76005;
  reg [31:0] p1_smul_76006;
  reg [31:0] p1_smul_76007;
  reg [31:0] p1_smul_76008;
  reg [31:0] p1_smul_76009;
  reg [31:0] p1_smul_76010;
  reg [31:0] p1_smul_76011;
  reg [31:0] p1_smul_76012;
  reg [31:0] p1_smul_76013;
  reg [31:0] p1_smul_76014;
  reg [31:0] p1_smul_76015;
  reg [31:0] p1_smul_76016;
  reg [31:0] p1_smul_76017;
  reg [31:0] p1_smul_76018;
  reg [31:0] p1_smul_76019;
  reg [31:0] p1_smul_76020;
  reg [31:0] p1_smul_76021;
  reg [31:0] p1_smul_76022;
  reg [31:0] p1_smul_76023;
  reg [31:0] p1_smul_76024;
  reg [31:0] p1_smul_76025;
  reg [31:0] p1_smul_76026;
  reg [31:0] p1_smul_76027;
  reg [31:0] p1_smul_76028;
  reg [31:0] p1_smul_76029;
  reg [31:0] p1_smul_76030;
  reg [31:0] p1_smul_76031;
  reg [31:0] p1_smul_76032;
  reg [31:0] p1_smul_76033;
  reg [31:0] p1_smul_76034;
  reg [31:0] p1_smul_76035;
  reg [31:0] p1_smul_76036;
  reg [31:0] p1_smul_76037;
  reg [31:0] p1_smul_76038;
  reg [31:0] p1_smul_76039;
  reg [31:0] p1_smul_76040;
  reg [31:0] p1_smul_76041;
  reg [31:0] p1_smul_76042;
  reg [31:0] p1_smul_76043;
  reg [31:0] p1_smul_76044;
  reg [31:0] p1_smul_76045;
  reg [31:0] p1_smul_76046;
  reg [31:0] p1_smul_76047;
  reg [31:0] p1_smul_76048;
  reg [31:0] p1_smul_76049;
  reg [31:0] p1_smul_76050;
  reg [31:0] p1_smul_76051;
  reg [31:0] p1_smul_76052;
  reg [31:0] p1_smul_76053;
  reg [31:0] p1_smul_76054;
  reg [31:0] p1_smul_76055;
  reg [31:0] p1_smul_76056;
  reg [31:0] p1_smul_76057;
  reg [31:0] p1_smul_76058;
  reg [31:0] p1_smul_76059;
  reg [31:0] p1_smul_76060;
  reg [31:0] p1_smul_76061;
  reg [31:0] p1_smul_76062;
  reg [31:0] p1_smul_76063;
  reg [31:0] p1_smul_76064;
  reg [31:0] p1_smul_76065;
  reg [31:0] p1_smul_76066;
  reg [31:0] p1_smul_76067;
  reg [31:0] p1_smul_76068;
  reg [31:0] p1_smul_76069;
  reg [31:0] p1_smul_76070;
  reg [31:0] p1_smul_76071;
  reg [31:0] p1_smul_76072;
  reg [31:0] p1_smul_76073;
  reg [31:0] p1_smul_76074;
  reg [31:0] p1_smul_76075;
  reg [31:0] p1_smul_76076;
  reg [31:0] p1_smul_76077;
  reg [31:0] p1_smul_76078;
  reg [31:0] p1_smul_76079;
  reg [31:0] p1_smul_76080;
  reg [31:0] p1_smul_76081;
  reg [31:0] p1_smul_76082;
  reg [31:0] p1_smul_76083;
  reg [31:0] p1_smul_76084;
  reg [31:0] p1_smul_76085;
  reg [31:0] p1_smul_76086;
  reg [31:0] p1_smul_76087;
  reg [31:0] p1_smul_76088;
  reg [31:0] p1_smul_76089;
  reg [31:0] p1_smul_76090;
  reg [31:0] p1_smul_76091;
  reg [31:0] p1_smul_76092;
  reg [31:0] p1_smul_76093;
  reg [31:0] p1_smul_76094;
  reg [31:0] p1_smul_76095;
  reg [31:0] p1_smul_76096;
  reg [31:0] p1_smul_76097;
  reg [31:0] p1_smul_76098;
  reg [31:0] p1_smul_76099;
  reg [31:0] p1_smul_76100;
  reg [31:0] p1_smul_76101;
  reg [31:0] p1_smul_76102;
  reg [31:0] p1_smul_76103;
  reg [31:0] p1_smul_76104;
  reg [31:0] p1_smul_76105;
  reg [31:0] p1_smul_76106;
  reg [31:0] p1_smul_76107;
  reg [31:0] p1_smul_76108;
  reg [31:0] p1_smul_76109;
  reg [31:0] p1_smul_76110;
  reg [31:0] p1_smul_76111;
  reg [31:0] p1_smul_76112;
  reg [31:0] p1_smul_76113;
  reg [31:0] p1_smul_76114;
  reg [31:0] p1_smul_76115;
  reg [31:0] p1_smul_76116;
  reg [31:0] p1_smul_76117;
  reg [31:0] p1_smul_76118;
  reg [31:0] p1_smul_76119;
  reg [31:0] p1_smul_76120;
  reg [31:0] p1_smul_76121;
  reg [31:0] p1_smul_76122;
  reg [31:0] p1_smul_76123;
  reg [31:0] p1_smul_76124;
  reg [31:0] p1_smul_76125;
  reg [31:0] p1_smul_76126;
  reg [31:0] p1_smul_76127;
  reg [31:0] p1_smul_76128;
  reg [31:0] p1_smul_76129;
  reg [31:0] p1_smul_76130;
  reg [31:0] p1_smul_76131;
  reg [31:0] p1_smul_76132;
  reg [31:0] p1_smul_76133;
  reg [31:0] p1_smul_76134;
  reg [31:0] p1_smul_76135;
  reg [31:0] p1_smul_76136;
  reg [31:0] p1_smul_76137;
  reg [31:0] p1_smul_76138;
  reg [31:0] p1_smul_76139;
  reg [31:0] p1_smul_76140;
  reg [31:0] p1_smul_76141;
  reg [31:0] p1_smul_76142;
  reg [31:0] p1_smul_76143;
  reg [31:0] p1_smul_76144;
  reg [31:0] p1_smul_76145;
  reg [31:0] p1_smul_76146;
  reg [31:0] p1_smul_76147;
  reg [31:0] p1_smul_76148;
  reg [31:0] p1_smul_76149;
  reg [31:0] p1_smul_76150;
  reg [31:0] p1_smul_76151;
  reg [31:0] p1_smul_76152;
  reg [31:0] p1_smul_76153;
  reg [31:0] p1_smul_76154;
  reg [31:0] p1_smul_76155;
  reg [31:0] p1_smul_76156;
  reg [31:0] p1_smul_76157;
  reg [31:0] p1_smul_76158;
  reg [31:0] p1_smul_76159;
  reg [31:0] p1_smul_76160;
  reg [31:0] p1_smul_76161;
  reg [31:0] p1_smul_76162;
  reg [31:0] p1_smul_76163;
  reg [31:0] p1_smul_76164;
  reg [31:0] p1_smul_76165;
  reg [31:0] p1_smul_76166;
  reg [31:0] p1_smul_76167;
  reg [31:0] p1_smul_76168;
  reg [31:0] p1_smul_76169;
  reg [31:0] p1_smul_76170;
  reg [31:0] p1_smul_76171;
  reg [31:0] p1_smul_76172;
  reg [31:0] p1_smul_76173;
  reg [31:0] p1_smul_76174;
  reg [31:0] p1_smul_76175;
  reg [31:0] p1_smul_76176;
  reg [31:0] p1_smul_76177;
  reg [31:0] p1_smul_76178;
  reg [31:0] p1_smul_76179;
  reg [31:0] p1_smul_76180;
  reg [31:0] p1_smul_76181;
  reg [31:0] p1_smul_76182;
  reg [31:0] p1_smul_76183;
  reg [31:0] p1_smul_76184;
  reg [31:0] p1_smul_76185;
  reg [31:0] p1_smul_76186;
  reg [31:0] p1_smul_76187;
  reg [31:0] p1_smul_76188;
  reg [31:0] p1_smul_76189;
  reg [31:0] p1_smul_76190;
  reg [31:0] p1_smul_76191;
  reg [31:0] p1_smul_76192;
  reg [31:0] p1_smul_76193;
  reg [31:0] p1_smul_76194;
  reg [31:0] p1_smul_76195;
  reg [31:0] p1_smul_76196;
  reg [31:0] p1_smul_76197;
  reg [31:0] p1_smul_76198;
  reg [31:0] p1_smul_76199;
  reg [31:0] p1_smul_76200;
  reg [31:0] p1_smul_76201;
  reg [31:0] p1_smul_76202;
  reg [31:0] p1_smul_76203;
  reg [31:0] p1_smul_76204;
  reg [31:0] p1_smul_76205;
  reg [31:0] p1_smul_76206;
  reg [31:0] p1_smul_76207;
  reg [31:0] p1_smul_76208;
  reg [31:0] p1_smul_76209;
  reg [31:0] p1_smul_76210;
  reg [31:0] p1_smul_76211;
  reg [31:0] p1_smul_76212;
  reg [31:0] p1_smul_76213;
  reg [31:0] p1_smul_76214;
  reg [31:0] p1_smul_76215;
  reg [31:0] p1_smul_76216;
  reg [31:0] p1_smul_76217;
  reg [31:0] p1_smul_76218;
  reg [31:0] p1_smul_76219;
  reg [31:0] p1_smul_76220;
  reg [31:0] p1_smul_76221;
  reg [31:0] p1_smul_76222;
  reg [31:0] p1_smul_76223;
  reg [31:0] p1_smul_76224;
  reg [31:0] p1_smul_76225;
  reg [31:0] p1_smul_76226;
  reg [31:0] p1_smul_76227;
  reg [31:0] p1_smul_76228;
  reg [31:0] p1_smul_76229;
  reg [31:0] p1_smul_76230;
  reg [31:0] p1_smul_76231;
  reg [31:0] p1_smul_76232;
  reg [31:0] p1_smul_76233;
  reg [31:0] p1_smul_76234;
  reg [31:0] p1_smul_76235;
  reg [31:0] p1_smul_76236;
  reg [31:0] p1_smul_76237;
  reg [31:0] p1_smul_76238;
  reg [31:0] p1_smul_76239;
  reg [31:0] p1_smul_76240;
  reg [31:0] p1_smul_76241;
  reg [31:0] p1_smul_76242;
  reg [31:0] p1_smul_76243;
  reg [31:0] p1_smul_76244;
  reg [31:0] p1_smul_76245;
  reg [31:0] p1_smul_76246;
  reg [31:0] p1_smul_76247;
  reg [31:0] p1_smul_76248;
  reg [31:0] p1_smul_76249;
  reg [31:0] p1_smul_76250;
  reg [31:0] p1_smul_76251;
  reg [31:0] p1_smul_76252;
  reg [31:0] p1_smul_76253;
  reg [31:0] p1_smul_76254;
  reg [31:0] p1_smul_76255;
  reg [31:0] p1_smul_76256;
  reg [31:0] p1_smul_76257;
  reg [31:0] p1_smul_76258;
  reg [31:0] p1_smul_76259;
  reg [31:0] p1_smul_76260;
  reg [31:0] p1_smul_76261;
  reg [31:0] p1_smul_76262;
  reg [31:0] p1_smul_76263;
  reg [31:0] p1_smul_76264;
  reg [31:0] p1_smul_76265;
  reg [31:0] p1_smul_76266;
  reg [31:0] p1_smul_76267;
  reg [31:0] p1_smul_76268;
  reg [31:0] p1_smul_76269;
  reg [31:0] p1_smul_76270;
  reg [31:0] p1_smul_76271;
  reg [31:0] p1_smul_76272;
  reg [31:0] p1_smul_76273;
  reg [31:0] p1_smul_76274;
  reg [31:0] p1_smul_76275;
  reg [31:0] p1_smul_76276;
  reg [31:0] p1_smul_76277;
  reg [31:0] p1_smul_76278;
  reg [31:0] p1_smul_76279;
  reg [31:0] p1_smul_76280;
  reg [31:0] p1_smul_76281;
  reg [31:0] p1_smul_76282;
  reg [31:0] p1_smul_76283;
  reg [31:0] p1_smul_76284;
  reg [31:0] p1_smul_76285;
  reg [31:0] p1_smul_76286;
  reg [31:0] p1_smul_76287;
  reg [31:0] p1_smul_76288;
  reg [31:0] p1_smul_76289;
  reg [31:0] p1_smul_76290;
  reg [31:0] p1_smul_76291;
  reg [31:0] p1_smul_76292;
  reg [31:0] p1_smul_76293;
  reg [31:0] p1_smul_76294;
  reg [31:0] p1_smul_76295;
  reg [31:0] p1_smul_76296;
  reg [31:0] p1_smul_76297;
  reg [31:0] p1_smul_76298;
  reg [31:0] p1_smul_76299;
  reg [31:0] p1_smul_76300;
  reg [31:0] p1_smul_76301;
  reg [31:0] p1_smul_76302;
  reg [31:0] p1_smul_76303;
  reg [31:0] p1_smul_76304;
  reg [31:0] p1_smul_76305;
  reg [31:0] p1_smul_76306;
  reg [31:0] p1_smul_76307;
  reg [31:0] p1_smul_76308;
  reg [31:0] p1_smul_76309;
  reg [31:0] p1_smul_76310;
  reg [31:0] p1_smul_76311;
  reg [31:0] p1_smul_76312;
  reg [31:0] p1_smul_76313;
  reg [31:0] p1_smul_76314;
  reg [31:0] p1_smul_76315;
  reg [31:0] p1_smul_76316;
  reg [31:0] p1_smul_76317;
  reg [31:0] p1_smul_76318;
  reg [31:0] p1_smul_76319;
  reg [31:0] p1_smul_76320;
  reg [31:0] p1_smul_76321;
  reg [31:0] p1_smul_76322;
  reg [31:0] p1_smul_76323;
  reg [31:0] p1_smul_76324;
  reg [31:0] p1_smul_76325;
  reg [31:0] p1_smul_76326;
  reg [31:0] p1_smul_76327;
  reg [31:0] p1_smul_76328;
  reg [31:0] p1_smul_76329;
  reg [31:0] p1_smul_76330;
  reg [31:0] p1_smul_76331;
  reg [31:0] p1_smul_76332;
  reg [31:0] p1_smul_76333;
  reg [31:0] p1_smul_76334;
  reg [31:0] p1_smul_76335;
  reg [31:0] p1_smul_76336;
  reg [31:0] p1_smul_76337;
  reg [31:0] p1_smul_76338;
  reg [31:0] p1_smul_76339;
  reg [31:0] p1_smul_76340;
  reg [31:0] p1_smul_76341;
  reg [31:0] p1_smul_76342;
  reg [31:0] p1_smul_76343;
  reg [31:0] p1_smul_76344;
  reg [31:0] p1_smul_76345;
  reg [31:0] p1_smul_76346;
  reg [31:0] p1_smul_76347;
  reg [31:0] p1_smul_76348;
  reg [31:0] p1_smul_76349;
  reg [31:0] p1_smul_76350;
  reg [31:0] p1_smul_76351;
  reg [31:0] p1_smul_76352;
  reg [31:0] p1_smul_76353;
  reg [31:0] p1_smul_76354;
  reg [31:0] p1_smul_76355;
  reg [31:0] p1_smul_76356;
  reg [31:0] p1_smul_76357;
  reg [31:0] p1_smul_76358;
  reg [31:0] p1_smul_76359;
  reg [31:0] p1_smul_76360;
  reg [31:0] p1_smul_76361;
  reg [31:0] p1_smul_76362;
  reg [31:0] p1_smul_76363;
  reg [31:0] p1_smul_76364;
  reg [31:0] p1_smul_76365;
  reg [31:0] p1_smul_76366;
  reg [31:0] p1_smul_76367;
  reg [31:0] p1_smul_76368;
  reg [31:0] p1_smul_76369;
  reg [31:0] p1_smul_76370;
  reg [31:0] p1_smul_76371;
  reg [31:0] p1_smul_76372;
  reg [31:0] p1_smul_76373;
  reg [31:0] p1_smul_76374;
  reg [31:0] p1_smul_76375;
  reg [31:0] p1_smul_76376;
  reg [31:0] p1_smul_76377;
  reg [31:0] p1_smul_76378;
  reg [31:0] p1_smul_76379;
  reg [31:0] p1_smul_76380;
  reg [31:0] p1_smul_76381;
  reg [31:0] p1_smul_76382;
  reg [31:0] p1_smul_76383;
  reg [31:0] p1_smul_76384;
  reg [31:0] p1_smul_76385;
  reg [31:0] p1_smul_76386;
  reg [31:0] p1_smul_76387;
  reg [31:0] p1_smul_76388;
  reg [31:0] p1_smul_76389;
  reg [31:0] p1_smul_76390;
  reg [31:0] p1_smul_76391;
  reg [31:0] p1_smul_76392;
  reg [31:0] p1_smul_76393;
  reg [31:0] p1_smul_76394;
  reg [31:0] p1_smul_76395;
  reg [31:0] p1_smul_76396;
  reg [31:0] p1_smul_76397;
  reg [31:0] p1_smul_76398;
  reg [31:0] p1_smul_76399;
  reg [31:0] p1_smul_76400;
  reg [31:0] p1_smul_76401;
  reg [31:0] p1_smul_76402;
  reg [31:0] p1_smul_76403;
  reg [31:0] p1_smul_76404;
  reg [31:0] p1_smul_76405;
  reg [31:0] p1_smul_76406;
  reg [31:0] p1_smul_76407;
  reg [31:0] p1_smul_76408;
  reg [31:0] p1_smul_76409;
  reg [31:0] p1_smul_76410;
  reg [31:0] p1_smul_76411;
  reg [31:0] p1_smul_76412;
  reg [31:0] p1_smul_76413;
  reg [31:0] p1_smul_76414;
  reg [31:0] p1_smul_76415;
  reg [31:0] p1_smul_76416;
  reg [31:0] p1_smul_76417;
  reg [31:0] p1_smul_76418;
  reg [31:0] p1_smul_76419;
  reg [31:0] p1_smul_76420;
  reg [31:0] p1_smul_76421;
  reg [31:0] p1_smul_76422;
  reg [31:0] p1_smul_76423;
  reg [31:0] p1_smul_76424;
  reg [31:0] p1_smul_76425;
  reg [31:0] p1_smul_76426;
  reg [31:0] p1_smul_76427;
  reg [31:0] p1_smul_76428;
  reg [31:0] p1_smul_76429;
  reg [31:0] p1_smul_76430;
  reg [31:0] p1_smul_76431;
  reg [31:0] p1_smul_76432;
  reg [31:0] p1_smul_76433;
  reg [31:0] p1_smul_76434;
  reg [31:0] p1_smul_76435;
  reg [31:0] p1_smul_76436;
  reg [31:0] p1_smul_76437;
  reg [31:0] p1_smul_76438;
  reg [31:0] p1_smul_76439;
  reg [31:0] p1_smul_76440;
  reg [31:0] p1_smul_76441;
  reg [31:0] p1_smul_76442;
  reg [31:0] p1_smul_76443;
  reg [31:0] p1_smul_76444;
  reg [31:0] p1_smul_76445;
  reg [31:0] p1_smul_76446;
  reg [31:0] p1_smul_76447;
  reg [31:0] p1_smul_76448;
  reg [31:0] p1_smul_76449;
  reg [31:0] p1_smul_76450;
  reg [31:0] p1_smul_76451;
  reg [31:0] p1_smul_76452;
  reg [31:0] p1_smul_76453;
  reg [31:0] p1_smul_76454;
  reg [31:0] p1_smul_76455;
  reg [31:0] p1_smul_76456;
  reg [31:0] p1_smul_76457;
  reg [31:0] p1_smul_76458;
  reg [31:0] p1_smul_76459;
  reg [31:0] p1_smul_76460;
  reg [31:0] p1_smul_76461;
  reg [31:0] p1_smul_76462;
  reg [31:0] p1_smul_76463;
  reg [31:0] p1_smul_76464;
  reg [31:0] p1_smul_76465;
  reg [31:0] p1_smul_76466;
  reg [31:0] p1_smul_76467;
  reg [31:0] p1_smul_76468;
  reg [31:0] p1_smul_76469;
  reg [31:0] p1_smul_76470;
  reg [31:0] p1_smul_76471;
  reg [31:0] p1_smul_76472;
  reg [31:0] p1_smul_76473;
  reg [31:0] p1_smul_76474;
  reg [31:0] p1_smul_76475;
  reg [31:0] p1_smul_76476;
  reg [31:0] p1_smul_76477;
  reg [31:0] p1_smul_76478;
  reg [31:0] p1_smul_76479;
  reg [31:0] p1_smul_76480;
  reg [31:0] p1_smul_76481;
  reg [31:0] p1_smul_76482;
  reg [31:0] p1_smul_76483;
  reg [31:0] p1_smul_76484;
  reg [31:0] p1_smul_76485;
  reg [31:0] p1_smul_76486;
  reg [31:0] p1_smul_76487;
  reg [31:0] p1_smul_76488;
  reg [31:0] p1_smul_76489;
  reg [31:0] p1_smul_76490;
  reg [31:0] p1_smul_76491;
  reg [31:0] p1_smul_76492;
  reg [31:0] p1_smul_76493;
  reg [31:0] p1_smul_76494;
  reg [31:0] p1_smul_76495;
  reg [31:0] p1_smul_76496;
  reg [31:0] p1_smul_76497;
  reg [31:0] p1_smul_76498;
  reg [31:0] p1_smul_76499;
  reg [31:0] p1_smul_76500;
  reg [31:0] p1_smul_76501;
  reg [31:0] p1_smul_76502;
  reg [31:0] p1_smul_76503;
  reg [31:0] p1_smul_76504;
  reg [31:0] p1_smul_76505;
  reg [31:0] p1_smul_76506;
  reg [31:0] p1_smul_76507;
  reg [31:0] p1_smul_76508;
  reg [31:0] p1_smul_76509;
  reg [31:0] p1_smul_76510;
  reg [31:0] p1_smul_76511;
  reg [31:0] p1_smul_76512;
  reg [31:0] p1_smul_76513;
  reg [31:0] p1_smul_76514;
  reg [31:0] p1_smul_76515;
  reg [31:0] p1_smul_76516;
  reg [31:0] p1_smul_76517;
  reg [31:0] p1_smul_76518;
  reg [31:0] p1_smul_76519;
  reg [31:0] p1_smul_76520;
  reg [31:0] p1_smul_76521;
  reg [31:0] p1_smul_76522;
  reg [31:0] p1_smul_76523;
  reg [31:0] p1_smul_76524;
  reg [31:0] p1_smul_76525;
  reg [31:0] p1_smul_76526;
  reg [31:0] p1_smul_76527;
  reg [31:0] p1_smul_76528;
  reg [31:0] p1_smul_76529;
  reg [31:0] p1_smul_76530;
  reg [31:0] p1_smul_76531;
  reg [31:0] p1_smul_76532;
  reg [31:0] p1_smul_76533;
  reg [31:0] p1_smul_76534;
  reg [31:0] p1_smul_76535;
  reg [31:0] p1_smul_76536;
  reg [31:0] p1_smul_76537;
  reg [31:0] p1_smul_76538;
  reg [31:0] p1_smul_76539;
  reg [31:0] p1_smul_76540;
  reg [31:0] p1_smul_76541;
  reg [31:0] p1_smul_76542;
  reg [31:0] p1_smul_76543;
  reg [31:0] p1_smul_76544;
  reg [31:0] p1_smul_76545;
  reg [31:0] p1_smul_76546;
  reg [31:0] p1_smul_76547;
  reg [31:0] p1_smul_76548;
  reg [31:0] p1_smul_76549;
  reg [31:0] p1_smul_76550;
  reg [31:0] p1_smul_76551;
  reg [31:0] p1_smul_76552;
  reg [31:0] p1_smul_76553;
  reg [31:0] p1_smul_76554;
  reg [31:0] p1_smul_76555;
  reg [31:0] p1_smul_76556;
  reg [31:0] p1_smul_76557;
  reg [31:0] p1_smul_76558;
  reg [31:0] p1_smul_76559;
  reg [31:0] p1_smul_76560;
  reg [31:0] p1_smul_76561;
  reg [31:0] p1_smul_76562;
  reg [31:0] p1_smul_76563;
  reg [31:0] p1_smul_76564;
  reg [31:0] p1_smul_76565;
  reg [31:0] p1_smul_76566;
  reg [31:0] p1_smul_76567;
  reg [31:0] p1_smul_76568;
  reg [31:0] p1_smul_76569;
  reg [31:0] p1_smul_76570;
  reg [31:0] p1_smul_76571;
  reg [31:0] p1_smul_76572;
  reg [31:0] p1_smul_76573;
  reg [31:0] p1_smul_76574;
  reg [31:0] p1_smul_76575;
  reg [31:0] p1_smul_76576;
  reg [31:0] p1_smul_76577;
  reg [31:0] p1_smul_76578;
  reg [31:0] p1_smul_76579;
  reg [31:0] p1_smul_76580;
  reg [31:0] p1_smul_76581;
  reg [31:0] p1_smul_76582;
  reg [31:0] p1_smul_76583;
  reg [31:0] p1_smul_76584;
  reg [31:0] p1_smul_76585;
  reg [31:0] p1_smul_76586;
  reg [31:0] p1_smul_76587;
  reg [31:0] p1_smul_76588;
  reg [31:0] p1_smul_76589;
  reg [31:0] p1_smul_76590;
  reg [31:0] p1_smul_76591;
  reg [31:0] p1_smul_76592;
  reg [31:0] p1_smul_76593;
  reg [31:0] p1_smul_76594;
  reg [31:0] p1_smul_76595;
  reg [31:0] p1_smul_76596;
  reg [31:0] p1_smul_76597;
  reg [31:0] p1_smul_76598;
  reg [31:0] p1_smul_76599;
  reg [31:0] p1_smul_76600;
  reg [31:0] p1_smul_76601;
  reg [31:0] p1_smul_76602;
  reg [31:0] p1_smul_76603;
  reg [31:0] p1_smul_76604;
  reg [31:0] p1_smul_76605;
  reg [31:0] p1_smul_76606;
  reg [31:0] p1_smul_76607;
  reg [31:0] p1_smul_76608;
  reg [31:0] p1_smul_76609;
  reg [31:0] p1_smul_76610;
  reg [31:0] p1_smul_76611;
  reg [31:0] p1_smul_76612;
  reg [31:0] p1_smul_76613;
  reg [31:0] p1_smul_76614;
  reg [31:0] p1_smul_76615;
  reg [31:0] p1_smul_76616;
  reg [31:0] p1_smul_76617;
  reg [31:0] p1_smul_76618;
  reg [31:0] p1_smul_76619;
  reg [31:0] p1_smul_76620;
  reg [31:0] p1_smul_76621;
  reg [31:0] p1_smul_76622;
  reg [31:0] p1_smul_76623;
  reg [31:0] p1_smul_76624;
  reg [31:0] p1_smul_76625;
  reg [31:0] p1_smul_76626;
  reg [31:0] p1_smul_76627;
  reg [31:0] p1_smul_76628;
  reg [31:0] p1_smul_76629;
  reg [31:0] p1_smul_76630;
  reg [31:0] p1_smul_76631;
  reg [31:0] p1_smul_76632;
  reg [31:0] p1_smul_76633;
  reg [31:0] p1_smul_76634;
  reg [31:0] p1_smul_76635;
  reg [31:0] p1_smul_76636;
  reg [31:0] p1_smul_76637;
  reg [31:0] p1_smul_76638;
  reg [31:0] p1_smul_76639;
  reg [31:0] p1_smul_76640;
  reg [31:0] p1_smul_76641;
  reg [31:0] p1_smul_76642;
  reg [31:0] p1_smul_76643;
  reg [31:0] p1_smul_76644;
  reg [31:0] p1_smul_76645;
  reg [31:0] p1_smul_76646;
  reg [31:0] p1_smul_76647;
  reg [31:0] p1_smul_76648;
  reg [31:0] p1_smul_76649;
  reg [31:0] p1_smul_76650;
  reg [31:0] p1_smul_76651;
  reg [31:0] p1_smul_76652;
  reg [31:0] p1_smul_76653;
  reg [31:0] p1_smul_76654;
  reg [31:0] p1_smul_76655;
  reg [31:0] p1_smul_76656;
  reg [31:0] p1_smul_76657;
  reg [31:0] p1_smul_76658;
  reg [31:0] p1_smul_76659;
  reg [31:0] p1_smul_76660;
  reg [31:0] p1_smul_76661;
  reg [31:0] p1_smul_76662;
  reg [31:0] p1_smul_76663;
  reg [31:0] p1_smul_76664;
  reg [31:0] p1_smul_76665;
  reg [31:0] p1_smul_76666;
  reg [31:0] p1_smul_76667;
  reg [31:0] p1_smul_76668;
  reg [31:0] p1_smul_76669;
  reg [31:0] p1_smul_76670;
  reg [31:0] p1_smul_76671;
  reg [31:0] p1_smul_76672;
  reg [31:0] p1_smul_76673;
  reg [31:0] p1_smul_76674;
  reg [31:0] p1_smul_76675;
  reg [31:0] p1_smul_76676;
  reg [31:0] p1_smul_76677;
  reg [31:0] p1_smul_76678;
  reg [31:0] p1_smul_76679;
  reg [31:0] p1_smul_76680;
  reg [31:0] p1_smul_76681;
  reg [31:0] p1_smul_76682;
  reg [31:0] p1_smul_76683;
  reg [31:0] p1_smul_76684;
  reg [31:0] p1_smul_76685;
  reg [31:0] p1_smul_76686;
  reg [31:0] p1_smul_76687;
  reg [31:0] p1_smul_76688;
  reg [31:0] p1_smul_76689;
  reg [31:0] p1_smul_76690;
  reg [31:0] p1_smul_76691;
  reg [31:0] p1_smul_76692;
  reg [31:0] p1_smul_76693;
  reg [31:0] p1_smul_76694;
  reg [31:0] p1_smul_76695;
  reg [31:0] p1_smul_76696;
  reg [31:0] p1_smul_76697;
  reg [31:0] p1_smul_76698;
  reg [31:0] p1_smul_76699;
  reg [31:0] p1_smul_76700;
  reg [31:0] p1_smul_76701;
  reg [31:0] p1_smul_76702;
  reg [31:0] p1_smul_76703;
  reg [31:0] p1_smul_76704;
  reg [31:0] p1_smul_76705;
  reg [31:0] p1_smul_76706;
  reg [31:0] p1_smul_76707;
  reg [31:0] p1_smul_76708;
  reg [31:0] p1_smul_76709;
  reg [31:0] p1_smul_76710;
  reg [31:0] p1_smul_76711;
  reg [31:0] p1_smul_76712;
  reg [31:0] p1_smul_76713;
  reg [31:0] p1_smul_76714;
  reg [31:0] p1_smul_76715;
  reg [31:0] p1_smul_76716;
  reg [31:0] p1_smul_76717;
  reg [31:0] p1_smul_76718;
  reg [31:0] p1_smul_76719;
  reg [31:0] p1_smul_76720;
  reg [31:0] p1_smul_76721;
  reg [31:0] p1_smul_76722;
  reg [31:0] p1_smul_76723;
  reg [31:0] p1_smul_76724;
  reg [31:0] p1_smul_76725;
  reg [31:0] p1_smul_76726;
  reg [31:0] p1_smul_76727;
  reg [31:0] p1_smul_76728;
  reg [31:0] p1_smul_76729;
  reg [31:0] p1_smul_76730;
  reg [31:0] p1_smul_76731;
  reg [31:0] p1_smul_76732;
  reg [31:0] p1_smul_76733;
  reg [31:0] p1_smul_76734;
  reg [31:0] p1_smul_76735;
  reg [31:0] p1_smul_76736;
  reg [31:0] p1_smul_76737;
  reg [31:0] p1_smul_76738;
  reg [31:0] p1_smul_76739;
  reg [31:0] p1_smul_76740;
  reg [31:0] p1_smul_76741;
  reg [31:0] p1_smul_76742;
  reg [31:0] p1_smul_76743;
  reg [31:0] p1_smul_76744;
  reg [31:0] p1_smul_76745;
  reg [31:0] p1_smul_76746;
  reg [31:0] p1_smul_76747;
  reg [31:0] p1_smul_76748;
  reg [31:0] p1_smul_76749;
  reg [31:0] p1_smul_76750;
  reg [31:0] p1_smul_76751;
  reg [31:0] p1_smul_76752;
  reg [31:0] p1_smul_76753;
  reg [31:0] p1_smul_76754;
  reg [31:0] p1_smul_76755;
  reg [31:0] p1_smul_76756;
  reg [31:0] p1_smul_76757;
  reg [31:0] p1_smul_76758;
  reg [31:0] p1_smul_76759;
  reg [31:0] p1_smul_76760;
  reg [31:0] p1_smul_76761;
  reg [31:0] p1_smul_76762;
  reg [31:0] p1_smul_76763;
  reg [31:0] p1_smul_76764;
  reg [31:0] p1_smul_76765;
  reg [31:0] p1_smul_76766;
  reg [31:0] p1_smul_76767;
  reg [31:0] p1_smul_76768;
  reg [31:0] p1_smul_76769;
  reg [31:0] p1_smul_76770;
  reg [31:0] p1_smul_76771;
  reg [31:0] p1_smul_76772;
  reg [31:0] p1_smul_76773;
  reg [31:0] p1_smul_76774;
  reg [31:0] p1_smul_76775;
  reg [31:0] p1_smul_76776;
  reg [31:0] p1_smul_76777;
  reg [31:0] p1_smul_76778;
  reg [31:0] p1_smul_76779;
  reg [31:0] p1_smul_76780;
  reg [31:0] p1_smul_76781;
  reg [31:0] p1_smul_76782;
  reg [31:0] p1_smul_76783;
  reg [31:0] p1_smul_76784;
  reg [31:0] p1_smul_76785;
  reg [31:0] p1_smul_76786;
  reg [31:0] p1_smul_76787;
  reg [31:0] p1_smul_76788;
  reg [31:0] p1_smul_76789;
  reg [31:0] p1_smul_76790;
  reg [31:0] p1_smul_76791;
  reg [31:0] p1_smul_76792;
  reg [31:0] p1_smul_76793;
  reg [31:0] p1_smul_76794;
  reg [31:0] p1_smul_76795;
  reg [31:0] p1_smul_76796;
  reg [31:0] p1_smul_76797;
  reg [31:0] p1_smul_76798;
  reg [31:0] p1_smul_76799;
  reg [31:0] p1_smul_76800;
  reg [31:0] p1_smul_76801;
  reg [31:0] p1_smul_76802;
  reg [31:0] p1_smul_76803;
  reg [31:0] p1_smul_76804;
  reg [31:0] p1_smul_76805;
  reg [31:0] p1_smul_76806;
  reg [31:0] p1_smul_76807;
  reg [31:0] p1_smul_76808;
  reg [31:0] p1_smul_76809;
  reg [31:0] p1_smul_76810;
  reg [31:0] p1_smul_76811;
  reg [31:0] p1_smul_76812;
  reg [31:0] p1_smul_76813;
  reg [31:0] p1_smul_76814;
  reg [31:0] p1_smul_76815;
  reg [31:0] p1_smul_76816;
  reg [31:0] p1_smul_76817;
  reg [31:0] p1_smul_76818;
  reg [31:0] p1_smul_76819;
  reg [31:0] p1_smul_76820;
  reg [31:0] p1_smul_76821;
  reg [31:0] p1_smul_76822;
  reg [31:0] p1_smul_76823;
  reg [31:0] p1_smul_76824;
  reg [31:0] p1_smul_76825;
  reg [31:0] p1_smul_76826;
  reg [31:0] p1_smul_76827;
  reg [31:0] p1_smul_76828;
  reg [31:0] p1_smul_76829;
  reg [31:0] p1_smul_76830;
  reg [31:0] p1_smul_76831;
  reg [31:0] p1_smul_76832;
  reg [31:0] p1_smul_76833;
  reg [31:0] p1_smul_76834;
  reg [31:0] p1_smul_76835;
  reg [31:0] p1_smul_76836;
  reg [31:0] p1_smul_76837;
  reg [31:0] p1_smul_76838;
  reg [31:0] p1_smul_76839;
  reg [31:0] p1_smul_76840;
  reg [31:0] p1_smul_76841;
  reg [31:0] p1_smul_76842;
  reg [31:0] p1_smul_76843;
  reg [31:0] p1_smul_76844;
  reg [31:0] p1_smul_76845;
  reg [31:0] p1_smul_76846;
  reg [31:0] p1_smul_76847;
  reg [31:0] p1_smul_76848;
  reg [31:0] p1_smul_76849;
  reg [31:0] p1_smul_76850;
  reg [31:0] p1_smul_76851;
  reg [31:0] p1_smul_76852;
  reg [31:0] p1_smul_76853;
  reg [31:0] p1_smul_76854;
  reg [31:0] p1_smul_76855;
  reg [31:0] p1_smul_76856;
  reg [31:0] p1_smul_76857;
  reg [31:0] p1_smul_76858;
  reg [31:0] p1_smul_76859;
  reg [31:0] p1_smul_76860;
  reg [31:0] p1_smul_76861;
  reg [31:0] p1_smul_76862;
  reg [31:0] p1_smul_76863;
  reg [31:0] p1_smul_76864;
  reg [31:0] p1_smul_76865;
  reg [31:0] p1_smul_76866;
  reg [31:0] p1_smul_76867;
  reg [31:0] p1_smul_76868;
  reg [31:0] p1_smul_76869;
  reg [31:0] p1_smul_76870;
  reg [31:0] p1_smul_76871;
  reg [31:0] p1_smul_76872;
  reg [31:0] p1_smul_76873;
  reg [31:0] p1_smul_76874;
  reg [31:0] p1_smul_76875;
  reg [31:0] p1_smul_76876;
  reg [31:0] p1_smul_76877;
  reg [31:0] p1_smul_76878;
  reg [31:0] p1_smul_76879;
  reg [31:0] p1_smul_76880;
  reg [31:0] p1_smul_76881;
  reg [31:0] p1_smul_76882;
  reg [31:0] p1_smul_76883;
  reg [31:0] p1_smul_76884;
  reg [31:0] p1_smul_76885;
  reg [31:0] p1_smul_76886;
  reg [31:0] p1_smul_76887;
  reg [31:0] p1_smul_76888;
  reg [31:0] p1_smul_76889;
  reg [31:0] p1_smul_76890;
  reg [31:0] p1_smul_76891;
  reg [31:0] p1_smul_76892;
  reg [31:0] p1_smul_76893;
  reg [31:0] p1_smul_76894;
  reg [31:0] p1_smul_76895;
  reg [31:0] p1_smul_76896;
  reg [31:0] p1_smul_76897;
  reg [31:0] p1_smul_76898;
  reg [31:0] p1_smul_76899;
  reg [31:0] p1_smul_76900;
  reg [31:0] p1_smul_76901;
  reg [31:0] p1_smul_76902;
  reg [31:0] p1_smul_76903;
  reg [31:0] p1_smul_76904;
  reg [31:0] p1_smul_76905;
  reg [31:0] p1_smul_76906;
  reg [31:0] p1_smul_76907;
  reg [31:0] p1_smul_76908;
  reg [31:0] p1_smul_76909;
  reg [31:0] p1_smul_76910;
  reg [31:0] p1_smul_76911;
  reg [31:0] p1_smul_76912;
  reg [31:0] p1_smul_76913;
  reg [31:0] p1_smul_76914;
  reg [31:0] p1_smul_76915;
  reg [31:0] p1_smul_76916;
  reg [31:0] p1_smul_76917;
  reg [31:0] p1_smul_76918;
  reg [31:0] p1_smul_76919;
  reg [31:0] p1_smul_76920;
  reg [31:0] p1_smul_76921;
  reg [31:0] p1_smul_76922;
  reg [31:0] p1_smul_76923;
  reg [31:0] p1_smul_76924;
  reg [31:0] p1_smul_76925;
  reg [31:0] p1_smul_76926;
  reg [31:0] p1_smul_76927;
  reg [31:0] p1_smul_76928;
  reg [31:0] p1_smul_76929;
  reg [31:0] p1_smul_76930;
  reg [31:0] p1_smul_76931;
  reg [31:0] p1_smul_76932;
  reg [31:0] p1_smul_76933;
  reg [31:0] p1_smul_76934;
  reg [31:0] p1_smul_76935;
  reg [31:0] p1_smul_76936;
  reg [31:0] p1_smul_76937;
  reg [31:0] p1_smul_76938;
  reg [31:0] p1_smul_76939;
  reg [31:0] p1_smul_76940;
  reg [31:0] p1_smul_76941;
  reg [31:0] p1_smul_76942;
  reg [31:0] p1_smul_76943;
  reg [31:0] p1_smul_76944;
  reg [31:0] p1_smul_76945;
  reg [31:0] p1_smul_76946;
  reg [31:0] p1_smul_76947;
  reg [31:0] p1_smul_76948;
  reg [31:0] p1_smul_76949;
  reg [31:0] p1_smul_76950;
  reg [31:0] p1_smul_76951;
  reg [31:0] p1_smul_76952;
  reg [31:0] p1_smul_76953;
  reg [31:0] p1_smul_76954;
  reg [31:0] p1_smul_76955;
  reg [31:0] p1_smul_76956;
  reg [31:0] p1_smul_76957;
  reg [31:0] p1_smul_76958;
  reg [31:0] p1_smul_76959;
  reg [31:0] p1_smul_76960;
  reg [31:0] p1_smul_76961;
  reg [31:0] p1_smul_76962;
  reg [31:0] p1_smul_76963;
  reg [31:0] p1_smul_76964;
  reg [31:0] p1_smul_76965;
  reg [31:0] p1_smul_76966;
  reg [31:0] p1_smul_76967;
  reg [31:0] p1_smul_76968;
  reg [31:0] p1_smul_76969;
  reg [31:0] p1_smul_76970;
  reg [31:0] p1_smul_76971;
  always_ff @ (posedge clk) begin
    p1_smul_75972 <= p1_smul_75972_comb;
    p1_smul_75973 <= p1_smul_75973_comb;
    p1_smul_75974 <= p1_smul_75974_comb;
    p1_smul_75975 <= p1_smul_75975_comb;
    p1_smul_75976 <= p1_smul_75976_comb;
    p1_smul_75977 <= p1_smul_75977_comb;
    p1_smul_75978 <= p1_smul_75978_comb;
    p1_smul_75979 <= p1_smul_75979_comb;
    p1_smul_75980 <= p1_smul_75980_comb;
    p1_smul_75981 <= p1_smul_75981_comb;
    p1_smul_75982 <= p1_smul_75982_comb;
    p1_smul_75983 <= p1_smul_75983_comb;
    p1_smul_75984 <= p1_smul_75984_comb;
    p1_smul_75985 <= p1_smul_75985_comb;
    p1_smul_75986 <= p1_smul_75986_comb;
    p1_smul_75987 <= p1_smul_75987_comb;
    p1_smul_75988 <= p1_smul_75988_comb;
    p1_smul_75989 <= p1_smul_75989_comb;
    p1_smul_75990 <= p1_smul_75990_comb;
    p1_smul_75991 <= p1_smul_75991_comb;
    p1_smul_75992 <= p1_smul_75992_comb;
    p1_smul_75993 <= p1_smul_75993_comb;
    p1_smul_75994 <= p1_smul_75994_comb;
    p1_smul_75995 <= p1_smul_75995_comb;
    p1_smul_75996 <= p1_smul_75996_comb;
    p1_smul_75997 <= p1_smul_75997_comb;
    p1_smul_75998 <= p1_smul_75998_comb;
    p1_smul_75999 <= p1_smul_75999_comb;
    p1_smul_76000 <= p1_smul_76000_comb;
    p1_smul_76001 <= p1_smul_76001_comb;
    p1_smul_76002 <= p1_smul_76002_comb;
    p1_smul_76003 <= p1_smul_76003_comb;
    p1_smul_76004 <= p1_smul_76004_comb;
    p1_smul_76005 <= p1_smul_76005_comb;
    p1_smul_76006 <= p1_smul_76006_comb;
    p1_smul_76007 <= p1_smul_76007_comb;
    p1_smul_76008 <= p1_smul_76008_comb;
    p1_smul_76009 <= p1_smul_76009_comb;
    p1_smul_76010 <= p1_smul_76010_comb;
    p1_smul_76011 <= p1_smul_76011_comb;
    p1_smul_76012 <= p1_smul_76012_comb;
    p1_smul_76013 <= p1_smul_76013_comb;
    p1_smul_76014 <= p1_smul_76014_comb;
    p1_smul_76015 <= p1_smul_76015_comb;
    p1_smul_76016 <= p1_smul_76016_comb;
    p1_smul_76017 <= p1_smul_76017_comb;
    p1_smul_76018 <= p1_smul_76018_comb;
    p1_smul_76019 <= p1_smul_76019_comb;
    p1_smul_76020 <= p1_smul_76020_comb;
    p1_smul_76021 <= p1_smul_76021_comb;
    p1_smul_76022 <= p1_smul_76022_comb;
    p1_smul_76023 <= p1_smul_76023_comb;
    p1_smul_76024 <= p1_smul_76024_comb;
    p1_smul_76025 <= p1_smul_76025_comb;
    p1_smul_76026 <= p1_smul_76026_comb;
    p1_smul_76027 <= p1_smul_76027_comb;
    p1_smul_76028 <= p1_smul_76028_comb;
    p1_smul_76029 <= p1_smul_76029_comb;
    p1_smul_76030 <= p1_smul_76030_comb;
    p1_smul_76031 <= p1_smul_76031_comb;
    p1_smul_76032 <= p1_smul_76032_comb;
    p1_smul_76033 <= p1_smul_76033_comb;
    p1_smul_76034 <= p1_smul_76034_comb;
    p1_smul_76035 <= p1_smul_76035_comb;
    p1_smul_76036 <= p1_smul_76036_comb;
    p1_smul_76037 <= p1_smul_76037_comb;
    p1_smul_76038 <= p1_smul_76038_comb;
    p1_smul_76039 <= p1_smul_76039_comb;
    p1_smul_76040 <= p1_smul_76040_comb;
    p1_smul_76041 <= p1_smul_76041_comb;
    p1_smul_76042 <= p1_smul_76042_comb;
    p1_smul_76043 <= p1_smul_76043_comb;
    p1_smul_76044 <= p1_smul_76044_comb;
    p1_smul_76045 <= p1_smul_76045_comb;
    p1_smul_76046 <= p1_smul_76046_comb;
    p1_smul_76047 <= p1_smul_76047_comb;
    p1_smul_76048 <= p1_smul_76048_comb;
    p1_smul_76049 <= p1_smul_76049_comb;
    p1_smul_76050 <= p1_smul_76050_comb;
    p1_smul_76051 <= p1_smul_76051_comb;
    p1_smul_76052 <= p1_smul_76052_comb;
    p1_smul_76053 <= p1_smul_76053_comb;
    p1_smul_76054 <= p1_smul_76054_comb;
    p1_smul_76055 <= p1_smul_76055_comb;
    p1_smul_76056 <= p1_smul_76056_comb;
    p1_smul_76057 <= p1_smul_76057_comb;
    p1_smul_76058 <= p1_smul_76058_comb;
    p1_smul_76059 <= p1_smul_76059_comb;
    p1_smul_76060 <= p1_smul_76060_comb;
    p1_smul_76061 <= p1_smul_76061_comb;
    p1_smul_76062 <= p1_smul_76062_comb;
    p1_smul_76063 <= p1_smul_76063_comb;
    p1_smul_76064 <= p1_smul_76064_comb;
    p1_smul_76065 <= p1_smul_76065_comb;
    p1_smul_76066 <= p1_smul_76066_comb;
    p1_smul_76067 <= p1_smul_76067_comb;
    p1_smul_76068 <= p1_smul_76068_comb;
    p1_smul_76069 <= p1_smul_76069_comb;
    p1_smul_76070 <= p1_smul_76070_comb;
    p1_smul_76071 <= p1_smul_76071_comb;
    p1_smul_76072 <= p1_smul_76072_comb;
    p1_smul_76073 <= p1_smul_76073_comb;
    p1_smul_76074 <= p1_smul_76074_comb;
    p1_smul_76075 <= p1_smul_76075_comb;
    p1_smul_76076 <= p1_smul_76076_comb;
    p1_smul_76077 <= p1_smul_76077_comb;
    p1_smul_76078 <= p1_smul_76078_comb;
    p1_smul_76079 <= p1_smul_76079_comb;
    p1_smul_76080 <= p1_smul_76080_comb;
    p1_smul_76081 <= p1_smul_76081_comb;
    p1_smul_76082 <= p1_smul_76082_comb;
    p1_smul_76083 <= p1_smul_76083_comb;
    p1_smul_76084 <= p1_smul_76084_comb;
    p1_smul_76085 <= p1_smul_76085_comb;
    p1_smul_76086 <= p1_smul_76086_comb;
    p1_smul_76087 <= p1_smul_76087_comb;
    p1_smul_76088 <= p1_smul_76088_comb;
    p1_smul_76089 <= p1_smul_76089_comb;
    p1_smul_76090 <= p1_smul_76090_comb;
    p1_smul_76091 <= p1_smul_76091_comb;
    p1_smul_76092 <= p1_smul_76092_comb;
    p1_smul_76093 <= p1_smul_76093_comb;
    p1_smul_76094 <= p1_smul_76094_comb;
    p1_smul_76095 <= p1_smul_76095_comb;
    p1_smul_76096 <= p1_smul_76096_comb;
    p1_smul_76097 <= p1_smul_76097_comb;
    p1_smul_76098 <= p1_smul_76098_comb;
    p1_smul_76099 <= p1_smul_76099_comb;
    p1_smul_76100 <= p1_smul_76100_comb;
    p1_smul_76101 <= p1_smul_76101_comb;
    p1_smul_76102 <= p1_smul_76102_comb;
    p1_smul_76103 <= p1_smul_76103_comb;
    p1_smul_76104 <= p1_smul_76104_comb;
    p1_smul_76105 <= p1_smul_76105_comb;
    p1_smul_76106 <= p1_smul_76106_comb;
    p1_smul_76107 <= p1_smul_76107_comb;
    p1_smul_76108 <= p1_smul_76108_comb;
    p1_smul_76109 <= p1_smul_76109_comb;
    p1_smul_76110 <= p1_smul_76110_comb;
    p1_smul_76111 <= p1_smul_76111_comb;
    p1_smul_76112 <= p1_smul_76112_comb;
    p1_smul_76113 <= p1_smul_76113_comb;
    p1_smul_76114 <= p1_smul_76114_comb;
    p1_smul_76115 <= p1_smul_76115_comb;
    p1_smul_76116 <= p1_smul_76116_comb;
    p1_smul_76117 <= p1_smul_76117_comb;
    p1_smul_76118 <= p1_smul_76118_comb;
    p1_smul_76119 <= p1_smul_76119_comb;
    p1_smul_76120 <= p1_smul_76120_comb;
    p1_smul_76121 <= p1_smul_76121_comb;
    p1_smul_76122 <= p1_smul_76122_comb;
    p1_smul_76123 <= p1_smul_76123_comb;
    p1_smul_76124 <= p1_smul_76124_comb;
    p1_smul_76125 <= p1_smul_76125_comb;
    p1_smul_76126 <= p1_smul_76126_comb;
    p1_smul_76127 <= p1_smul_76127_comb;
    p1_smul_76128 <= p1_smul_76128_comb;
    p1_smul_76129 <= p1_smul_76129_comb;
    p1_smul_76130 <= p1_smul_76130_comb;
    p1_smul_76131 <= p1_smul_76131_comb;
    p1_smul_76132 <= p1_smul_76132_comb;
    p1_smul_76133 <= p1_smul_76133_comb;
    p1_smul_76134 <= p1_smul_76134_comb;
    p1_smul_76135 <= p1_smul_76135_comb;
    p1_smul_76136 <= p1_smul_76136_comb;
    p1_smul_76137 <= p1_smul_76137_comb;
    p1_smul_76138 <= p1_smul_76138_comb;
    p1_smul_76139 <= p1_smul_76139_comb;
    p1_smul_76140 <= p1_smul_76140_comb;
    p1_smul_76141 <= p1_smul_76141_comb;
    p1_smul_76142 <= p1_smul_76142_comb;
    p1_smul_76143 <= p1_smul_76143_comb;
    p1_smul_76144 <= p1_smul_76144_comb;
    p1_smul_76145 <= p1_smul_76145_comb;
    p1_smul_76146 <= p1_smul_76146_comb;
    p1_smul_76147 <= p1_smul_76147_comb;
    p1_smul_76148 <= p1_smul_76148_comb;
    p1_smul_76149 <= p1_smul_76149_comb;
    p1_smul_76150 <= p1_smul_76150_comb;
    p1_smul_76151 <= p1_smul_76151_comb;
    p1_smul_76152 <= p1_smul_76152_comb;
    p1_smul_76153 <= p1_smul_76153_comb;
    p1_smul_76154 <= p1_smul_76154_comb;
    p1_smul_76155 <= p1_smul_76155_comb;
    p1_smul_76156 <= p1_smul_76156_comb;
    p1_smul_76157 <= p1_smul_76157_comb;
    p1_smul_76158 <= p1_smul_76158_comb;
    p1_smul_76159 <= p1_smul_76159_comb;
    p1_smul_76160 <= p1_smul_76160_comb;
    p1_smul_76161 <= p1_smul_76161_comb;
    p1_smul_76162 <= p1_smul_76162_comb;
    p1_smul_76163 <= p1_smul_76163_comb;
    p1_smul_76164 <= p1_smul_76164_comb;
    p1_smul_76165 <= p1_smul_76165_comb;
    p1_smul_76166 <= p1_smul_76166_comb;
    p1_smul_76167 <= p1_smul_76167_comb;
    p1_smul_76168 <= p1_smul_76168_comb;
    p1_smul_76169 <= p1_smul_76169_comb;
    p1_smul_76170 <= p1_smul_76170_comb;
    p1_smul_76171 <= p1_smul_76171_comb;
    p1_smul_76172 <= p1_smul_76172_comb;
    p1_smul_76173 <= p1_smul_76173_comb;
    p1_smul_76174 <= p1_smul_76174_comb;
    p1_smul_76175 <= p1_smul_76175_comb;
    p1_smul_76176 <= p1_smul_76176_comb;
    p1_smul_76177 <= p1_smul_76177_comb;
    p1_smul_76178 <= p1_smul_76178_comb;
    p1_smul_76179 <= p1_smul_76179_comb;
    p1_smul_76180 <= p1_smul_76180_comb;
    p1_smul_76181 <= p1_smul_76181_comb;
    p1_smul_76182 <= p1_smul_76182_comb;
    p1_smul_76183 <= p1_smul_76183_comb;
    p1_smul_76184 <= p1_smul_76184_comb;
    p1_smul_76185 <= p1_smul_76185_comb;
    p1_smul_76186 <= p1_smul_76186_comb;
    p1_smul_76187 <= p1_smul_76187_comb;
    p1_smul_76188 <= p1_smul_76188_comb;
    p1_smul_76189 <= p1_smul_76189_comb;
    p1_smul_76190 <= p1_smul_76190_comb;
    p1_smul_76191 <= p1_smul_76191_comb;
    p1_smul_76192 <= p1_smul_76192_comb;
    p1_smul_76193 <= p1_smul_76193_comb;
    p1_smul_76194 <= p1_smul_76194_comb;
    p1_smul_76195 <= p1_smul_76195_comb;
    p1_smul_76196 <= p1_smul_76196_comb;
    p1_smul_76197 <= p1_smul_76197_comb;
    p1_smul_76198 <= p1_smul_76198_comb;
    p1_smul_76199 <= p1_smul_76199_comb;
    p1_smul_76200 <= p1_smul_76200_comb;
    p1_smul_76201 <= p1_smul_76201_comb;
    p1_smul_76202 <= p1_smul_76202_comb;
    p1_smul_76203 <= p1_smul_76203_comb;
    p1_smul_76204 <= p1_smul_76204_comb;
    p1_smul_76205 <= p1_smul_76205_comb;
    p1_smul_76206 <= p1_smul_76206_comb;
    p1_smul_76207 <= p1_smul_76207_comb;
    p1_smul_76208 <= p1_smul_76208_comb;
    p1_smul_76209 <= p1_smul_76209_comb;
    p1_smul_76210 <= p1_smul_76210_comb;
    p1_smul_76211 <= p1_smul_76211_comb;
    p1_smul_76212 <= p1_smul_76212_comb;
    p1_smul_76213 <= p1_smul_76213_comb;
    p1_smul_76214 <= p1_smul_76214_comb;
    p1_smul_76215 <= p1_smul_76215_comb;
    p1_smul_76216 <= p1_smul_76216_comb;
    p1_smul_76217 <= p1_smul_76217_comb;
    p1_smul_76218 <= p1_smul_76218_comb;
    p1_smul_76219 <= p1_smul_76219_comb;
    p1_smul_76220 <= p1_smul_76220_comb;
    p1_smul_76221 <= p1_smul_76221_comb;
    p1_smul_76222 <= p1_smul_76222_comb;
    p1_smul_76223 <= p1_smul_76223_comb;
    p1_smul_76224 <= p1_smul_76224_comb;
    p1_smul_76225 <= p1_smul_76225_comb;
    p1_smul_76226 <= p1_smul_76226_comb;
    p1_smul_76227 <= p1_smul_76227_comb;
    p1_smul_76228 <= p1_smul_76228_comb;
    p1_smul_76229 <= p1_smul_76229_comb;
    p1_smul_76230 <= p1_smul_76230_comb;
    p1_smul_76231 <= p1_smul_76231_comb;
    p1_smul_76232 <= p1_smul_76232_comb;
    p1_smul_76233 <= p1_smul_76233_comb;
    p1_smul_76234 <= p1_smul_76234_comb;
    p1_smul_76235 <= p1_smul_76235_comb;
    p1_smul_76236 <= p1_smul_76236_comb;
    p1_smul_76237 <= p1_smul_76237_comb;
    p1_smul_76238 <= p1_smul_76238_comb;
    p1_smul_76239 <= p1_smul_76239_comb;
    p1_smul_76240 <= p1_smul_76240_comb;
    p1_smul_76241 <= p1_smul_76241_comb;
    p1_smul_76242 <= p1_smul_76242_comb;
    p1_smul_76243 <= p1_smul_76243_comb;
    p1_smul_76244 <= p1_smul_76244_comb;
    p1_smul_76245 <= p1_smul_76245_comb;
    p1_smul_76246 <= p1_smul_76246_comb;
    p1_smul_76247 <= p1_smul_76247_comb;
    p1_smul_76248 <= p1_smul_76248_comb;
    p1_smul_76249 <= p1_smul_76249_comb;
    p1_smul_76250 <= p1_smul_76250_comb;
    p1_smul_76251 <= p1_smul_76251_comb;
    p1_smul_76252 <= p1_smul_76252_comb;
    p1_smul_76253 <= p1_smul_76253_comb;
    p1_smul_76254 <= p1_smul_76254_comb;
    p1_smul_76255 <= p1_smul_76255_comb;
    p1_smul_76256 <= p1_smul_76256_comb;
    p1_smul_76257 <= p1_smul_76257_comb;
    p1_smul_76258 <= p1_smul_76258_comb;
    p1_smul_76259 <= p1_smul_76259_comb;
    p1_smul_76260 <= p1_smul_76260_comb;
    p1_smul_76261 <= p1_smul_76261_comb;
    p1_smul_76262 <= p1_smul_76262_comb;
    p1_smul_76263 <= p1_smul_76263_comb;
    p1_smul_76264 <= p1_smul_76264_comb;
    p1_smul_76265 <= p1_smul_76265_comb;
    p1_smul_76266 <= p1_smul_76266_comb;
    p1_smul_76267 <= p1_smul_76267_comb;
    p1_smul_76268 <= p1_smul_76268_comb;
    p1_smul_76269 <= p1_smul_76269_comb;
    p1_smul_76270 <= p1_smul_76270_comb;
    p1_smul_76271 <= p1_smul_76271_comb;
    p1_smul_76272 <= p1_smul_76272_comb;
    p1_smul_76273 <= p1_smul_76273_comb;
    p1_smul_76274 <= p1_smul_76274_comb;
    p1_smul_76275 <= p1_smul_76275_comb;
    p1_smul_76276 <= p1_smul_76276_comb;
    p1_smul_76277 <= p1_smul_76277_comb;
    p1_smul_76278 <= p1_smul_76278_comb;
    p1_smul_76279 <= p1_smul_76279_comb;
    p1_smul_76280 <= p1_smul_76280_comb;
    p1_smul_76281 <= p1_smul_76281_comb;
    p1_smul_76282 <= p1_smul_76282_comb;
    p1_smul_76283 <= p1_smul_76283_comb;
    p1_smul_76284 <= p1_smul_76284_comb;
    p1_smul_76285 <= p1_smul_76285_comb;
    p1_smul_76286 <= p1_smul_76286_comb;
    p1_smul_76287 <= p1_smul_76287_comb;
    p1_smul_76288 <= p1_smul_76288_comb;
    p1_smul_76289 <= p1_smul_76289_comb;
    p1_smul_76290 <= p1_smul_76290_comb;
    p1_smul_76291 <= p1_smul_76291_comb;
    p1_smul_76292 <= p1_smul_76292_comb;
    p1_smul_76293 <= p1_smul_76293_comb;
    p1_smul_76294 <= p1_smul_76294_comb;
    p1_smul_76295 <= p1_smul_76295_comb;
    p1_smul_76296 <= p1_smul_76296_comb;
    p1_smul_76297 <= p1_smul_76297_comb;
    p1_smul_76298 <= p1_smul_76298_comb;
    p1_smul_76299 <= p1_smul_76299_comb;
    p1_smul_76300 <= p1_smul_76300_comb;
    p1_smul_76301 <= p1_smul_76301_comb;
    p1_smul_76302 <= p1_smul_76302_comb;
    p1_smul_76303 <= p1_smul_76303_comb;
    p1_smul_76304 <= p1_smul_76304_comb;
    p1_smul_76305 <= p1_smul_76305_comb;
    p1_smul_76306 <= p1_smul_76306_comb;
    p1_smul_76307 <= p1_smul_76307_comb;
    p1_smul_76308 <= p1_smul_76308_comb;
    p1_smul_76309 <= p1_smul_76309_comb;
    p1_smul_76310 <= p1_smul_76310_comb;
    p1_smul_76311 <= p1_smul_76311_comb;
    p1_smul_76312 <= p1_smul_76312_comb;
    p1_smul_76313 <= p1_smul_76313_comb;
    p1_smul_76314 <= p1_smul_76314_comb;
    p1_smul_76315 <= p1_smul_76315_comb;
    p1_smul_76316 <= p1_smul_76316_comb;
    p1_smul_76317 <= p1_smul_76317_comb;
    p1_smul_76318 <= p1_smul_76318_comb;
    p1_smul_76319 <= p1_smul_76319_comb;
    p1_smul_76320 <= p1_smul_76320_comb;
    p1_smul_76321 <= p1_smul_76321_comb;
    p1_smul_76322 <= p1_smul_76322_comb;
    p1_smul_76323 <= p1_smul_76323_comb;
    p1_smul_76324 <= p1_smul_76324_comb;
    p1_smul_76325 <= p1_smul_76325_comb;
    p1_smul_76326 <= p1_smul_76326_comb;
    p1_smul_76327 <= p1_smul_76327_comb;
    p1_smul_76328 <= p1_smul_76328_comb;
    p1_smul_76329 <= p1_smul_76329_comb;
    p1_smul_76330 <= p1_smul_76330_comb;
    p1_smul_76331 <= p1_smul_76331_comb;
    p1_smul_76332 <= p1_smul_76332_comb;
    p1_smul_76333 <= p1_smul_76333_comb;
    p1_smul_76334 <= p1_smul_76334_comb;
    p1_smul_76335 <= p1_smul_76335_comb;
    p1_smul_76336 <= p1_smul_76336_comb;
    p1_smul_76337 <= p1_smul_76337_comb;
    p1_smul_76338 <= p1_smul_76338_comb;
    p1_smul_76339 <= p1_smul_76339_comb;
    p1_smul_76340 <= p1_smul_76340_comb;
    p1_smul_76341 <= p1_smul_76341_comb;
    p1_smul_76342 <= p1_smul_76342_comb;
    p1_smul_76343 <= p1_smul_76343_comb;
    p1_smul_76344 <= p1_smul_76344_comb;
    p1_smul_76345 <= p1_smul_76345_comb;
    p1_smul_76346 <= p1_smul_76346_comb;
    p1_smul_76347 <= p1_smul_76347_comb;
    p1_smul_76348 <= p1_smul_76348_comb;
    p1_smul_76349 <= p1_smul_76349_comb;
    p1_smul_76350 <= p1_smul_76350_comb;
    p1_smul_76351 <= p1_smul_76351_comb;
    p1_smul_76352 <= p1_smul_76352_comb;
    p1_smul_76353 <= p1_smul_76353_comb;
    p1_smul_76354 <= p1_smul_76354_comb;
    p1_smul_76355 <= p1_smul_76355_comb;
    p1_smul_76356 <= p1_smul_76356_comb;
    p1_smul_76357 <= p1_smul_76357_comb;
    p1_smul_76358 <= p1_smul_76358_comb;
    p1_smul_76359 <= p1_smul_76359_comb;
    p1_smul_76360 <= p1_smul_76360_comb;
    p1_smul_76361 <= p1_smul_76361_comb;
    p1_smul_76362 <= p1_smul_76362_comb;
    p1_smul_76363 <= p1_smul_76363_comb;
    p1_smul_76364 <= p1_smul_76364_comb;
    p1_smul_76365 <= p1_smul_76365_comb;
    p1_smul_76366 <= p1_smul_76366_comb;
    p1_smul_76367 <= p1_smul_76367_comb;
    p1_smul_76368 <= p1_smul_76368_comb;
    p1_smul_76369 <= p1_smul_76369_comb;
    p1_smul_76370 <= p1_smul_76370_comb;
    p1_smul_76371 <= p1_smul_76371_comb;
    p1_smul_76372 <= p1_smul_76372_comb;
    p1_smul_76373 <= p1_smul_76373_comb;
    p1_smul_76374 <= p1_smul_76374_comb;
    p1_smul_76375 <= p1_smul_76375_comb;
    p1_smul_76376 <= p1_smul_76376_comb;
    p1_smul_76377 <= p1_smul_76377_comb;
    p1_smul_76378 <= p1_smul_76378_comb;
    p1_smul_76379 <= p1_smul_76379_comb;
    p1_smul_76380 <= p1_smul_76380_comb;
    p1_smul_76381 <= p1_smul_76381_comb;
    p1_smul_76382 <= p1_smul_76382_comb;
    p1_smul_76383 <= p1_smul_76383_comb;
    p1_smul_76384 <= p1_smul_76384_comb;
    p1_smul_76385 <= p1_smul_76385_comb;
    p1_smul_76386 <= p1_smul_76386_comb;
    p1_smul_76387 <= p1_smul_76387_comb;
    p1_smul_76388 <= p1_smul_76388_comb;
    p1_smul_76389 <= p1_smul_76389_comb;
    p1_smul_76390 <= p1_smul_76390_comb;
    p1_smul_76391 <= p1_smul_76391_comb;
    p1_smul_76392 <= p1_smul_76392_comb;
    p1_smul_76393 <= p1_smul_76393_comb;
    p1_smul_76394 <= p1_smul_76394_comb;
    p1_smul_76395 <= p1_smul_76395_comb;
    p1_smul_76396 <= p1_smul_76396_comb;
    p1_smul_76397 <= p1_smul_76397_comb;
    p1_smul_76398 <= p1_smul_76398_comb;
    p1_smul_76399 <= p1_smul_76399_comb;
    p1_smul_76400 <= p1_smul_76400_comb;
    p1_smul_76401 <= p1_smul_76401_comb;
    p1_smul_76402 <= p1_smul_76402_comb;
    p1_smul_76403 <= p1_smul_76403_comb;
    p1_smul_76404 <= p1_smul_76404_comb;
    p1_smul_76405 <= p1_smul_76405_comb;
    p1_smul_76406 <= p1_smul_76406_comb;
    p1_smul_76407 <= p1_smul_76407_comb;
    p1_smul_76408 <= p1_smul_76408_comb;
    p1_smul_76409 <= p1_smul_76409_comb;
    p1_smul_76410 <= p1_smul_76410_comb;
    p1_smul_76411 <= p1_smul_76411_comb;
    p1_smul_76412 <= p1_smul_76412_comb;
    p1_smul_76413 <= p1_smul_76413_comb;
    p1_smul_76414 <= p1_smul_76414_comb;
    p1_smul_76415 <= p1_smul_76415_comb;
    p1_smul_76416 <= p1_smul_76416_comb;
    p1_smul_76417 <= p1_smul_76417_comb;
    p1_smul_76418 <= p1_smul_76418_comb;
    p1_smul_76419 <= p1_smul_76419_comb;
    p1_smul_76420 <= p1_smul_76420_comb;
    p1_smul_76421 <= p1_smul_76421_comb;
    p1_smul_76422 <= p1_smul_76422_comb;
    p1_smul_76423 <= p1_smul_76423_comb;
    p1_smul_76424 <= p1_smul_76424_comb;
    p1_smul_76425 <= p1_smul_76425_comb;
    p1_smul_76426 <= p1_smul_76426_comb;
    p1_smul_76427 <= p1_smul_76427_comb;
    p1_smul_76428 <= p1_smul_76428_comb;
    p1_smul_76429 <= p1_smul_76429_comb;
    p1_smul_76430 <= p1_smul_76430_comb;
    p1_smul_76431 <= p1_smul_76431_comb;
    p1_smul_76432 <= p1_smul_76432_comb;
    p1_smul_76433 <= p1_smul_76433_comb;
    p1_smul_76434 <= p1_smul_76434_comb;
    p1_smul_76435 <= p1_smul_76435_comb;
    p1_smul_76436 <= p1_smul_76436_comb;
    p1_smul_76437 <= p1_smul_76437_comb;
    p1_smul_76438 <= p1_smul_76438_comb;
    p1_smul_76439 <= p1_smul_76439_comb;
    p1_smul_76440 <= p1_smul_76440_comb;
    p1_smul_76441 <= p1_smul_76441_comb;
    p1_smul_76442 <= p1_smul_76442_comb;
    p1_smul_76443 <= p1_smul_76443_comb;
    p1_smul_76444 <= p1_smul_76444_comb;
    p1_smul_76445 <= p1_smul_76445_comb;
    p1_smul_76446 <= p1_smul_76446_comb;
    p1_smul_76447 <= p1_smul_76447_comb;
    p1_smul_76448 <= p1_smul_76448_comb;
    p1_smul_76449 <= p1_smul_76449_comb;
    p1_smul_76450 <= p1_smul_76450_comb;
    p1_smul_76451 <= p1_smul_76451_comb;
    p1_smul_76452 <= p1_smul_76452_comb;
    p1_smul_76453 <= p1_smul_76453_comb;
    p1_smul_76454 <= p1_smul_76454_comb;
    p1_smul_76455 <= p1_smul_76455_comb;
    p1_smul_76456 <= p1_smul_76456_comb;
    p1_smul_76457 <= p1_smul_76457_comb;
    p1_smul_76458 <= p1_smul_76458_comb;
    p1_smul_76459 <= p1_smul_76459_comb;
    p1_smul_76460 <= p1_smul_76460_comb;
    p1_smul_76461 <= p1_smul_76461_comb;
    p1_smul_76462 <= p1_smul_76462_comb;
    p1_smul_76463 <= p1_smul_76463_comb;
    p1_smul_76464 <= p1_smul_76464_comb;
    p1_smul_76465 <= p1_smul_76465_comb;
    p1_smul_76466 <= p1_smul_76466_comb;
    p1_smul_76467 <= p1_smul_76467_comb;
    p1_smul_76468 <= p1_smul_76468_comb;
    p1_smul_76469 <= p1_smul_76469_comb;
    p1_smul_76470 <= p1_smul_76470_comb;
    p1_smul_76471 <= p1_smul_76471_comb;
    p1_smul_76472 <= p1_smul_76472_comb;
    p1_smul_76473 <= p1_smul_76473_comb;
    p1_smul_76474 <= p1_smul_76474_comb;
    p1_smul_76475 <= p1_smul_76475_comb;
    p1_smul_76476 <= p1_smul_76476_comb;
    p1_smul_76477 <= p1_smul_76477_comb;
    p1_smul_76478 <= p1_smul_76478_comb;
    p1_smul_76479 <= p1_smul_76479_comb;
    p1_smul_76480 <= p1_smul_76480_comb;
    p1_smul_76481 <= p1_smul_76481_comb;
    p1_smul_76482 <= p1_smul_76482_comb;
    p1_smul_76483 <= p1_smul_76483_comb;
    p1_smul_76484 <= p1_smul_76484_comb;
    p1_smul_76485 <= p1_smul_76485_comb;
    p1_smul_76486 <= p1_smul_76486_comb;
    p1_smul_76487 <= p1_smul_76487_comb;
    p1_smul_76488 <= p1_smul_76488_comb;
    p1_smul_76489 <= p1_smul_76489_comb;
    p1_smul_76490 <= p1_smul_76490_comb;
    p1_smul_76491 <= p1_smul_76491_comb;
    p1_smul_76492 <= p1_smul_76492_comb;
    p1_smul_76493 <= p1_smul_76493_comb;
    p1_smul_76494 <= p1_smul_76494_comb;
    p1_smul_76495 <= p1_smul_76495_comb;
    p1_smul_76496 <= p1_smul_76496_comb;
    p1_smul_76497 <= p1_smul_76497_comb;
    p1_smul_76498 <= p1_smul_76498_comb;
    p1_smul_76499 <= p1_smul_76499_comb;
    p1_smul_76500 <= p1_smul_76500_comb;
    p1_smul_76501 <= p1_smul_76501_comb;
    p1_smul_76502 <= p1_smul_76502_comb;
    p1_smul_76503 <= p1_smul_76503_comb;
    p1_smul_76504 <= p1_smul_76504_comb;
    p1_smul_76505 <= p1_smul_76505_comb;
    p1_smul_76506 <= p1_smul_76506_comb;
    p1_smul_76507 <= p1_smul_76507_comb;
    p1_smul_76508 <= p1_smul_76508_comb;
    p1_smul_76509 <= p1_smul_76509_comb;
    p1_smul_76510 <= p1_smul_76510_comb;
    p1_smul_76511 <= p1_smul_76511_comb;
    p1_smul_76512 <= p1_smul_76512_comb;
    p1_smul_76513 <= p1_smul_76513_comb;
    p1_smul_76514 <= p1_smul_76514_comb;
    p1_smul_76515 <= p1_smul_76515_comb;
    p1_smul_76516 <= p1_smul_76516_comb;
    p1_smul_76517 <= p1_smul_76517_comb;
    p1_smul_76518 <= p1_smul_76518_comb;
    p1_smul_76519 <= p1_smul_76519_comb;
    p1_smul_76520 <= p1_smul_76520_comb;
    p1_smul_76521 <= p1_smul_76521_comb;
    p1_smul_76522 <= p1_smul_76522_comb;
    p1_smul_76523 <= p1_smul_76523_comb;
    p1_smul_76524 <= p1_smul_76524_comb;
    p1_smul_76525 <= p1_smul_76525_comb;
    p1_smul_76526 <= p1_smul_76526_comb;
    p1_smul_76527 <= p1_smul_76527_comb;
    p1_smul_76528 <= p1_smul_76528_comb;
    p1_smul_76529 <= p1_smul_76529_comb;
    p1_smul_76530 <= p1_smul_76530_comb;
    p1_smul_76531 <= p1_smul_76531_comb;
    p1_smul_76532 <= p1_smul_76532_comb;
    p1_smul_76533 <= p1_smul_76533_comb;
    p1_smul_76534 <= p1_smul_76534_comb;
    p1_smul_76535 <= p1_smul_76535_comb;
    p1_smul_76536 <= p1_smul_76536_comb;
    p1_smul_76537 <= p1_smul_76537_comb;
    p1_smul_76538 <= p1_smul_76538_comb;
    p1_smul_76539 <= p1_smul_76539_comb;
    p1_smul_76540 <= p1_smul_76540_comb;
    p1_smul_76541 <= p1_smul_76541_comb;
    p1_smul_76542 <= p1_smul_76542_comb;
    p1_smul_76543 <= p1_smul_76543_comb;
    p1_smul_76544 <= p1_smul_76544_comb;
    p1_smul_76545 <= p1_smul_76545_comb;
    p1_smul_76546 <= p1_smul_76546_comb;
    p1_smul_76547 <= p1_smul_76547_comb;
    p1_smul_76548 <= p1_smul_76548_comb;
    p1_smul_76549 <= p1_smul_76549_comb;
    p1_smul_76550 <= p1_smul_76550_comb;
    p1_smul_76551 <= p1_smul_76551_comb;
    p1_smul_76552 <= p1_smul_76552_comb;
    p1_smul_76553 <= p1_smul_76553_comb;
    p1_smul_76554 <= p1_smul_76554_comb;
    p1_smul_76555 <= p1_smul_76555_comb;
    p1_smul_76556 <= p1_smul_76556_comb;
    p1_smul_76557 <= p1_smul_76557_comb;
    p1_smul_76558 <= p1_smul_76558_comb;
    p1_smul_76559 <= p1_smul_76559_comb;
    p1_smul_76560 <= p1_smul_76560_comb;
    p1_smul_76561 <= p1_smul_76561_comb;
    p1_smul_76562 <= p1_smul_76562_comb;
    p1_smul_76563 <= p1_smul_76563_comb;
    p1_smul_76564 <= p1_smul_76564_comb;
    p1_smul_76565 <= p1_smul_76565_comb;
    p1_smul_76566 <= p1_smul_76566_comb;
    p1_smul_76567 <= p1_smul_76567_comb;
    p1_smul_76568 <= p1_smul_76568_comb;
    p1_smul_76569 <= p1_smul_76569_comb;
    p1_smul_76570 <= p1_smul_76570_comb;
    p1_smul_76571 <= p1_smul_76571_comb;
    p1_smul_76572 <= p1_smul_76572_comb;
    p1_smul_76573 <= p1_smul_76573_comb;
    p1_smul_76574 <= p1_smul_76574_comb;
    p1_smul_76575 <= p1_smul_76575_comb;
    p1_smul_76576 <= p1_smul_76576_comb;
    p1_smul_76577 <= p1_smul_76577_comb;
    p1_smul_76578 <= p1_smul_76578_comb;
    p1_smul_76579 <= p1_smul_76579_comb;
    p1_smul_76580 <= p1_smul_76580_comb;
    p1_smul_76581 <= p1_smul_76581_comb;
    p1_smul_76582 <= p1_smul_76582_comb;
    p1_smul_76583 <= p1_smul_76583_comb;
    p1_smul_76584 <= p1_smul_76584_comb;
    p1_smul_76585 <= p1_smul_76585_comb;
    p1_smul_76586 <= p1_smul_76586_comb;
    p1_smul_76587 <= p1_smul_76587_comb;
    p1_smul_76588 <= p1_smul_76588_comb;
    p1_smul_76589 <= p1_smul_76589_comb;
    p1_smul_76590 <= p1_smul_76590_comb;
    p1_smul_76591 <= p1_smul_76591_comb;
    p1_smul_76592 <= p1_smul_76592_comb;
    p1_smul_76593 <= p1_smul_76593_comb;
    p1_smul_76594 <= p1_smul_76594_comb;
    p1_smul_76595 <= p1_smul_76595_comb;
    p1_smul_76596 <= p1_smul_76596_comb;
    p1_smul_76597 <= p1_smul_76597_comb;
    p1_smul_76598 <= p1_smul_76598_comb;
    p1_smul_76599 <= p1_smul_76599_comb;
    p1_smul_76600 <= p1_smul_76600_comb;
    p1_smul_76601 <= p1_smul_76601_comb;
    p1_smul_76602 <= p1_smul_76602_comb;
    p1_smul_76603 <= p1_smul_76603_comb;
    p1_smul_76604 <= p1_smul_76604_comb;
    p1_smul_76605 <= p1_smul_76605_comb;
    p1_smul_76606 <= p1_smul_76606_comb;
    p1_smul_76607 <= p1_smul_76607_comb;
    p1_smul_76608 <= p1_smul_76608_comb;
    p1_smul_76609 <= p1_smul_76609_comb;
    p1_smul_76610 <= p1_smul_76610_comb;
    p1_smul_76611 <= p1_smul_76611_comb;
    p1_smul_76612 <= p1_smul_76612_comb;
    p1_smul_76613 <= p1_smul_76613_comb;
    p1_smul_76614 <= p1_smul_76614_comb;
    p1_smul_76615 <= p1_smul_76615_comb;
    p1_smul_76616 <= p1_smul_76616_comb;
    p1_smul_76617 <= p1_smul_76617_comb;
    p1_smul_76618 <= p1_smul_76618_comb;
    p1_smul_76619 <= p1_smul_76619_comb;
    p1_smul_76620 <= p1_smul_76620_comb;
    p1_smul_76621 <= p1_smul_76621_comb;
    p1_smul_76622 <= p1_smul_76622_comb;
    p1_smul_76623 <= p1_smul_76623_comb;
    p1_smul_76624 <= p1_smul_76624_comb;
    p1_smul_76625 <= p1_smul_76625_comb;
    p1_smul_76626 <= p1_smul_76626_comb;
    p1_smul_76627 <= p1_smul_76627_comb;
    p1_smul_76628 <= p1_smul_76628_comb;
    p1_smul_76629 <= p1_smul_76629_comb;
    p1_smul_76630 <= p1_smul_76630_comb;
    p1_smul_76631 <= p1_smul_76631_comb;
    p1_smul_76632 <= p1_smul_76632_comb;
    p1_smul_76633 <= p1_smul_76633_comb;
    p1_smul_76634 <= p1_smul_76634_comb;
    p1_smul_76635 <= p1_smul_76635_comb;
    p1_smul_76636 <= p1_smul_76636_comb;
    p1_smul_76637 <= p1_smul_76637_comb;
    p1_smul_76638 <= p1_smul_76638_comb;
    p1_smul_76639 <= p1_smul_76639_comb;
    p1_smul_76640 <= p1_smul_76640_comb;
    p1_smul_76641 <= p1_smul_76641_comb;
    p1_smul_76642 <= p1_smul_76642_comb;
    p1_smul_76643 <= p1_smul_76643_comb;
    p1_smul_76644 <= p1_smul_76644_comb;
    p1_smul_76645 <= p1_smul_76645_comb;
    p1_smul_76646 <= p1_smul_76646_comb;
    p1_smul_76647 <= p1_smul_76647_comb;
    p1_smul_76648 <= p1_smul_76648_comb;
    p1_smul_76649 <= p1_smul_76649_comb;
    p1_smul_76650 <= p1_smul_76650_comb;
    p1_smul_76651 <= p1_smul_76651_comb;
    p1_smul_76652 <= p1_smul_76652_comb;
    p1_smul_76653 <= p1_smul_76653_comb;
    p1_smul_76654 <= p1_smul_76654_comb;
    p1_smul_76655 <= p1_smul_76655_comb;
    p1_smul_76656 <= p1_smul_76656_comb;
    p1_smul_76657 <= p1_smul_76657_comb;
    p1_smul_76658 <= p1_smul_76658_comb;
    p1_smul_76659 <= p1_smul_76659_comb;
    p1_smul_76660 <= p1_smul_76660_comb;
    p1_smul_76661 <= p1_smul_76661_comb;
    p1_smul_76662 <= p1_smul_76662_comb;
    p1_smul_76663 <= p1_smul_76663_comb;
    p1_smul_76664 <= p1_smul_76664_comb;
    p1_smul_76665 <= p1_smul_76665_comb;
    p1_smul_76666 <= p1_smul_76666_comb;
    p1_smul_76667 <= p1_smul_76667_comb;
    p1_smul_76668 <= p1_smul_76668_comb;
    p1_smul_76669 <= p1_smul_76669_comb;
    p1_smul_76670 <= p1_smul_76670_comb;
    p1_smul_76671 <= p1_smul_76671_comb;
    p1_smul_76672 <= p1_smul_76672_comb;
    p1_smul_76673 <= p1_smul_76673_comb;
    p1_smul_76674 <= p1_smul_76674_comb;
    p1_smul_76675 <= p1_smul_76675_comb;
    p1_smul_76676 <= p1_smul_76676_comb;
    p1_smul_76677 <= p1_smul_76677_comb;
    p1_smul_76678 <= p1_smul_76678_comb;
    p1_smul_76679 <= p1_smul_76679_comb;
    p1_smul_76680 <= p1_smul_76680_comb;
    p1_smul_76681 <= p1_smul_76681_comb;
    p1_smul_76682 <= p1_smul_76682_comb;
    p1_smul_76683 <= p1_smul_76683_comb;
    p1_smul_76684 <= p1_smul_76684_comb;
    p1_smul_76685 <= p1_smul_76685_comb;
    p1_smul_76686 <= p1_smul_76686_comb;
    p1_smul_76687 <= p1_smul_76687_comb;
    p1_smul_76688 <= p1_smul_76688_comb;
    p1_smul_76689 <= p1_smul_76689_comb;
    p1_smul_76690 <= p1_smul_76690_comb;
    p1_smul_76691 <= p1_smul_76691_comb;
    p1_smul_76692 <= p1_smul_76692_comb;
    p1_smul_76693 <= p1_smul_76693_comb;
    p1_smul_76694 <= p1_smul_76694_comb;
    p1_smul_76695 <= p1_smul_76695_comb;
    p1_smul_76696 <= p1_smul_76696_comb;
    p1_smul_76697 <= p1_smul_76697_comb;
    p1_smul_76698 <= p1_smul_76698_comb;
    p1_smul_76699 <= p1_smul_76699_comb;
    p1_smul_76700 <= p1_smul_76700_comb;
    p1_smul_76701 <= p1_smul_76701_comb;
    p1_smul_76702 <= p1_smul_76702_comb;
    p1_smul_76703 <= p1_smul_76703_comb;
    p1_smul_76704 <= p1_smul_76704_comb;
    p1_smul_76705 <= p1_smul_76705_comb;
    p1_smul_76706 <= p1_smul_76706_comb;
    p1_smul_76707 <= p1_smul_76707_comb;
    p1_smul_76708 <= p1_smul_76708_comb;
    p1_smul_76709 <= p1_smul_76709_comb;
    p1_smul_76710 <= p1_smul_76710_comb;
    p1_smul_76711 <= p1_smul_76711_comb;
    p1_smul_76712 <= p1_smul_76712_comb;
    p1_smul_76713 <= p1_smul_76713_comb;
    p1_smul_76714 <= p1_smul_76714_comb;
    p1_smul_76715 <= p1_smul_76715_comb;
    p1_smul_76716 <= p1_smul_76716_comb;
    p1_smul_76717 <= p1_smul_76717_comb;
    p1_smul_76718 <= p1_smul_76718_comb;
    p1_smul_76719 <= p1_smul_76719_comb;
    p1_smul_76720 <= p1_smul_76720_comb;
    p1_smul_76721 <= p1_smul_76721_comb;
    p1_smul_76722 <= p1_smul_76722_comb;
    p1_smul_76723 <= p1_smul_76723_comb;
    p1_smul_76724 <= p1_smul_76724_comb;
    p1_smul_76725 <= p1_smul_76725_comb;
    p1_smul_76726 <= p1_smul_76726_comb;
    p1_smul_76727 <= p1_smul_76727_comb;
    p1_smul_76728 <= p1_smul_76728_comb;
    p1_smul_76729 <= p1_smul_76729_comb;
    p1_smul_76730 <= p1_smul_76730_comb;
    p1_smul_76731 <= p1_smul_76731_comb;
    p1_smul_76732 <= p1_smul_76732_comb;
    p1_smul_76733 <= p1_smul_76733_comb;
    p1_smul_76734 <= p1_smul_76734_comb;
    p1_smul_76735 <= p1_smul_76735_comb;
    p1_smul_76736 <= p1_smul_76736_comb;
    p1_smul_76737 <= p1_smul_76737_comb;
    p1_smul_76738 <= p1_smul_76738_comb;
    p1_smul_76739 <= p1_smul_76739_comb;
    p1_smul_76740 <= p1_smul_76740_comb;
    p1_smul_76741 <= p1_smul_76741_comb;
    p1_smul_76742 <= p1_smul_76742_comb;
    p1_smul_76743 <= p1_smul_76743_comb;
    p1_smul_76744 <= p1_smul_76744_comb;
    p1_smul_76745 <= p1_smul_76745_comb;
    p1_smul_76746 <= p1_smul_76746_comb;
    p1_smul_76747 <= p1_smul_76747_comb;
    p1_smul_76748 <= p1_smul_76748_comb;
    p1_smul_76749 <= p1_smul_76749_comb;
    p1_smul_76750 <= p1_smul_76750_comb;
    p1_smul_76751 <= p1_smul_76751_comb;
    p1_smul_76752 <= p1_smul_76752_comb;
    p1_smul_76753 <= p1_smul_76753_comb;
    p1_smul_76754 <= p1_smul_76754_comb;
    p1_smul_76755 <= p1_smul_76755_comb;
    p1_smul_76756 <= p1_smul_76756_comb;
    p1_smul_76757 <= p1_smul_76757_comb;
    p1_smul_76758 <= p1_smul_76758_comb;
    p1_smul_76759 <= p1_smul_76759_comb;
    p1_smul_76760 <= p1_smul_76760_comb;
    p1_smul_76761 <= p1_smul_76761_comb;
    p1_smul_76762 <= p1_smul_76762_comb;
    p1_smul_76763 <= p1_smul_76763_comb;
    p1_smul_76764 <= p1_smul_76764_comb;
    p1_smul_76765 <= p1_smul_76765_comb;
    p1_smul_76766 <= p1_smul_76766_comb;
    p1_smul_76767 <= p1_smul_76767_comb;
    p1_smul_76768 <= p1_smul_76768_comb;
    p1_smul_76769 <= p1_smul_76769_comb;
    p1_smul_76770 <= p1_smul_76770_comb;
    p1_smul_76771 <= p1_smul_76771_comb;
    p1_smul_76772 <= p1_smul_76772_comb;
    p1_smul_76773 <= p1_smul_76773_comb;
    p1_smul_76774 <= p1_smul_76774_comb;
    p1_smul_76775 <= p1_smul_76775_comb;
    p1_smul_76776 <= p1_smul_76776_comb;
    p1_smul_76777 <= p1_smul_76777_comb;
    p1_smul_76778 <= p1_smul_76778_comb;
    p1_smul_76779 <= p1_smul_76779_comb;
    p1_smul_76780 <= p1_smul_76780_comb;
    p1_smul_76781 <= p1_smul_76781_comb;
    p1_smul_76782 <= p1_smul_76782_comb;
    p1_smul_76783 <= p1_smul_76783_comb;
    p1_smul_76784 <= p1_smul_76784_comb;
    p1_smul_76785 <= p1_smul_76785_comb;
    p1_smul_76786 <= p1_smul_76786_comb;
    p1_smul_76787 <= p1_smul_76787_comb;
    p1_smul_76788 <= p1_smul_76788_comb;
    p1_smul_76789 <= p1_smul_76789_comb;
    p1_smul_76790 <= p1_smul_76790_comb;
    p1_smul_76791 <= p1_smul_76791_comb;
    p1_smul_76792 <= p1_smul_76792_comb;
    p1_smul_76793 <= p1_smul_76793_comb;
    p1_smul_76794 <= p1_smul_76794_comb;
    p1_smul_76795 <= p1_smul_76795_comb;
    p1_smul_76796 <= p1_smul_76796_comb;
    p1_smul_76797 <= p1_smul_76797_comb;
    p1_smul_76798 <= p1_smul_76798_comb;
    p1_smul_76799 <= p1_smul_76799_comb;
    p1_smul_76800 <= p1_smul_76800_comb;
    p1_smul_76801 <= p1_smul_76801_comb;
    p1_smul_76802 <= p1_smul_76802_comb;
    p1_smul_76803 <= p1_smul_76803_comb;
    p1_smul_76804 <= p1_smul_76804_comb;
    p1_smul_76805 <= p1_smul_76805_comb;
    p1_smul_76806 <= p1_smul_76806_comb;
    p1_smul_76807 <= p1_smul_76807_comb;
    p1_smul_76808 <= p1_smul_76808_comb;
    p1_smul_76809 <= p1_smul_76809_comb;
    p1_smul_76810 <= p1_smul_76810_comb;
    p1_smul_76811 <= p1_smul_76811_comb;
    p1_smul_76812 <= p1_smul_76812_comb;
    p1_smul_76813 <= p1_smul_76813_comb;
    p1_smul_76814 <= p1_smul_76814_comb;
    p1_smul_76815 <= p1_smul_76815_comb;
    p1_smul_76816 <= p1_smul_76816_comb;
    p1_smul_76817 <= p1_smul_76817_comb;
    p1_smul_76818 <= p1_smul_76818_comb;
    p1_smul_76819 <= p1_smul_76819_comb;
    p1_smul_76820 <= p1_smul_76820_comb;
    p1_smul_76821 <= p1_smul_76821_comb;
    p1_smul_76822 <= p1_smul_76822_comb;
    p1_smul_76823 <= p1_smul_76823_comb;
    p1_smul_76824 <= p1_smul_76824_comb;
    p1_smul_76825 <= p1_smul_76825_comb;
    p1_smul_76826 <= p1_smul_76826_comb;
    p1_smul_76827 <= p1_smul_76827_comb;
    p1_smul_76828 <= p1_smul_76828_comb;
    p1_smul_76829 <= p1_smul_76829_comb;
    p1_smul_76830 <= p1_smul_76830_comb;
    p1_smul_76831 <= p1_smul_76831_comb;
    p1_smul_76832 <= p1_smul_76832_comb;
    p1_smul_76833 <= p1_smul_76833_comb;
    p1_smul_76834 <= p1_smul_76834_comb;
    p1_smul_76835 <= p1_smul_76835_comb;
    p1_smul_76836 <= p1_smul_76836_comb;
    p1_smul_76837 <= p1_smul_76837_comb;
    p1_smul_76838 <= p1_smul_76838_comb;
    p1_smul_76839 <= p1_smul_76839_comb;
    p1_smul_76840 <= p1_smul_76840_comb;
    p1_smul_76841 <= p1_smul_76841_comb;
    p1_smul_76842 <= p1_smul_76842_comb;
    p1_smul_76843 <= p1_smul_76843_comb;
    p1_smul_76844 <= p1_smul_76844_comb;
    p1_smul_76845 <= p1_smul_76845_comb;
    p1_smul_76846 <= p1_smul_76846_comb;
    p1_smul_76847 <= p1_smul_76847_comb;
    p1_smul_76848 <= p1_smul_76848_comb;
    p1_smul_76849 <= p1_smul_76849_comb;
    p1_smul_76850 <= p1_smul_76850_comb;
    p1_smul_76851 <= p1_smul_76851_comb;
    p1_smul_76852 <= p1_smul_76852_comb;
    p1_smul_76853 <= p1_smul_76853_comb;
    p1_smul_76854 <= p1_smul_76854_comb;
    p1_smul_76855 <= p1_smul_76855_comb;
    p1_smul_76856 <= p1_smul_76856_comb;
    p1_smul_76857 <= p1_smul_76857_comb;
    p1_smul_76858 <= p1_smul_76858_comb;
    p1_smul_76859 <= p1_smul_76859_comb;
    p1_smul_76860 <= p1_smul_76860_comb;
    p1_smul_76861 <= p1_smul_76861_comb;
    p1_smul_76862 <= p1_smul_76862_comb;
    p1_smul_76863 <= p1_smul_76863_comb;
    p1_smul_76864 <= p1_smul_76864_comb;
    p1_smul_76865 <= p1_smul_76865_comb;
    p1_smul_76866 <= p1_smul_76866_comb;
    p1_smul_76867 <= p1_smul_76867_comb;
    p1_smul_76868 <= p1_smul_76868_comb;
    p1_smul_76869 <= p1_smul_76869_comb;
    p1_smul_76870 <= p1_smul_76870_comb;
    p1_smul_76871 <= p1_smul_76871_comb;
    p1_smul_76872 <= p1_smul_76872_comb;
    p1_smul_76873 <= p1_smul_76873_comb;
    p1_smul_76874 <= p1_smul_76874_comb;
    p1_smul_76875 <= p1_smul_76875_comb;
    p1_smul_76876 <= p1_smul_76876_comb;
    p1_smul_76877 <= p1_smul_76877_comb;
    p1_smul_76878 <= p1_smul_76878_comb;
    p1_smul_76879 <= p1_smul_76879_comb;
    p1_smul_76880 <= p1_smul_76880_comb;
    p1_smul_76881 <= p1_smul_76881_comb;
    p1_smul_76882 <= p1_smul_76882_comb;
    p1_smul_76883 <= p1_smul_76883_comb;
    p1_smul_76884 <= p1_smul_76884_comb;
    p1_smul_76885 <= p1_smul_76885_comb;
    p1_smul_76886 <= p1_smul_76886_comb;
    p1_smul_76887 <= p1_smul_76887_comb;
    p1_smul_76888 <= p1_smul_76888_comb;
    p1_smul_76889 <= p1_smul_76889_comb;
    p1_smul_76890 <= p1_smul_76890_comb;
    p1_smul_76891 <= p1_smul_76891_comb;
    p1_smul_76892 <= p1_smul_76892_comb;
    p1_smul_76893 <= p1_smul_76893_comb;
    p1_smul_76894 <= p1_smul_76894_comb;
    p1_smul_76895 <= p1_smul_76895_comb;
    p1_smul_76896 <= p1_smul_76896_comb;
    p1_smul_76897 <= p1_smul_76897_comb;
    p1_smul_76898 <= p1_smul_76898_comb;
    p1_smul_76899 <= p1_smul_76899_comb;
    p1_smul_76900 <= p1_smul_76900_comb;
    p1_smul_76901 <= p1_smul_76901_comb;
    p1_smul_76902 <= p1_smul_76902_comb;
    p1_smul_76903 <= p1_smul_76903_comb;
    p1_smul_76904 <= p1_smul_76904_comb;
    p1_smul_76905 <= p1_smul_76905_comb;
    p1_smul_76906 <= p1_smul_76906_comb;
    p1_smul_76907 <= p1_smul_76907_comb;
    p1_smul_76908 <= p1_smul_76908_comb;
    p1_smul_76909 <= p1_smul_76909_comb;
    p1_smul_76910 <= p1_smul_76910_comb;
    p1_smul_76911 <= p1_smul_76911_comb;
    p1_smul_76912 <= p1_smul_76912_comb;
    p1_smul_76913 <= p1_smul_76913_comb;
    p1_smul_76914 <= p1_smul_76914_comb;
    p1_smul_76915 <= p1_smul_76915_comb;
    p1_smul_76916 <= p1_smul_76916_comb;
    p1_smul_76917 <= p1_smul_76917_comb;
    p1_smul_76918 <= p1_smul_76918_comb;
    p1_smul_76919 <= p1_smul_76919_comb;
    p1_smul_76920 <= p1_smul_76920_comb;
    p1_smul_76921 <= p1_smul_76921_comb;
    p1_smul_76922 <= p1_smul_76922_comb;
    p1_smul_76923 <= p1_smul_76923_comb;
    p1_smul_76924 <= p1_smul_76924_comb;
    p1_smul_76925 <= p1_smul_76925_comb;
    p1_smul_76926 <= p1_smul_76926_comb;
    p1_smul_76927 <= p1_smul_76927_comb;
    p1_smul_76928 <= p1_smul_76928_comb;
    p1_smul_76929 <= p1_smul_76929_comb;
    p1_smul_76930 <= p1_smul_76930_comb;
    p1_smul_76931 <= p1_smul_76931_comb;
    p1_smul_76932 <= p1_smul_76932_comb;
    p1_smul_76933 <= p1_smul_76933_comb;
    p1_smul_76934 <= p1_smul_76934_comb;
    p1_smul_76935 <= p1_smul_76935_comb;
    p1_smul_76936 <= p1_smul_76936_comb;
    p1_smul_76937 <= p1_smul_76937_comb;
    p1_smul_76938 <= p1_smul_76938_comb;
    p1_smul_76939 <= p1_smul_76939_comb;
    p1_smul_76940 <= p1_smul_76940_comb;
    p1_smul_76941 <= p1_smul_76941_comb;
    p1_smul_76942 <= p1_smul_76942_comb;
    p1_smul_76943 <= p1_smul_76943_comb;
    p1_smul_76944 <= p1_smul_76944_comb;
    p1_smul_76945 <= p1_smul_76945_comb;
    p1_smul_76946 <= p1_smul_76946_comb;
    p1_smul_76947 <= p1_smul_76947_comb;
    p1_smul_76948 <= p1_smul_76948_comb;
    p1_smul_76949 <= p1_smul_76949_comb;
    p1_smul_76950 <= p1_smul_76950_comb;
    p1_smul_76951 <= p1_smul_76951_comb;
    p1_smul_76952 <= p1_smul_76952_comb;
    p1_smul_76953 <= p1_smul_76953_comb;
    p1_smul_76954 <= p1_smul_76954_comb;
    p1_smul_76955 <= p1_smul_76955_comb;
    p1_smul_76956 <= p1_smul_76956_comb;
    p1_smul_76957 <= p1_smul_76957_comb;
    p1_smul_76958 <= p1_smul_76958_comb;
    p1_smul_76959 <= p1_smul_76959_comb;
    p1_smul_76960 <= p1_smul_76960_comb;
    p1_smul_76961 <= p1_smul_76961_comb;
    p1_smul_76962 <= p1_smul_76962_comb;
    p1_smul_76963 <= p1_smul_76963_comb;
    p1_smul_76964 <= p1_smul_76964_comb;
    p1_smul_76965 <= p1_smul_76965_comb;
    p1_smul_76966 <= p1_smul_76966_comb;
    p1_smul_76967 <= p1_smul_76967_comb;
    p1_smul_76968 <= p1_smul_76968_comb;
    p1_smul_76969 <= p1_smul_76969_comb;
    p1_smul_76970 <= p1_smul_76970_comb;
    p1_smul_76971 <= p1_smul_76971_comb;
  end

  // ===== Pipe stage 2:
  wire [31:0] p2_add_78986_comb;
  wire [31:0] p2_add_78987_comb;
  wire [31:0] p2_add_78988_comb;
  wire [31:0] p2_add_78989_comb;
  wire [31:0] p2_add_78990_comb;
  wire [31:0] p2_add_78991_comb;
  wire [31:0] p2_add_78992_comb;
  wire [31:0] p2_add_78993_comb;
  wire [31:0] p2_add_78994_comb;
  wire [31:0] p2_add_78995_comb;
  wire [31:0] p2_add_78996_comb;
  wire [31:0] p2_add_78997_comb;
  wire [31:0] p2_add_78998_comb;
  wire [31:0] p2_add_78999_comb;
  wire [31:0] p2_add_79000_comb;
  wire [31:0] p2_add_79001_comb;
  wire [31:0] p2_add_79002_comb;
  wire [31:0] p2_add_79003_comb;
  wire [31:0] p2_add_79004_comb;
  wire [31:0] p2_add_79005_comb;
  wire [31:0] p2_add_79006_comb;
  wire [31:0] p2_add_79007_comb;
  wire [31:0] p2_add_79008_comb;
  wire [31:0] p2_add_79009_comb;
  wire [31:0] p2_add_79010_comb;
  wire [31:0] p2_add_79011_comb;
  wire [31:0] p2_add_79012_comb;
  wire [31:0] p2_add_79013_comb;
  wire [31:0] p2_add_79014_comb;
  wire [31:0] p2_add_79015_comb;
  wire [31:0] p2_add_79016_comb;
  wire [31:0] p2_add_79017_comb;
  wire [31:0] p2_add_79018_comb;
  wire [31:0] p2_add_79019_comb;
  wire [31:0] p2_add_79020_comb;
  wire [31:0] p2_add_79021_comb;
  wire [31:0] p2_add_79022_comb;
  wire [31:0] p2_add_79023_comb;
  wire [31:0] p2_add_79024_comb;
  wire [31:0] p2_add_79025_comb;
  wire [31:0] p2_add_79026_comb;
  wire [31:0] p2_add_79027_comb;
  wire [31:0] p2_add_79028_comb;
  wire [31:0] p2_add_79029_comb;
  wire [31:0] p2_add_79030_comb;
  wire [31:0] p2_add_79031_comb;
  wire [31:0] p2_add_79032_comb;
  wire [31:0] p2_add_79033_comb;
  wire [31:0] p2_add_79034_comb;
  wire [31:0] p2_add_79035_comb;
  wire [31:0] p2_add_79036_comb;
  wire [31:0] p2_add_79037_comb;
  wire [31:0] p2_add_79038_comb;
  wire [31:0] p2_add_79039_comb;
  wire [31:0] p2_add_79040_comb;
  wire [31:0] p2_add_79041_comb;
  wire [31:0] p2_add_79042_comb;
  wire [31:0] p2_add_79043_comb;
  wire [31:0] p2_add_79044_comb;
  wire [31:0] p2_add_79045_comb;
  wire [31:0] p2_add_79046_comb;
  wire [31:0] p2_add_79047_comb;
  wire [31:0] p2_add_79048_comb;
  wire [31:0] p2_add_79049_comb;
  wire [31:0] p2_add_79050_comb;
  wire [31:0] p2_add_79051_comb;
  wire [31:0] p2_add_79052_comb;
  wire [31:0] p2_add_79053_comb;
  wire [31:0] p2_add_79054_comb;
  wire [31:0] p2_add_79055_comb;
  wire [31:0] p2_add_79056_comb;
  wire [31:0] p2_add_79057_comb;
  wire [31:0] p2_add_79058_comb;
  wire [31:0] p2_add_79059_comb;
  wire [31:0] p2_add_79060_comb;
  wire [31:0] p2_add_79061_comb;
  wire [31:0] p2_add_79062_comb;
  wire [31:0] p2_add_79063_comb;
  wire [31:0] p2_add_79064_comb;
  wire [31:0] p2_add_79065_comb;
  wire [31:0] p2_add_79066_comb;
  wire [31:0] p2_add_79067_comb;
  wire [31:0] p2_add_79068_comb;
  wire [31:0] p2_add_79069_comb;
  wire [31:0] p2_add_79070_comb;
  wire [31:0] p2_add_79071_comb;
  wire [31:0] p2_add_79072_comb;
  wire [31:0] p2_add_79073_comb;
  wire [31:0] p2_add_79074_comb;
  wire [31:0] p2_add_79075_comb;
  wire [31:0] p2_add_79076_comb;
  wire [31:0] p2_add_79077_comb;
  wire [31:0] p2_add_79078_comb;
  wire [31:0] p2_add_79079_comb;
  wire [31:0] p2_add_79080_comb;
  wire [31:0] p2_add_79081_comb;
  wire [31:0] p2_add_79082_comb;
  wire [31:0] p2_add_79083_comb;
  wire [31:0] p2_add_79084_comb;
  wire [31:0] p2_add_79085_comb;
  wire [31:0] p2_add_79086_comb;
  wire [31:0] p2_add_79087_comb;
  wire [31:0] p2_add_79088_comb;
  wire [31:0] p2_add_79089_comb;
  wire [31:0] p2_add_79090_comb;
  wire [31:0] p2_add_79091_comb;
  wire [31:0] p2_add_79092_comb;
  wire [31:0] p2_add_79093_comb;
  wire [31:0] p2_add_79094_comb;
  wire [31:0] p2_add_79095_comb;
  wire [31:0] p2_add_79096_comb;
  wire [31:0] p2_add_79097_comb;
  wire [31:0] p2_add_79098_comb;
  wire [31:0] p2_add_79099_comb;
  wire [31:0] p2_add_79100_comb;
  wire [31:0] p2_add_79101_comb;
  wire [31:0] p2_add_79102_comb;
  wire [31:0] p2_add_79103_comb;
  wire [31:0] p2_add_79104_comb;
  wire [31:0] p2_add_79105_comb;
  wire [31:0] p2_add_79106_comb;
  wire [31:0] p2_add_79107_comb;
  wire [31:0] p2_add_79108_comb;
  wire [31:0] p2_add_79109_comb;
  wire [31:0] p2_add_79110_comb;
  wire [31:0] p2_add_79111_comb;
  wire [31:0] p2_add_79112_comb;
  wire [31:0] p2_add_79113_comb;
  wire [31:0] p2_add_79114_comb;
  wire [31:0] p2_add_79115_comb;
  wire [31:0] p2_add_79116_comb;
  wire [31:0] p2_add_79117_comb;
  wire [31:0] p2_add_79118_comb;
  wire [31:0] p2_add_79119_comb;
  wire [31:0] p2_add_79120_comb;
  wire [31:0] p2_add_79121_comb;
  wire [31:0] p2_add_79122_comb;
  wire [31:0] p2_add_79123_comb;
  wire [31:0] p2_add_79124_comb;
  wire [31:0] p2_add_79125_comb;
  wire [31:0] p2_add_79126_comb;
  wire [31:0] p2_add_79127_comb;
  wire [31:0] p2_add_79128_comb;
  wire [31:0] p2_add_79129_comb;
  wire [31:0] p2_add_79130_comb;
  wire [31:0] p2_add_79131_comb;
  wire [31:0] p2_add_79132_comb;
  wire [31:0] p2_add_79133_comb;
  wire [31:0] p2_add_79134_comb;
  wire [31:0] p2_add_79135_comb;
  wire [31:0] p2_add_79136_comb;
  wire [31:0] p2_add_79137_comb;
  wire [31:0] p2_add_79138_comb;
  wire [31:0] p2_add_79139_comb;
  wire [31:0] p2_add_79140_comb;
  wire [31:0] p2_add_79141_comb;
  wire [31:0] p2_add_79142_comb;
  wire [31:0] p2_add_79143_comb;
  wire [31:0] p2_add_79144_comb;
  wire [31:0] p2_add_79145_comb;
  wire [31:0] p2_add_79146_comb;
  wire [31:0] p2_add_79147_comb;
  wire [31:0] p2_add_79148_comb;
  wire [31:0] p2_add_79149_comb;
  wire [31:0] p2_add_79150_comb;
  wire [31:0] p2_add_79151_comb;
  wire [31:0] p2_add_79152_comb;
  wire [31:0] p2_add_79153_comb;
  wire [31:0] p2_add_79154_comb;
  wire [31:0] p2_add_79155_comb;
  wire [31:0] p2_add_79156_comb;
  wire [31:0] p2_add_79157_comb;
  wire [31:0] p2_add_79158_comb;
  wire [31:0] p2_add_79159_comb;
  wire [31:0] p2_add_79160_comb;
  wire [31:0] p2_add_79161_comb;
  wire [31:0] p2_add_79162_comb;
  wire [31:0] p2_add_79163_comb;
  wire [31:0] p2_add_79164_comb;
  wire [31:0] p2_add_79165_comb;
  wire [31:0] p2_add_79166_comb;
  wire [31:0] p2_add_79167_comb;
  wire [31:0] p2_add_79168_comb;
  wire [31:0] p2_add_79169_comb;
  wire [31:0] p2_add_79170_comb;
  wire [31:0] p2_add_79171_comb;
  wire [31:0] p2_add_79172_comb;
  wire [31:0] p2_add_79173_comb;
  wire [31:0] p2_add_79174_comb;
  wire [31:0] p2_add_79175_comb;
  wire [31:0] p2_add_79176_comb;
  wire [31:0] p2_add_79177_comb;
  wire [31:0] p2_add_79178_comb;
  wire [31:0] p2_add_79179_comb;
  wire [31:0] p2_add_79180_comb;
  wire [31:0] p2_add_79181_comb;
  wire [31:0] p2_add_79182_comb;
  wire [31:0] p2_add_79183_comb;
  wire [31:0] p2_add_79184_comb;
  wire [31:0] p2_add_79185_comb;
  wire [31:0] p2_add_79188_comb;
  wire [31:0] p2_add_79189_comb;
  wire [31:0] p2_add_79192_comb;
  wire [31:0] p2_add_79193_comb;
  wire [31:0] p2_add_79196_comb;
  wire [31:0] p2_add_79197_comb;
  wire [31:0] p2_add_79200_comb;
  wire [31:0] p2_add_79201_comb;
  wire [31:0] p2_add_79204_comb;
  wire [31:0] p2_add_79205_comb;
  wire [31:0] p2_add_79208_comb;
  wire [31:0] p2_add_79209_comb;
  wire [31:0] p2_add_79212_comb;
  wire [31:0] p2_add_79213_comb;
  wire [31:0] p2_add_79216_comb;
  wire [31:0] p2_add_79217_comb;
  wire [31:0] p2_add_79220_comb;
  wire [31:0] p2_add_79221_comb;
  wire [31:0] p2_add_79224_comb;
  wire [31:0] p2_add_79225_comb;
  wire [31:0] p2_add_79228_comb;
  wire [31:0] p2_add_79229_comb;
  wire [31:0] p2_add_79232_comb;
  wire [31:0] p2_add_79233_comb;
  wire [31:0] p2_add_79236_comb;
  wire [31:0] p2_add_79237_comb;
  wire [31:0] p2_add_79240_comb;
  wire [31:0] p2_add_79241_comb;
  wire [31:0] p2_add_79244_comb;
  wire [31:0] p2_add_79245_comb;
  wire [31:0] p2_add_79248_comb;
  wire [31:0] p2_add_79249_comb;
  wire [31:0] p2_add_79252_comb;
  wire [31:0] p2_add_79253_comb;
  wire [31:0] p2_add_79256_comb;
  wire [31:0] p2_add_79257_comb;
  wire [31:0] p2_add_79260_comb;
  wire [31:0] p2_add_79261_comb;
  wire [31:0] p2_add_79264_comb;
  wire [31:0] p2_add_79265_comb;
  wire [31:0] p2_add_79268_comb;
  wire [31:0] p2_add_79269_comb;
  wire [31:0] p2_add_79272_comb;
  wire [31:0] p2_add_79273_comb;
  wire [31:0] p2_add_79276_comb;
  wire [31:0] p2_add_79277_comb;
  wire [31:0] p2_add_79280_comb;
  wire [31:0] p2_add_79281_comb;
  wire [31:0] p2_add_79284_comb;
  wire [31:0] p2_add_79285_comb;
  wire [31:0] p2_add_79288_comb;
  wire [31:0] p2_add_79289_comb;
  wire [31:0] p2_add_79292_comb;
  wire [31:0] p2_add_79293_comb;
  wire [31:0] p2_add_79296_comb;
  wire [31:0] p2_add_79297_comb;
  wire [31:0] p2_add_79300_comb;
  wire [31:0] p2_add_79301_comb;
  wire [31:0] p2_add_79304_comb;
  wire [31:0] p2_add_79305_comb;
  wire [31:0] p2_add_79308_comb;
  wire [31:0] p2_add_79309_comb;
  wire [31:0] p2_add_79312_comb;
  wire [31:0] p2_add_79313_comb;
  wire [31:0] p2_add_79316_comb;
  wire [31:0] p2_add_79317_comb;
  wire [31:0] p2_add_79320_comb;
  wire [31:0] p2_add_79321_comb;
  wire [31:0] p2_add_79324_comb;
  wire [31:0] p2_add_79325_comb;
  wire [31:0] p2_add_79328_comb;
  wire [31:0] p2_add_79329_comb;
  wire [31:0] p2_add_79332_comb;
  wire [31:0] p2_add_79333_comb;
  wire [31:0] p2_add_79336_comb;
  wire [31:0] p2_add_79337_comb;
  wire [31:0] p2_add_79340_comb;
  wire [31:0] p2_add_79341_comb;
  wire [31:0] p2_add_79344_comb;
  wire [31:0] p2_add_79345_comb;
  wire [31:0] p2_add_79348_comb;
  wire [31:0] p2_add_79349_comb;
  wire [31:0] p2_add_79352_comb;
  wire [31:0] p2_add_79353_comb;
  wire [31:0] p2_add_79356_comb;
  wire [31:0] p2_add_79357_comb;
  wire [31:0] p2_add_79360_comb;
  wire [31:0] p2_add_79361_comb;
  wire [31:0] p2_add_79364_comb;
  wire [31:0] p2_add_79365_comb;
  wire [31:0] p2_add_79368_comb;
  wire [31:0] p2_add_79369_comb;
  wire [31:0] p2_add_79372_comb;
  wire [31:0] p2_add_79373_comb;
  wire [31:0] p2_add_79376_comb;
  wire [31:0] p2_add_79377_comb;
  wire [31:0] p2_add_79380_comb;
  wire [31:0] p2_add_79381_comb;
  wire [31:0] p2_add_79384_comb;
  wire [31:0] p2_add_79385_comb;
  wire [31:0] p2_add_79388_comb;
  wire [31:0] p2_add_79389_comb;
  wire [31:0] p2_add_79392_comb;
  wire [31:0] p2_add_79393_comb;
  wire [31:0] p2_add_79396_comb;
  wire [31:0] p2_add_79397_comb;
  wire [31:0] p2_add_79400_comb;
  wire [31:0] p2_add_79401_comb;
  wire [31:0] p2_add_79404_comb;
  wire [31:0] p2_add_79405_comb;
  wire [31:0] p2_add_79408_comb;
  wire [31:0] p2_add_79409_comb;
  wire [31:0] p2_add_79412_comb;
  wire [31:0] p2_add_79413_comb;
  wire [31:0] p2_add_79416_comb;
  wire [31:0] p2_add_79417_comb;
  wire [31:0] p2_add_79420_comb;
  wire [31:0] p2_add_79421_comb;
  wire [31:0] p2_add_79424_comb;
  wire [31:0] p2_add_79425_comb;
  wire [31:0] p2_add_79428_comb;
  wire [31:0] p2_add_79429_comb;
  wire [31:0] p2_add_79432_comb;
  wire [31:0] p2_add_79433_comb;
  wire [31:0] p2_add_79436_comb;
  wire [31:0] p2_add_79437_comb;
  wire [31:0] p2_add_79440_comb;
  wire [31:0] p2_add_79441_comb;
  wire [31:0] p2_add_79444_comb;
  wire [31:0] p2_add_79445_comb;
  wire [31:0] p2_add_79448_comb;
  wire [31:0] p2_add_79449_comb;
  wire [31:0] p2_add_79452_comb;
  wire [31:0] p2_add_79453_comb;
  wire [31:0] p2_add_79456_comb;
  wire [31:0] p2_add_79457_comb;
  wire [31:0] p2_add_79460_comb;
  wire [31:0] p2_add_79461_comb;
  wire [31:0] p2_add_79464_comb;
  wire [31:0] p2_add_79465_comb;
  wire [31:0] p2_add_79468_comb;
  wire [31:0] p2_add_79469_comb;
  wire [31:0] p2_add_79472_comb;
  wire [31:0] p2_add_79473_comb;
  wire [31:0] p2_add_79476_comb;
  wire [31:0] p2_add_79477_comb;
  wire [31:0] p2_add_79480_comb;
  wire [31:0] p2_add_79481_comb;
  wire [31:0] p2_add_79484_comb;
  wire [31:0] p2_add_79485_comb;
  wire [31:0] p2_add_79488_comb;
  wire [31:0] p2_add_79489_comb;
  wire [31:0] p2_add_79492_comb;
  wire [31:0] p2_add_79493_comb;
  wire [31:0] p2_add_79496_comb;
  wire [31:0] p2_add_79497_comb;
  wire [31:0] p2_add_79500_comb;
  wire [31:0] p2_add_79501_comb;
  wire [31:0] p2_add_79504_comb;
  wire [31:0] p2_add_79505_comb;
  wire [31:0] p2_add_79508_comb;
  wire [31:0] p2_add_79509_comb;
  wire [31:0] p2_add_79512_comb;
  wire [31:0] p2_add_79513_comb;
  wire [31:0] p2_add_79516_comb;
  wire [31:0] p2_add_79517_comb;
  wire [31:0] p2_add_79520_comb;
  wire [31:0] p2_add_79521_comb;
  wire [31:0] p2_add_79524_comb;
  wire [31:0] p2_add_79525_comb;
  wire [31:0] p2_add_79528_comb;
  wire [31:0] p2_add_79529_comb;
  wire [31:0] p2_add_79532_comb;
  wire [31:0] p2_add_79533_comb;
  wire [31:0] p2_add_79536_comb;
  wire [31:0] p2_add_79537_comb;
  wire [31:0] p2_add_79540_comb;
  wire [31:0] p2_add_79541_comb;
  wire [31:0] p2_add_79544_comb;
  wire [31:0] p2_add_79545_comb;
  wire [31:0] p2_add_79548_comb;
  wire [31:0] p2_add_79549_comb;
  wire [31:0] p2_add_79552_comb;
  wire [31:0] p2_add_79553_comb;
  wire [31:0] p2_add_79556_comb;
  wire [31:0] p2_add_79557_comb;
  wire [31:0] p2_add_79560_comb;
  wire [31:0] p2_add_79561_comb;
  wire [31:0] p2_add_79564_comb;
  wire [31:0] p2_add_79565_comb;
  wire [31:0] p2_add_79568_comb;
  wire [31:0] p2_add_79569_comb;
  wire [31:0] p2_add_79572_comb;
  wire [31:0] p2_add_79573_comb;
  wire [31:0] p2_add_79576_comb;
  wire [31:0] p2_add_79577_comb;
  wire [31:0] p2_add_79580_comb;
  wire [31:0] p2_add_79581_comb;
  wire [31:0] p2_add_79584_comb;
  wire [31:0] p2_add_79585_comb;
  wire [31:0] p2_add_79186_comb;
  wire [31:0] p2_add_79187_comb;
  wire [31:0] p2_add_79190_comb;
  wire [31:0] p2_add_79191_comb;
  wire [31:0] p2_add_79194_comb;
  wire [31:0] p2_add_79195_comb;
  wire [31:0] p2_add_79198_comb;
  wire [31:0] p2_add_79199_comb;
  wire [31:0] p2_add_79202_comb;
  wire [31:0] p2_add_79203_comb;
  wire [31:0] p2_add_79206_comb;
  wire [31:0] p2_add_79207_comb;
  wire [31:0] p2_add_79210_comb;
  wire [31:0] p2_add_79211_comb;
  wire [31:0] p2_add_79214_comb;
  wire [31:0] p2_add_79215_comb;
  wire [31:0] p2_add_79218_comb;
  wire [31:0] p2_add_79219_comb;
  wire [31:0] p2_add_79222_comb;
  wire [31:0] p2_add_79223_comb;
  wire [31:0] p2_add_79226_comb;
  wire [31:0] p2_add_79227_comb;
  wire [31:0] p2_add_79230_comb;
  wire [31:0] p2_add_79231_comb;
  wire [31:0] p2_add_79234_comb;
  wire [31:0] p2_add_79235_comb;
  wire [31:0] p2_add_79238_comb;
  wire [31:0] p2_add_79239_comb;
  wire [31:0] p2_add_79242_comb;
  wire [31:0] p2_add_79243_comb;
  wire [31:0] p2_add_79246_comb;
  wire [31:0] p2_add_79247_comb;
  wire [31:0] p2_add_79250_comb;
  wire [31:0] p2_add_79251_comb;
  wire [31:0] p2_add_79254_comb;
  wire [31:0] p2_add_79255_comb;
  wire [31:0] p2_add_79258_comb;
  wire [31:0] p2_add_79259_comb;
  wire [31:0] p2_add_79262_comb;
  wire [31:0] p2_add_79263_comb;
  wire [31:0] p2_add_79266_comb;
  wire [31:0] p2_add_79267_comb;
  wire [31:0] p2_add_79270_comb;
  wire [31:0] p2_add_79271_comb;
  wire [31:0] p2_add_79274_comb;
  wire [31:0] p2_add_79275_comb;
  wire [31:0] p2_add_79278_comb;
  wire [31:0] p2_add_79279_comb;
  wire [31:0] p2_add_79282_comb;
  wire [31:0] p2_add_79283_comb;
  wire [31:0] p2_add_79286_comb;
  wire [31:0] p2_add_79287_comb;
  wire [31:0] p2_add_79290_comb;
  wire [31:0] p2_add_79291_comb;
  wire [31:0] p2_add_79294_comb;
  wire [31:0] p2_add_79295_comb;
  wire [31:0] p2_add_79298_comb;
  wire [31:0] p2_add_79299_comb;
  wire [31:0] p2_add_79302_comb;
  wire [31:0] p2_add_79303_comb;
  wire [31:0] p2_add_79306_comb;
  wire [31:0] p2_add_79307_comb;
  wire [31:0] p2_add_79310_comb;
  wire [31:0] p2_add_79311_comb;
  wire [31:0] p2_add_79314_comb;
  wire [31:0] p2_add_79315_comb;
  wire [31:0] p2_add_79318_comb;
  wire [31:0] p2_add_79319_comb;
  wire [31:0] p2_add_79322_comb;
  wire [31:0] p2_add_79323_comb;
  wire [31:0] p2_add_79326_comb;
  wire [31:0] p2_add_79327_comb;
  wire [31:0] p2_add_79330_comb;
  wire [31:0] p2_add_79331_comb;
  wire [31:0] p2_add_79334_comb;
  wire [31:0] p2_add_79335_comb;
  wire [31:0] p2_add_79338_comb;
  wire [31:0] p2_add_79339_comb;
  wire [31:0] p2_add_79342_comb;
  wire [31:0] p2_add_79343_comb;
  wire [31:0] p2_add_79346_comb;
  wire [31:0] p2_add_79347_comb;
  wire [31:0] p2_add_79350_comb;
  wire [31:0] p2_add_79351_comb;
  wire [31:0] p2_add_79354_comb;
  wire [31:0] p2_add_79355_comb;
  wire [31:0] p2_add_79358_comb;
  wire [31:0] p2_add_79359_comb;
  wire [31:0] p2_add_79362_comb;
  wire [31:0] p2_add_79363_comb;
  wire [31:0] p2_add_79366_comb;
  wire [31:0] p2_add_79367_comb;
  wire [31:0] p2_add_79370_comb;
  wire [31:0] p2_add_79371_comb;
  wire [31:0] p2_add_79374_comb;
  wire [31:0] p2_add_79375_comb;
  wire [31:0] p2_add_79378_comb;
  wire [31:0] p2_add_79379_comb;
  wire [31:0] p2_add_79382_comb;
  wire [31:0] p2_add_79383_comb;
  wire [31:0] p2_add_79386_comb;
  wire [31:0] p2_add_79387_comb;
  wire [31:0] p2_add_79390_comb;
  wire [31:0] p2_add_79391_comb;
  wire [31:0] p2_add_79394_comb;
  wire [31:0] p2_add_79395_comb;
  wire [31:0] p2_add_79398_comb;
  wire [31:0] p2_add_79399_comb;
  wire [31:0] p2_add_79402_comb;
  wire [31:0] p2_add_79403_comb;
  wire [31:0] p2_add_79406_comb;
  wire [31:0] p2_add_79407_comb;
  wire [31:0] p2_add_79410_comb;
  wire [31:0] p2_add_79411_comb;
  wire [31:0] p2_add_79414_comb;
  wire [31:0] p2_add_79415_comb;
  wire [31:0] p2_add_79418_comb;
  wire [31:0] p2_add_79419_comb;
  wire [31:0] p2_add_79422_comb;
  wire [31:0] p2_add_79423_comb;
  wire [31:0] p2_add_79426_comb;
  wire [31:0] p2_add_79427_comb;
  wire [31:0] p2_add_79430_comb;
  wire [31:0] p2_add_79431_comb;
  wire [31:0] p2_add_79434_comb;
  wire [31:0] p2_add_79435_comb;
  wire [31:0] p2_add_79438_comb;
  wire [31:0] p2_add_79439_comb;
  wire [31:0] p2_add_79442_comb;
  wire [31:0] p2_add_79443_comb;
  wire [31:0] p2_add_79446_comb;
  wire [31:0] p2_add_79447_comb;
  wire [31:0] p2_add_79450_comb;
  wire [31:0] p2_add_79451_comb;
  wire [31:0] p2_add_79454_comb;
  wire [31:0] p2_add_79455_comb;
  wire [31:0] p2_add_79458_comb;
  wire [31:0] p2_add_79459_comb;
  wire [31:0] p2_add_79462_comb;
  wire [31:0] p2_add_79463_comb;
  wire [31:0] p2_add_79466_comb;
  wire [31:0] p2_add_79467_comb;
  wire [31:0] p2_add_79470_comb;
  wire [31:0] p2_add_79471_comb;
  wire [31:0] p2_add_79474_comb;
  wire [31:0] p2_add_79475_comb;
  wire [31:0] p2_add_79478_comb;
  wire [31:0] p2_add_79479_comb;
  wire [31:0] p2_add_79482_comb;
  wire [31:0] p2_add_79483_comb;
  wire [31:0] p2_add_79486_comb;
  wire [31:0] p2_add_79487_comb;
  wire [31:0] p2_add_79490_comb;
  wire [31:0] p2_add_79491_comb;
  wire [31:0] p2_add_79494_comb;
  wire [31:0] p2_add_79495_comb;
  wire [31:0] p2_add_79498_comb;
  wire [31:0] p2_add_79499_comb;
  wire [31:0] p2_add_79502_comb;
  wire [31:0] p2_add_79503_comb;
  wire [31:0] p2_add_79506_comb;
  wire [31:0] p2_add_79507_comb;
  wire [31:0] p2_add_79510_comb;
  wire [31:0] p2_add_79511_comb;
  wire [31:0] p2_add_79514_comb;
  wire [31:0] p2_add_79515_comb;
  wire [31:0] p2_add_79518_comb;
  wire [31:0] p2_add_79519_comb;
  wire [31:0] p2_add_79522_comb;
  wire [31:0] p2_add_79523_comb;
  wire [31:0] p2_add_79526_comb;
  wire [31:0] p2_add_79527_comb;
  wire [31:0] p2_add_79530_comb;
  wire [31:0] p2_add_79531_comb;
  wire [31:0] p2_add_79534_comb;
  wire [31:0] p2_add_79535_comb;
  wire [31:0] p2_add_79538_comb;
  wire [31:0] p2_add_79539_comb;
  wire [31:0] p2_add_79542_comb;
  wire [31:0] p2_add_79543_comb;
  wire [31:0] p2_add_79546_comb;
  wire [31:0] p2_add_79547_comb;
  wire [31:0] p2_add_79550_comb;
  wire [31:0] p2_add_79551_comb;
  wire [31:0] p2_add_79554_comb;
  wire [31:0] p2_add_79555_comb;
  wire [31:0] p2_add_79558_comb;
  wire [31:0] p2_add_79559_comb;
  wire [31:0] p2_add_79562_comb;
  wire [31:0] p2_add_79563_comb;
  wire [31:0] p2_add_79566_comb;
  wire [31:0] p2_add_79567_comb;
  wire [31:0] p2_add_79570_comb;
  wire [31:0] p2_add_79571_comb;
  wire [31:0] p2_add_79574_comb;
  wire [31:0] p2_add_79575_comb;
  wire [31:0] p2_add_79578_comb;
  wire [31:0] p2_add_79579_comb;
  wire [31:0] p2_add_79582_comb;
  wire [31:0] p2_add_79583_comb;
  wire [31:0] p2_add_79586_comb;
  wire [31:0] p2_add_79587_comb;
  wire [31:0] p2_add_79588_comb;
  wire [31:0] p2_add_79589_comb;
  wire [31:0] p2_add_79590_comb;
  wire [31:0] p2_add_79591_comb;
  wire [31:0] p2_add_79592_comb;
  wire [31:0] p2_add_79593_comb;
  wire [31:0] p2_add_79594_comb;
  wire [31:0] p2_add_79595_comb;
  wire [31:0] p2_add_79596_comb;
  wire [31:0] p2_add_79597_comb;
  wire [31:0] p2_add_79598_comb;
  wire [31:0] p2_add_79599_comb;
  wire [31:0] p2_add_79600_comb;
  wire [31:0] p2_add_79601_comb;
  wire [31:0] p2_add_79602_comb;
  wire [31:0] p2_add_79603_comb;
  wire [31:0] p2_add_79604_comb;
  wire [31:0] p2_add_79605_comb;
  wire [31:0] p2_add_79606_comb;
  wire [31:0] p2_add_79607_comb;
  wire [31:0] p2_add_79608_comb;
  wire [31:0] p2_add_79609_comb;
  wire [31:0] p2_add_79610_comb;
  wire [31:0] p2_add_79611_comb;
  wire [31:0] p2_add_79612_comb;
  wire [31:0] p2_add_79613_comb;
  wire [31:0] p2_add_79614_comb;
  wire [31:0] p2_add_79615_comb;
  wire [31:0] p2_add_79616_comb;
  wire [31:0] p2_add_79617_comb;
  wire [31:0] p2_add_79618_comb;
  wire [31:0] p2_add_79619_comb;
  wire [31:0] p2_add_79620_comb;
  wire [31:0] p2_add_79621_comb;
  wire [31:0] p2_add_79622_comb;
  wire [31:0] p2_add_79623_comb;
  wire [31:0] p2_add_79624_comb;
  wire [31:0] p2_add_79625_comb;
  wire [31:0] p2_add_79626_comb;
  wire [31:0] p2_add_79627_comb;
  wire [31:0] p2_add_79628_comb;
  wire [31:0] p2_add_79629_comb;
  wire [31:0] p2_add_79630_comb;
  wire [31:0] p2_add_79631_comb;
  wire [31:0] p2_add_79632_comb;
  wire [31:0] p2_add_79633_comb;
  wire [31:0] p2_add_79634_comb;
  wire [31:0] p2_add_79635_comb;
  wire [31:0] p2_add_79636_comb;
  wire [31:0] p2_add_79637_comb;
  wire [31:0] p2_add_79638_comb;
  wire [31:0] p2_add_79639_comb;
  wire [31:0] p2_add_79640_comb;
  wire [31:0] p2_add_79641_comb;
  wire [31:0] p2_add_79642_comb;
  wire [31:0] p2_add_79643_comb;
  wire [31:0] p2_add_79644_comb;
  wire [31:0] p2_add_79645_comb;
  wire [31:0] p2_add_79646_comb;
  wire [31:0] p2_add_79647_comb;
  wire [31:0] p2_add_79648_comb;
  wire [31:0] p2_add_79649_comb;
  wire [31:0] p2_add_79650_comb;
  wire [31:0] p2_add_79651_comb;
  wire [31:0] p2_add_79652_comb;
  wire [31:0] p2_add_79653_comb;
  wire [31:0] p2_add_79654_comb;
  wire [31:0] p2_add_79655_comb;
  wire [31:0] p2_add_79656_comb;
  wire [31:0] p2_add_79657_comb;
  wire [31:0] p2_add_79658_comb;
  wire [31:0] p2_add_79659_comb;
  wire [31:0] p2_add_79660_comb;
  wire [31:0] p2_add_79661_comb;
  wire [31:0] p2_add_79662_comb;
  wire [31:0] p2_add_79663_comb;
  wire [31:0] p2_add_79664_comb;
  wire [31:0] p2_add_79665_comb;
  wire [31:0] p2_add_79666_comb;
  wire [31:0] p2_add_79667_comb;
  wire [31:0] p2_add_79668_comb;
  wire [31:0] p2_add_79669_comb;
  wire [31:0] p2_add_79670_comb;
  wire [31:0] p2_add_79671_comb;
  wire [31:0] p2_add_79672_comb;
  wire [31:0] p2_add_79673_comb;
  wire [31:0] p2_add_79674_comb;
  wire [31:0] p2_add_79675_comb;
  wire [31:0] p2_add_79676_comb;
  wire [31:0] p2_add_79677_comb;
  wire [31:0] p2_add_79678_comb;
  wire [31:0] p2_add_79679_comb;
  wire [31:0] p2_add_79680_comb;
  wire [31:0] p2_add_79681_comb;
  wire [31:0] p2_add_79682_comb;
  wire [31:0] p2_add_79683_comb;
  wire [31:0] p2_add_79684_comb;
  wire [31:0] p2_add_79685_comb;
  assign p2_add_78986_comb = p1_smul_75972 + p1_smul_75973;
  assign p2_add_78987_comb = p1_smul_75974 + p1_smul_75975;
  assign p2_add_78988_comb = p1_smul_75976 + p1_smul_75977;
  assign p2_add_78989_comb = p1_smul_75978 + p1_smul_75979;
  assign p2_add_78990_comb = p1_smul_75980 + p1_smul_75981;
  assign p2_add_78991_comb = p1_smul_75982 + p1_smul_75983;
  assign p2_add_78992_comb = p1_smul_75984 + p1_smul_75985;
  assign p2_add_78993_comb = p1_smul_75986 + p1_smul_75987;
  assign p2_add_78994_comb = p1_smul_75988 + p1_smul_75989;
  assign p2_add_78995_comb = p1_smul_75990 + p1_smul_75991;
  assign p2_add_78996_comb = p1_smul_75992 + p1_smul_75993;
  assign p2_add_78997_comb = p1_smul_75994 + p1_smul_75995;
  assign p2_add_78998_comb = p1_smul_75996 + p1_smul_75997;
  assign p2_add_78999_comb = p1_smul_75998 + p1_smul_75999;
  assign p2_add_79000_comb = p1_smul_76000 + p1_smul_76001;
  assign p2_add_79001_comb = p1_smul_76002 + p1_smul_76003;
  assign p2_add_79002_comb = p1_smul_76004 + p1_smul_76005;
  assign p2_add_79003_comb = p1_smul_76006 + p1_smul_76007;
  assign p2_add_79004_comb = p1_smul_76008 + p1_smul_76009;
  assign p2_add_79005_comb = p1_smul_76010 + p1_smul_76011;
  assign p2_add_79006_comb = p1_smul_76012 + p1_smul_76013;
  assign p2_add_79007_comb = p1_smul_76014 + p1_smul_76015;
  assign p2_add_79008_comb = p1_smul_76016 + p1_smul_76017;
  assign p2_add_79009_comb = p1_smul_76018 + p1_smul_76019;
  assign p2_add_79010_comb = p1_smul_76020 + p1_smul_76021;
  assign p2_add_79011_comb = p1_smul_76022 + p1_smul_76023;
  assign p2_add_79012_comb = p1_smul_76024 + p1_smul_76025;
  assign p2_add_79013_comb = p1_smul_76026 + p1_smul_76027;
  assign p2_add_79014_comb = p1_smul_76028 + p1_smul_76029;
  assign p2_add_79015_comb = p1_smul_76030 + p1_smul_76031;
  assign p2_add_79016_comb = p1_smul_76032 + p1_smul_76033;
  assign p2_add_79017_comb = p1_smul_76034 + p1_smul_76035;
  assign p2_add_79018_comb = p1_smul_76036 + p1_smul_76037;
  assign p2_add_79019_comb = p1_smul_76038 + p1_smul_76039;
  assign p2_add_79020_comb = p1_smul_76040 + p1_smul_76041;
  assign p2_add_79021_comb = p1_smul_76042 + p1_smul_76043;
  assign p2_add_79022_comb = p1_smul_76044 + p1_smul_76045;
  assign p2_add_79023_comb = p1_smul_76046 + p1_smul_76047;
  assign p2_add_79024_comb = p1_smul_76048 + p1_smul_76049;
  assign p2_add_79025_comb = p1_smul_76050 + p1_smul_76051;
  assign p2_add_79026_comb = p1_smul_76052 + p1_smul_76053;
  assign p2_add_79027_comb = p1_smul_76054 + p1_smul_76055;
  assign p2_add_79028_comb = p1_smul_76056 + p1_smul_76057;
  assign p2_add_79029_comb = p1_smul_76058 + p1_smul_76059;
  assign p2_add_79030_comb = p1_smul_76060 + p1_smul_76061;
  assign p2_add_79031_comb = p1_smul_76062 + p1_smul_76063;
  assign p2_add_79032_comb = p1_smul_76064 + p1_smul_76065;
  assign p2_add_79033_comb = p1_smul_76066 + p1_smul_76067;
  assign p2_add_79034_comb = p1_smul_76068 + p1_smul_76069;
  assign p2_add_79035_comb = p1_smul_76070 + p1_smul_76071;
  assign p2_add_79036_comb = p1_smul_76072 + p1_smul_76073;
  assign p2_add_79037_comb = p1_smul_76074 + p1_smul_76075;
  assign p2_add_79038_comb = p1_smul_76076 + p1_smul_76077;
  assign p2_add_79039_comb = p1_smul_76078 + p1_smul_76079;
  assign p2_add_79040_comb = p1_smul_76080 + p1_smul_76081;
  assign p2_add_79041_comb = p1_smul_76082 + p1_smul_76083;
  assign p2_add_79042_comb = p1_smul_76084 + p1_smul_76085;
  assign p2_add_79043_comb = p1_smul_76086 + p1_smul_76087;
  assign p2_add_79044_comb = p1_smul_76088 + p1_smul_76089;
  assign p2_add_79045_comb = p1_smul_76090 + p1_smul_76091;
  assign p2_add_79046_comb = p1_smul_76092 + p1_smul_76093;
  assign p2_add_79047_comb = p1_smul_76094 + p1_smul_76095;
  assign p2_add_79048_comb = p1_smul_76096 + p1_smul_76097;
  assign p2_add_79049_comb = p1_smul_76098 + p1_smul_76099;
  assign p2_add_79050_comb = p1_smul_76100 + p1_smul_76101;
  assign p2_add_79051_comb = p1_smul_76102 + p1_smul_76103;
  assign p2_add_79052_comb = p1_smul_76104 + p1_smul_76105;
  assign p2_add_79053_comb = p1_smul_76106 + p1_smul_76107;
  assign p2_add_79054_comb = p1_smul_76108 + p1_smul_76109;
  assign p2_add_79055_comb = p1_smul_76110 + p1_smul_76111;
  assign p2_add_79056_comb = p1_smul_76112 + p1_smul_76113;
  assign p2_add_79057_comb = p1_smul_76114 + p1_smul_76115;
  assign p2_add_79058_comb = p1_smul_76116 + p1_smul_76117;
  assign p2_add_79059_comb = p1_smul_76118 + p1_smul_76119;
  assign p2_add_79060_comb = p1_smul_76120 + p1_smul_76121;
  assign p2_add_79061_comb = p1_smul_76122 + p1_smul_76123;
  assign p2_add_79062_comb = p1_smul_76124 + p1_smul_76125;
  assign p2_add_79063_comb = p1_smul_76126 + p1_smul_76127;
  assign p2_add_79064_comb = p1_smul_76128 + p1_smul_76129;
  assign p2_add_79065_comb = p1_smul_76130 + p1_smul_76131;
  assign p2_add_79066_comb = p1_smul_76132 + p1_smul_76133;
  assign p2_add_79067_comb = p1_smul_76134 + p1_smul_76135;
  assign p2_add_79068_comb = p1_smul_76136 + p1_smul_76137;
  assign p2_add_79069_comb = p1_smul_76138 + p1_smul_76139;
  assign p2_add_79070_comb = p1_smul_76140 + p1_smul_76141;
  assign p2_add_79071_comb = p1_smul_76142 + p1_smul_76143;
  assign p2_add_79072_comb = p1_smul_76144 + p1_smul_76145;
  assign p2_add_79073_comb = p1_smul_76146 + p1_smul_76147;
  assign p2_add_79074_comb = p1_smul_76148 + p1_smul_76149;
  assign p2_add_79075_comb = p1_smul_76150 + p1_smul_76151;
  assign p2_add_79076_comb = p1_smul_76152 + p1_smul_76153;
  assign p2_add_79077_comb = p1_smul_76154 + p1_smul_76155;
  assign p2_add_79078_comb = p1_smul_76156 + p1_smul_76157;
  assign p2_add_79079_comb = p1_smul_76158 + p1_smul_76159;
  assign p2_add_79080_comb = p1_smul_76160 + p1_smul_76161;
  assign p2_add_79081_comb = p1_smul_76162 + p1_smul_76163;
  assign p2_add_79082_comb = p1_smul_76164 + p1_smul_76165;
  assign p2_add_79083_comb = p1_smul_76166 + p1_smul_76167;
  assign p2_add_79084_comb = p1_smul_76168 + p1_smul_76169;
  assign p2_add_79085_comb = p1_smul_76170 + p1_smul_76171;
  assign p2_add_79086_comb = p1_smul_76172 + p1_smul_76173;
  assign p2_add_79087_comb = p1_smul_76174 + p1_smul_76175;
  assign p2_add_79088_comb = p1_smul_76176 + p1_smul_76177;
  assign p2_add_79089_comb = p1_smul_76178 + p1_smul_76179;
  assign p2_add_79090_comb = p1_smul_76180 + p1_smul_76181;
  assign p2_add_79091_comb = p1_smul_76182 + p1_smul_76183;
  assign p2_add_79092_comb = p1_smul_76184 + p1_smul_76185;
  assign p2_add_79093_comb = p1_smul_76186 + p1_smul_76187;
  assign p2_add_79094_comb = p1_smul_76188 + p1_smul_76189;
  assign p2_add_79095_comb = p1_smul_76190 + p1_smul_76191;
  assign p2_add_79096_comb = p1_smul_76192 + p1_smul_76193;
  assign p2_add_79097_comb = p1_smul_76194 + p1_smul_76195;
  assign p2_add_79098_comb = p1_smul_76196 + p1_smul_76197;
  assign p2_add_79099_comb = p1_smul_76198 + p1_smul_76199;
  assign p2_add_79100_comb = p1_smul_76200 + p1_smul_76201;
  assign p2_add_79101_comb = p1_smul_76202 + p1_smul_76203;
  assign p2_add_79102_comb = p1_smul_76204 + p1_smul_76205;
  assign p2_add_79103_comb = p1_smul_76206 + p1_smul_76207;
  assign p2_add_79104_comb = p1_smul_76208 + p1_smul_76209;
  assign p2_add_79105_comb = p1_smul_76210 + p1_smul_76211;
  assign p2_add_79106_comb = p1_smul_76212 + p1_smul_76213;
  assign p2_add_79107_comb = p1_smul_76214 + p1_smul_76215;
  assign p2_add_79108_comb = p1_smul_76216 + p1_smul_76217;
  assign p2_add_79109_comb = p1_smul_76218 + p1_smul_76219;
  assign p2_add_79110_comb = p1_smul_76220 + p1_smul_76221;
  assign p2_add_79111_comb = p1_smul_76222 + p1_smul_76223;
  assign p2_add_79112_comb = p1_smul_76224 + p1_smul_76225;
  assign p2_add_79113_comb = p1_smul_76226 + p1_smul_76227;
  assign p2_add_79114_comb = p1_smul_76228 + p1_smul_76229;
  assign p2_add_79115_comb = p1_smul_76230 + p1_smul_76231;
  assign p2_add_79116_comb = p1_smul_76232 + p1_smul_76233;
  assign p2_add_79117_comb = p1_smul_76234 + p1_smul_76235;
  assign p2_add_79118_comb = p1_smul_76236 + p1_smul_76237;
  assign p2_add_79119_comb = p1_smul_76238 + p1_smul_76239;
  assign p2_add_79120_comb = p1_smul_76240 + p1_smul_76241;
  assign p2_add_79121_comb = p1_smul_76242 + p1_smul_76243;
  assign p2_add_79122_comb = p1_smul_76244 + p1_smul_76245;
  assign p2_add_79123_comb = p1_smul_76246 + p1_smul_76247;
  assign p2_add_79124_comb = p1_smul_76248 + p1_smul_76249;
  assign p2_add_79125_comb = p1_smul_76250 + p1_smul_76251;
  assign p2_add_79126_comb = p1_smul_76252 + p1_smul_76253;
  assign p2_add_79127_comb = p1_smul_76254 + p1_smul_76255;
  assign p2_add_79128_comb = p1_smul_76256 + p1_smul_76257;
  assign p2_add_79129_comb = p1_smul_76258 + p1_smul_76259;
  assign p2_add_79130_comb = p1_smul_76260 + p1_smul_76261;
  assign p2_add_79131_comb = p1_smul_76262 + p1_smul_76263;
  assign p2_add_79132_comb = p1_smul_76264 + p1_smul_76265;
  assign p2_add_79133_comb = p1_smul_76266 + p1_smul_76267;
  assign p2_add_79134_comb = p1_smul_76268 + p1_smul_76269;
  assign p2_add_79135_comb = p1_smul_76270 + p1_smul_76271;
  assign p2_add_79136_comb = p1_smul_76272 + p1_smul_76273;
  assign p2_add_79137_comb = p1_smul_76274 + p1_smul_76275;
  assign p2_add_79138_comb = p1_smul_76276 + p1_smul_76277;
  assign p2_add_79139_comb = p1_smul_76278 + p1_smul_76279;
  assign p2_add_79140_comb = p1_smul_76280 + p1_smul_76281;
  assign p2_add_79141_comb = p1_smul_76282 + p1_smul_76283;
  assign p2_add_79142_comb = p1_smul_76284 + p1_smul_76285;
  assign p2_add_79143_comb = p1_smul_76286 + p1_smul_76287;
  assign p2_add_79144_comb = p1_smul_76288 + p1_smul_76289;
  assign p2_add_79145_comb = p1_smul_76290 + p1_smul_76291;
  assign p2_add_79146_comb = p1_smul_76292 + p1_smul_76293;
  assign p2_add_79147_comb = p1_smul_76294 + p1_smul_76295;
  assign p2_add_79148_comb = p1_smul_76296 + p1_smul_76297;
  assign p2_add_79149_comb = p1_smul_76298 + p1_smul_76299;
  assign p2_add_79150_comb = p1_smul_76300 + p1_smul_76301;
  assign p2_add_79151_comb = p1_smul_76302 + p1_smul_76303;
  assign p2_add_79152_comb = p1_smul_76304 + p1_smul_76305;
  assign p2_add_79153_comb = p1_smul_76306 + p1_smul_76307;
  assign p2_add_79154_comb = p1_smul_76308 + p1_smul_76309;
  assign p2_add_79155_comb = p1_smul_76310 + p1_smul_76311;
  assign p2_add_79156_comb = p1_smul_76312 + p1_smul_76313;
  assign p2_add_79157_comb = p1_smul_76314 + p1_smul_76315;
  assign p2_add_79158_comb = p1_smul_76316 + p1_smul_76317;
  assign p2_add_79159_comb = p1_smul_76318 + p1_smul_76319;
  assign p2_add_79160_comb = p1_smul_76320 + p1_smul_76321;
  assign p2_add_79161_comb = p1_smul_76322 + p1_smul_76323;
  assign p2_add_79162_comb = p1_smul_76324 + p1_smul_76325;
  assign p2_add_79163_comb = p1_smul_76326 + p1_smul_76327;
  assign p2_add_79164_comb = p1_smul_76328 + p1_smul_76329;
  assign p2_add_79165_comb = p1_smul_76330 + p1_smul_76331;
  assign p2_add_79166_comb = p1_smul_76332 + p1_smul_76333;
  assign p2_add_79167_comb = p1_smul_76334 + p1_smul_76335;
  assign p2_add_79168_comb = p1_smul_76336 + p1_smul_76337;
  assign p2_add_79169_comb = p1_smul_76338 + p1_smul_76339;
  assign p2_add_79170_comb = p1_smul_76340 + p1_smul_76341;
  assign p2_add_79171_comb = p1_smul_76342 + p1_smul_76343;
  assign p2_add_79172_comb = p1_smul_76344 + p1_smul_76345;
  assign p2_add_79173_comb = p1_smul_76346 + p1_smul_76347;
  assign p2_add_79174_comb = p1_smul_76348 + p1_smul_76349;
  assign p2_add_79175_comb = p1_smul_76350 + p1_smul_76351;
  assign p2_add_79176_comb = p1_smul_76352 + p1_smul_76353;
  assign p2_add_79177_comb = p1_smul_76354 + p1_smul_76355;
  assign p2_add_79178_comb = p1_smul_76356 + p1_smul_76357;
  assign p2_add_79179_comb = p1_smul_76358 + p1_smul_76359;
  assign p2_add_79180_comb = p1_smul_76360 + p1_smul_76361;
  assign p2_add_79181_comb = p1_smul_76362 + p1_smul_76363;
  assign p2_add_79182_comb = p1_smul_76364 + p1_smul_76365;
  assign p2_add_79183_comb = p1_smul_76366 + p1_smul_76367;
  assign p2_add_79184_comb = p1_smul_76368 + p1_smul_76369;
  assign p2_add_79185_comb = p1_smul_76370 + p1_smul_76371;
  assign p2_add_79188_comb = p1_smul_76374 + p1_smul_76375;
  assign p2_add_79189_comb = p1_smul_76376 + p1_smul_76377;
  assign p2_add_79192_comb = p1_smul_76380 + p1_smul_76381;
  assign p2_add_79193_comb = p1_smul_76382 + p1_smul_76383;
  assign p2_add_79196_comb = p1_smul_76386 + p1_smul_76387;
  assign p2_add_79197_comb = p1_smul_76388 + p1_smul_76389;
  assign p2_add_79200_comb = p1_smul_76392 + p1_smul_76393;
  assign p2_add_79201_comb = p1_smul_76394 + p1_smul_76395;
  assign p2_add_79204_comb = p1_smul_76398 + p1_smul_76399;
  assign p2_add_79205_comb = p1_smul_76400 + p1_smul_76401;
  assign p2_add_79208_comb = p1_smul_76404 + p1_smul_76405;
  assign p2_add_79209_comb = p1_smul_76406 + p1_smul_76407;
  assign p2_add_79212_comb = p1_smul_76410 + p1_smul_76411;
  assign p2_add_79213_comb = p1_smul_76412 + p1_smul_76413;
  assign p2_add_79216_comb = p1_smul_76416 + p1_smul_76417;
  assign p2_add_79217_comb = p1_smul_76418 + p1_smul_76419;
  assign p2_add_79220_comb = p1_smul_76422 + p1_smul_76423;
  assign p2_add_79221_comb = p1_smul_76424 + p1_smul_76425;
  assign p2_add_79224_comb = p1_smul_76428 + p1_smul_76429;
  assign p2_add_79225_comb = p1_smul_76430 + p1_smul_76431;
  assign p2_add_79228_comb = p1_smul_76434 + p1_smul_76435;
  assign p2_add_79229_comb = p1_smul_76436 + p1_smul_76437;
  assign p2_add_79232_comb = p1_smul_76440 + p1_smul_76441;
  assign p2_add_79233_comb = p1_smul_76442 + p1_smul_76443;
  assign p2_add_79236_comb = p1_smul_76446 + p1_smul_76447;
  assign p2_add_79237_comb = p1_smul_76448 + p1_smul_76449;
  assign p2_add_79240_comb = p1_smul_76452 + p1_smul_76453;
  assign p2_add_79241_comb = p1_smul_76454 + p1_smul_76455;
  assign p2_add_79244_comb = p1_smul_76458 + p1_smul_76459;
  assign p2_add_79245_comb = p1_smul_76460 + p1_smul_76461;
  assign p2_add_79248_comb = p1_smul_76464 + p1_smul_76465;
  assign p2_add_79249_comb = p1_smul_76466 + p1_smul_76467;
  assign p2_add_79252_comb = p1_smul_76470 + p1_smul_76471;
  assign p2_add_79253_comb = p1_smul_76472 + p1_smul_76473;
  assign p2_add_79256_comb = p1_smul_76476 + p1_smul_76477;
  assign p2_add_79257_comb = p1_smul_76478 + p1_smul_76479;
  assign p2_add_79260_comb = p1_smul_76482 + p1_smul_76483;
  assign p2_add_79261_comb = p1_smul_76484 + p1_smul_76485;
  assign p2_add_79264_comb = p1_smul_76488 + p1_smul_76489;
  assign p2_add_79265_comb = p1_smul_76490 + p1_smul_76491;
  assign p2_add_79268_comb = p1_smul_76494 + p1_smul_76495;
  assign p2_add_79269_comb = p1_smul_76496 + p1_smul_76497;
  assign p2_add_79272_comb = p1_smul_76500 + p1_smul_76501;
  assign p2_add_79273_comb = p1_smul_76502 + p1_smul_76503;
  assign p2_add_79276_comb = p1_smul_76506 + p1_smul_76507;
  assign p2_add_79277_comb = p1_smul_76508 + p1_smul_76509;
  assign p2_add_79280_comb = p1_smul_76512 + p1_smul_76513;
  assign p2_add_79281_comb = p1_smul_76514 + p1_smul_76515;
  assign p2_add_79284_comb = p1_smul_76518 + p1_smul_76519;
  assign p2_add_79285_comb = p1_smul_76520 + p1_smul_76521;
  assign p2_add_79288_comb = p1_smul_76524 + p1_smul_76525;
  assign p2_add_79289_comb = p1_smul_76526 + p1_smul_76527;
  assign p2_add_79292_comb = p1_smul_76530 + p1_smul_76531;
  assign p2_add_79293_comb = p1_smul_76532 + p1_smul_76533;
  assign p2_add_79296_comb = p1_smul_76536 + p1_smul_76537;
  assign p2_add_79297_comb = p1_smul_76538 + p1_smul_76539;
  assign p2_add_79300_comb = p1_smul_76542 + p1_smul_76543;
  assign p2_add_79301_comb = p1_smul_76544 + p1_smul_76545;
  assign p2_add_79304_comb = p1_smul_76548 + p1_smul_76549;
  assign p2_add_79305_comb = p1_smul_76550 + p1_smul_76551;
  assign p2_add_79308_comb = p1_smul_76554 + p1_smul_76555;
  assign p2_add_79309_comb = p1_smul_76556 + p1_smul_76557;
  assign p2_add_79312_comb = p1_smul_76560 + p1_smul_76561;
  assign p2_add_79313_comb = p1_smul_76562 + p1_smul_76563;
  assign p2_add_79316_comb = p1_smul_76566 + p1_smul_76567;
  assign p2_add_79317_comb = p1_smul_76568 + p1_smul_76569;
  assign p2_add_79320_comb = p1_smul_76572 + p1_smul_76573;
  assign p2_add_79321_comb = p1_smul_76574 + p1_smul_76575;
  assign p2_add_79324_comb = p1_smul_76578 + p1_smul_76579;
  assign p2_add_79325_comb = p1_smul_76580 + p1_smul_76581;
  assign p2_add_79328_comb = p1_smul_76584 + p1_smul_76585;
  assign p2_add_79329_comb = p1_smul_76586 + p1_smul_76587;
  assign p2_add_79332_comb = p1_smul_76590 + p1_smul_76591;
  assign p2_add_79333_comb = p1_smul_76592 + p1_smul_76593;
  assign p2_add_79336_comb = p1_smul_76596 + p1_smul_76597;
  assign p2_add_79337_comb = p1_smul_76598 + p1_smul_76599;
  assign p2_add_79340_comb = p1_smul_76602 + p1_smul_76603;
  assign p2_add_79341_comb = p1_smul_76604 + p1_smul_76605;
  assign p2_add_79344_comb = p1_smul_76608 + p1_smul_76609;
  assign p2_add_79345_comb = p1_smul_76610 + p1_smul_76611;
  assign p2_add_79348_comb = p1_smul_76614 + p1_smul_76615;
  assign p2_add_79349_comb = p1_smul_76616 + p1_smul_76617;
  assign p2_add_79352_comb = p1_smul_76620 + p1_smul_76621;
  assign p2_add_79353_comb = p1_smul_76622 + p1_smul_76623;
  assign p2_add_79356_comb = p1_smul_76626 + p1_smul_76627;
  assign p2_add_79357_comb = p1_smul_76628 + p1_smul_76629;
  assign p2_add_79360_comb = p1_smul_76632 + p1_smul_76633;
  assign p2_add_79361_comb = p1_smul_76634 + p1_smul_76635;
  assign p2_add_79364_comb = p1_smul_76638 + p1_smul_76639;
  assign p2_add_79365_comb = p1_smul_76640 + p1_smul_76641;
  assign p2_add_79368_comb = p1_smul_76644 + p1_smul_76645;
  assign p2_add_79369_comb = p1_smul_76646 + p1_smul_76647;
  assign p2_add_79372_comb = p1_smul_76650 + p1_smul_76651;
  assign p2_add_79373_comb = p1_smul_76652 + p1_smul_76653;
  assign p2_add_79376_comb = p1_smul_76656 + p1_smul_76657;
  assign p2_add_79377_comb = p1_smul_76658 + p1_smul_76659;
  assign p2_add_79380_comb = p1_smul_76662 + p1_smul_76663;
  assign p2_add_79381_comb = p1_smul_76664 + p1_smul_76665;
  assign p2_add_79384_comb = p1_smul_76668 + p1_smul_76669;
  assign p2_add_79385_comb = p1_smul_76670 + p1_smul_76671;
  assign p2_add_79388_comb = p1_smul_76674 + p1_smul_76675;
  assign p2_add_79389_comb = p1_smul_76676 + p1_smul_76677;
  assign p2_add_79392_comb = p1_smul_76680 + p1_smul_76681;
  assign p2_add_79393_comb = p1_smul_76682 + p1_smul_76683;
  assign p2_add_79396_comb = p1_smul_76686 + p1_smul_76687;
  assign p2_add_79397_comb = p1_smul_76688 + p1_smul_76689;
  assign p2_add_79400_comb = p1_smul_76692 + p1_smul_76693;
  assign p2_add_79401_comb = p1_smul_76694 + p1_smul_76695;
  assign p2_add_79404_comb = p1_smul_76698 + p1_smul_76699;
  assign p2_add_79405_comb = p1_smul_76700 + p1_smul_76701;
  assign p2_add_79408_comb = p1_smul_76704 + p1_smul_76705;
  assign p2_add_79409_comb = p1_smul_76706 + p1_smul_76707;
  assign p2_add_79412_comb = p1_smul_76710 + p1_smul_76711;
  assign p2_add_79413_comb = p1_smul_76712 + p1_smul_76713;
  assign p2_add_79416_comb = p1_smul_76716 + p1_smul_76717;
  assign p2_add_79417_comb = p1_smul_76718 + p1_smul_76719;
  assign p2_add_79420_comb = p1_smul_76722 + p1_smul_76723;
  assign p2_add_79421_comb = p1_smul_76724 + p1_smul_76725;
  assign p2_add_79424_comb = p1_smul_76728 + p1_smul_76729;
  assign p2_add_79425_comb = p1_smul_76730 + p1_smul_76731;
  assign p2_add_79428_comb = p1_smul_76734 + p1_smul_76735;
  assign p2_add_79429_comb = p1_smul_76736 + p1_smul_76737;
  assign p2_add_79432_comb = p1_smul_76740 + p1_smul_76741;
  assign p2_add_79433_comb = p1_smul_76742 + p1_smul_76743;
  assign p2_add_79436_comb = p1_smul_76746 + p1_smul_76747;
  assign p2_add_79437_comb = p1_smul_76748 + p1_smul_76749;
  assign p2_add_79440_comb = p1_smul_76752 + p1_smul_76753;
  assign p2_add_79441_comb = p1_smul_76754 + p1_smul_76755;
  assign p2_add_79444_comb = p1_smul_76758 + p1_smul_76759;
  assign p2_add_79445_comb = p1_smul_76760 + p1_smul_76761;
  assign p2_add_79448_comb = p1_smul_76764 + p1_smul_76765;
  assign p2_add_79449_comb = p1_smul_76766 + p1_smul_76767;
  assign p2_add_79452_comb = p1_smul_76770 + p1_smul_76771;
  assign p2_add_79453_comb = p1_smul_76772 + p1_smul_76773;
  assign p2_add_79456_comb = p1_smul_76776 + p1_smul_76777;
  assign p2_add_79457_comb = p1_smul_76778 + p1_smul_76779;
  assign p2_add_79460_comb = p1_smul_76782 + p1_smul_76783;
  assign p2_add_79461_comb = p1_smul_76784 + p1_smul_76785;
  assign p2_add_79464_comb = p1_smul_76788 + p1_smul_76789;
  assign p2_add_79465_comb = p1_smul_76790 + p1_smul_76791;
  assign p2_add_79468_comb = p1_smul_76794 + p1_smul_76795;
  assign p2_add_79469_comb = p1_smul_76796 + p1_smul_76797;
  assign p2_add_79472_comb = p1_smul_76800 + p1_smul_76801;
  assign p2_add_79473_comb = p1_smul_76802 + p1_smul_76803;
  assign p2_add_79476_comb = p1_smul_76806 + p1_smul_76807;
  assign p2_add_79477_comb = p1_smul_76808 + p1_smul_76809;
  assign p2_add_79480_comb = p1_smul_76812 + p1_smul_76813;
  assign p2_add_79481_comb = p1_smul_76814 + p1_smul_76815;
  assign p2_add_79484_comb = p1_smul_76818 + p1_smul_76819;
  assign p2_add_79485_comb = p1_smul_76820 + p1_smul_76821;
  assign p2_add_79488_comb = p1_smul_76824 + p1_smul_76825;
  assign p2_add_79489_comb = p1_smul_76826 + p1_smul_76827;
  assign p2_add_79492_comb = p1_smul_76830 + p1_smul_76831;
  assign p2_add_79493_comb = p1_smul_76832 + p1_smul_76833;
  assign p2_add_79496_comb = p1_smul_76836 + p1_smul_76837;
  assign p2_add_79497_comb = p1_smul_76838 + p1_smul_76839;
  assign p2_add_79500_comb = p1_smul_76842 + p1_smul_76843;
  assign p2_add_79501_comb = p1_smul_76844 + p1_smul_76845;
  assign p2_add_79504_comb = p1_smul_76848 + p1_smul_76849;
  assign p2_add_79505_comb = p1_smul_76850 + p1_smul_76851;
  assign p2_add_79508_comb = p1_smul_76854 + p1_smul_76855;
  assign p2_add_79509_comb = p1_smul_76856 + p1_smul_76857;
  assign p2_add_79512_comb = p1_smul_76860 + p1_smul_76861;
  assign p2_add_79513_comb = p1_smul_76862 + p1_smul_76863;
  assign p2_add_79516_comb = p1_smul_76866 + p1_smul_76867;
  assign p2_add_79517_comb = p1_smul_76868 + p1_smul_76869;
  assign p2_add_79520_comb = p1_smul_76872 + p1_smul_76873;
  assign p2_add_79521_comb = p1_smul_76874 + p1_smul_76875;
  assign p2_add_79524_comb = p1_smul_76878 + p1_smul_76879;
  assign p2_add_79525_comb = p1_smul_76880 + p1_smul_76881;
  assign p2_add_79528_comb = p1_smul_76884 + p1_smul_76885;
  assign p2_add_79529_comb = p1_smul_76886 + p1_smul_76887;
  assign p2_add_79532_comb = p1_smul_76890 + p1_smul_76891;
  assign p2_add_79533_comb = p1_smul_76892 + p1_smul_76893;
  assign p2_add_79536_comb = p1_smul_76896 + p1_smul_76897;
  assign p2_add_79537_comb = p1_smul_76898 + p1_smul_76899;
  assign p2_add_79540_comb = p1_smul_76902 + p1_smul_76903;
  assign p2_add_79541_comb = p1_smul_76904 + p1_smul_76905;
  assign p2_add_79544_comb = p1_smul_76908 + p1_smul_76909;
  assign p2_add_79545_comb = p1_smul_76910 + p1_smul_76911;
  assign p2_add_79548_comb = p1_smul_76914 + p1_smul_76915;
  assign p2_add_79549_comb = p1_smul_76916 + p1_smul_76917;
  assign p2_add_79552_comb = p1_smul_76920 + p1_smul_76921;
  assign p2_add_79553_comb = p1_smul_76922 + p1_smul_76923;
  assign p2_add_79556_comb = p1_smul_76926 + p1_smul_76927;
  assign p2_add_79557_comb = p1_smul_76928 + p1_smul_76929;
  assign p2_add_79560_comb = p1_smul_76932 + p1_smul_76933;
  assign p2_add_79561_comb = p1_smul_76934 + p1_smul_76935;
  assign p2_add_79564_comb = p1_smul_76938 + p1_smul_76939;
  assign p2_add_79565_comb = p1_smul_76940 + p1_smul_76941;
  assign p2_add_79568_comb = p1_smul_76944 + p1_smul_76945;
  assign p2_add_79569_comb = p1_smul_76946 + p1_smul_76947;
  assign p2_add_79572_comb = p1_smul_76950 + p1_smul_76951;
  assign p2_add_79573_comb = p1_smul_76952 + p1_smul_76953;
  assign p2_add_79576_comb = p1_smul_76956 + p1_smul_76957;
  assign p2_add_79577_comb = p1_smul_76958 + p1_smul_76959;
  assign p2_add_79580_comb = p1_smul_76962 + p1_smul_76963;
  assign p2_add_79581_comb = p1_smul_76964 + p1_smul_76965;
  assign p2_add_79584_comb = p1_smul_76968 + p1_smul_76969;
  assign p2_add_79585_comb = p1_smul_76970 + p1_smul_76971;
  assign p2_add_79186_comb = p2_add_78986_comb + p2_add_78987_comb;
  assign p2_add_79187_comb = p1_smul_76372 + p1_smul_76373;
  assign p2_add_79190_comb = p2_add_78988_comb + p2_add_78989_comb;
  assign p2_add_79191_comb = p1_smul_76378 + p1_smul_76379;
  assign p2_add_79194_comb = p2_add_78990_comb + p2_add_78991_comb;
  assign p2_add_79195_comb = p1_smul_76384 + p1_smul_76385;
  assign p2_add_79198_comb = p2_add_78992_comb + p2_add_78993_comb;
  assign p2_add_79199_comb = p1_smul_76390 + p1_smul_76391;
  assign p2_add_79202_comb = p2_add_78994_comb + p2_add_78995_comb;
  assign p2_add_79203_comb = p1_smul_76396 + p1_smul_76397;
  assign p2_add_79206_comb = p2_add_78996_comb + p2_add_78997_comb;
  assign p2_add_79207_comb = p1_smul_76402 + p1_smul_76403;
  assign p2_add_79210_comb = p2_add_78998_comb + p2_add_78999_comb;
  assign p2_add_79211_comb = p1_smul_76408 + p1_smul_76409;
  assign p2_add_79214_comb = p2_add_79000_comb + p2_add_79001_comb;
  assign p2_add_79215_comb = p1_smul_76414 + p1_smul_76415;
  assign p2_add_79218_comb = p2_add_79002_comb + p2_add_79003_comb;
  assign p2_add_79219_comb = p1_smul_76420 + p1_smul_76421;
  assign p2_add_79222_comb = p2_add_79004_comb + p2_add_79005_comb;
  assign p2_add_79223_comb = p1_smul_76426 + p1_smul_76427;
  assign p2_add_79226_comb = p2_add_79006_comb + p2_add_79007_comb;
  assign p2_add_79227_comb = p1_smul_76432 + p1_smul_76433;
  assign p2_add_79230_comb = p2_add_79008_comb + p2_add_79009_comb;
  assign p2_add_79231_comb = p1_smul_76438 + p1_smul_76439;
  assign p2_add_79234_comb = p2_add_79010_comb + p2_add_79011_comb;
  assign p2_add_79235_comb = p1_smul_76444 + p1_smul_76445;
  assign p2_add_79238_comb = p2_add_79012_comb + p2_add_79013_comb;
  assign p2_add_79239_comb = p1_smul_76450 + p1_smul_76451;
  assign p2_add_79242_comb = p2_add_79014_comb + p2_add_79015_comb;
  assign p2_add_79243_comb = p1_smul_76456 + p1_smul_76457;
  assign p2_add_79246_comb = p2_add_79016_comb + p2_add_79017_comb;
  assign p2_add_79247_comb = p1_smul_76462 + p1_smul_76463;
  assign p2_add_79250_comb = p2_add_79018_comb + p2_add_79019_comb;
  assign p2_add_79251_comb = p1_smul_76468 + p1_smul_76469;
  assign p2_add_79254_comb = p2_add_79020_comb + p2_add_79021_comb;
  assign p2_add_79255_comb = p1_smul_76474 + p1_smul_76475;
  assign p2_add_79258_comb = p2_add_79022_comb + p2_add_79023_comb;
  assign p2_add_79259_comb = p1_smul_76480 + p1_smul_76481;
  assign p2_add_79262_comb = p2_add_79024_comb + p2_add_79025_comb;
  assign p2_add_79263_comb = p1_smul_76486 + p1_smul_76487;
  assign p2_add_79266_comb = p2_add_79026_comb + p2_add_79027_comb;
  assign p2_add_79267_comb = p1_smul_76492 + p1_smul_76493;
  assign p2_add_79270_comb = p2_add_79028_comb + p2_add_79029_comb;
  assign p2_add_79271_comb = p1_smul_76498 + p1_smul_76499;
  assign p2_add_79274_comb = p2_add_79030_comb + p2_add_79031_comb;
  assign p2_add_79275_comb = p1_smul_76504 + p1_smul_76505;
  assign p2_add_79278_comb = p2_add_79032_comb + p2_add_79033_comb;
  assign p2_add_79279_comb = p1_smul_76510 + p1_smul_76511;
  assign p2_add_79282_comb = p2_add_79034_comb + p2_add_79035_comb;
  assign p2_add_79283_comb = p1_smul_76516 + p1_smul_76517;
  assign p2_add_79286_comb = p2_add_79036_comb + p2_add_79037_comb;
  assign p2_add_79287_comb = p1_smul_76522 + p1_smul_76523;
  assign p2_add_79290_comb = p2_add_79038_comb + p2_add_79039_comb;
  assign p2_add_79291_comb = p1_smul_76528 + p1_smul_76529;
  assign p2_add_79294_comb = p2_add_79040_comb + p2_add_79041_comb;
  assign p2_add_79295_comb = p1_smul_76534 + p1_smul_76535;
  assign p2_add_79298_comb = p2_add_79042_comb + p2_add_79043_comb;
  assign p2_add_79299_comb = p1_smul_76540 + p1_smul_76541;
  assign p2_add_79302_comb = p2_add_79044_comb + p2_add_79045_comb;
  assign p2_add_79303_comb = p1_smul_76546 + p1_smul_76547;
  assign p2_add_79306_comb = p2_add_79046_comb + p2_add_79047_comb;
  assign p2_add_79307_comb = p1_smul_76552 + p1_smul_76553;
  assign p2_add_79310_comb = p2_add_79048_comb + p2_add_79049_comb;
  assign p2_add_79311_comb = p1_smul_76558 + p1_smul_76559;
  assign p2_add_79314_comb = p2_add_79050_comb + p2_add_79051_comb;
  assign p2_add_79315_comb = p1_smul_76564 + p1_smul_76565;
  assign p2_add_79318_comb = p2_add_79052_comb + p2_add_79053_comb;
  assign p2_add_79319_comb = p1_smul_76570 + p1_smul_76571;
  assign p2_add_79322_comb = p2_add_79054_comb + p2_add_79055_comb;
  assign p2_add_79323_comb = p1_smul_76576 + p1_smul_76577;
  assign p2_add_79326_comb = p2_add_79056_comb + p2_add_79057_comb;
  assign p2_add_79327_comb = p1_smul_76582 + p1_smul_76583;
  assign p2_add_79330_comb = p2_add_79058_comb + p2_add_79059_comb;
  assign p2_add_79331_comb = p1_smul_76588 + p1_smul_76589;
  assign p2_add_79334_comb = p2_add_79060_comb + p2_add_79061_comb;
  assign p2_add_79335_comb = p1_smul_76594 + p1_smul_76595;
  assign p2_add_79338_comb = p2_add_79062_comb + p2_add_79063_comb;
  assign p2_add_79339_comb = p1_smul_76600 + p1_smul_76601;
  assign p2_add_79342_comb = p2_add_79064_comb + p2_add_79065_comb;
  assign p2_add_79343_comb = p1_smul_76606 + p1_smul_76607;
  assign p2_add_79346_comb = p2_add_79066_comb + p2_add_79067_comb;
  assign p2_add_79347_comb = p1_smul_76612 + p1_smul_76613;
  assign p2_add_79350_comb = p2_add_79068_comb + p2_add_79069_comb;
  assign p2_add_79351_comb = p1_smul_76618 + p1_smul_76619;
  assign p2_add_79354_comb = p2_add_79070_comb + p2_add_79071_comb;
  assign p2_add_79355_comb = p1_smul_76624 + p1_smul_76625;
  assign p2_add_79358_comb = p2_add_79072_comb + p2_add_79073_comb;
  assign p2_add_79359_comb = p1_smul_76630 + p1_smul_76631;
  assign p2_add_79362_comb = p2_add_79074_comb + p2_add_79075_comb;
  assign p2_add_79363_comb = p1_smul_76636 + p1_smul_76637;
  assign p2_add_79366_comb = p2_add_79076_comb + p2_add_79077_comb;
  assign p2_add_79367_comb = p1_smul_76642 + p1_smul_76643;
  assign p2_add_79370_comb = p2_add_79078_comb + p2_add_79079_comb;
  assign p2_add_79371_comb = p1_smul_76648 + p1_smul_76649;
  assign p2_add_79374_comb = p2_add_79080_comb + p2_add_79081_comb;
  assign p2_add_79375_comb = p1_smul_76654 + p1_smul_76655;
  assign p2_add_79378_comb = p2_add_79082_comb + p2_add_79083_comb;
  assign p2_add_79379_comb = p1_smul_76660 + p1_smul_76661;
  assign p2_add_79382_comb = p2_add_79084_comb + p2_add_79085_comb;
  assign p2_add_79383_comb = p1_smul_76666 + p1_smul_76667;
  assign p2_add_79386_comb = p2_add_79086_comb + p2_add_79087_comb;
  assign p2_add_79387_comb = p1_smul_76672 + p1_smul_76673;
  assign p2_add_79390_comb = p2_add_79088_comb + p2_add_79089_comb;
  assign p2_add_79391_comb = p1_smul_76678 + p1_smul_76679;
  assign p2_add_79394_comb = p2_add_79090_comb + p2_add_79091_comb;
  assign p2_add_79395_comb = p1_smul_76684 + p1_smul_76685;
  assign p2_add_79398_comb = p2_add_79092_comb + p2_add_79093_comb;
  assign p2_add_79399_comb = p1_smul_76690 + p1_smul_76691;
  assign p2_add_79402_comb = p2_add_79094_comb + p2_add_79095_comb;
  assign p2_add_79403_comb = p1_smul_76696 + p1_smul_76697;
  assign p2_add_79406_comb = p2_add_79096_comb + p2_add_79097_comb;
  assign p2_add_79407_comb = p1_smul_76702 + p1_smul_76703;
  assign p2_add_79410_comb = p2_add_79098_comb + p2_add_79099_comb;
  assign p2_add_79411_comb = p1_smul_76708 + p1_smul_76709;
  assign p2_add_79414_comb = p2_add_79100_comb + p2_add_79101_comb;
  assign p2_add_79415_comb = p1_smul_76714 + p1_smul_76715;
  assign p2_add_79418_comb = p2_add_79102_comb + p2_add_79103_comb;
  assign p2_add_79419_comb = p1_smul_76720 + p1_smul_76721;
  assign p2_add_79422_comb = p2_add_79104_comb + p2_add_79105_comb;
  assign p2_add_79423_comb = p1_smul_76726 + p1_smul_76727;
  assign p2_add_79426_comb = p2_add_79106_comb + p2_add_79107_comb;
  assign p2_add_79427_comb = p1_smul_76732 + p1_smul_76733;
  assign p2_add_79430_comb = p2_add_79108_comb + p2_add_79109_comb;
  assign p2_add_79431_comb = p1_smul_76738 + p1_smul_76739;
  assign p2_add_79434_comb = p2_add_79110_comb + p2_add_79111_comb;
  assign p2_add_79435_comb = p1_smul_76744 + p1_smul_76745;
  assign p2_add_79438_comb = p2_add_79112_comb + p2_add_79113_comb;
  assign p2_add_79439_comb = p1_smul_76750 + p1_smul_76751;
  assign p2_add_79442_comb = p2_add_79114_comb + p2_add_79115_comb;
  assign p2_add_79443_comb = p1_smul_76756 + p1_smul_76757;
  assign p2_add_79446_comb = p2_add_79116_comb + p2_add_79117_comb;
  assign p2_add_79447_comb = p1_smul_76762 + p1_smul_76763;
  assign p2_add_79450_comb = p2_add_79118_comb + p2_add_79119_comb;
  assign p2_add_79451_comb = p1_smul_76768 + p1_smul_76769;
  assign p2_add_79454_comb = p2_add_79120_comb + p2_add_79121_comb;
  assign p2_add_79455_comb = p1_smul_76774 + p1_smul_76775;
  assign p2_add_79458_comb = p2_add_79122_comb + p2_add_79123_comb;
  assign p2_add_79459_comb = p1_smul_76780 + p1_smul_76781;
  assign p2_add_79462_comb = p2_add_79124_comb + p2_add_79125_comb;
  assign p2_add_79463_comb = p1_smul_76786 + p1_smul_76787;
  assign p2_add_79466_comb = p2_add_79126_comb + p2_add_79127_comb;
  assign p2_add_79467_comb = p1_smul_76792 + p1_smul_76793;
  assign p2_add_79470_comb = p2_add_79128_comb + p2_add_79129_comb;
  assign p2_add_79471_comb = p1_smul_76798 + p1_smul_76799;
  assign p2_add_79474_comb = p2_add_79130_comb + p2_add_79131_comb;
  assign p2_add_79475_comb = p1_smul_76804 + p1_smul_76805;
  assign p2_add_79478_comb = p2_add_79132_comb + p2_add_79133_comb;
  assign p2_add_79479_comb = p1_smul_76810 + p1_smul_76811;
  assign p2_add_79482_comb = p2_add_79134_comb + p2_add_79135_comb;
  assign p2_add_79483_comb = p1_smul_76816 + p1_smul_76817;
  assign p2_add_79486_comb = p2_add_79136_comb + p2_add_79137_comb;
  assign p2_add_79487_comb = p1_smul_76822 + p1_smul_76823;
  assign p2_add_79490_comb = p2_add_79138_comb + p2_add_79139_comb;
  assign p2_add_79491_comb = p1_smul_76828 + p1_smul_76829;
  assign p2_add_79494_comb = p2_add_79140_comb + p2_add_79141_comb;
  assign p2_add_79495_comb = p1_smul_76834 + p1_smul_76835;
  assign p2_add_79498_comb = p2_add_79142_comb + p2_add_79143_comb;
  assign p2_add_79499_comb = p1_smul_76840 + p1_smul_76841;
  assign p2_add_79502_comb = p2_add_79144_comb + p2_add_79145_comb;
  assign p2_add_79503_comb = p1_smul_76846 + p1_smul_76847;
  assign p2_add_79506_comb = p2_add_79146_comb + p2_add_79147_comb;
  assign p2_add_79507_comb = p1_smul_76852 + p1_smul_76853;
  assign p2_add_79510_comb = p2_add_79148_comb + p2_add_79149_comb;
  assign p2_add_79511_comb = p1_smul_76858 + p1_smul_76859;
  assign p2_add_79514_comb = p2_add_79150_comb + p2_add_79151_comb;
  assign p2_add_79515_comb = p1_smul_76864 + p1_smul_76865;
  assign p2_add_79518_comb = p2_add_79152_comb + p2_add_79153_comb;
  assign p2_add_79519_comb = p1_smul_76870 + p1_smul_76871;
  assign p2_add_79522_comb = p2_add_79154_comb + p2_add_79155_comb;
  assign p2_add_79523_comb = p1_smul_76876 + p1_smul_76877;
  assign p2_add_79526_comb = p2_add_79156_comb + p2_add_79157_comb;
  assign p2_add_79527_comb = p1_smul_76882 + p1_smul_76883;
  assign p2_add_79530_comb = p2_add_79158_comb + p2_add_79159_comb;
  assign p2_add_79531_comb = p1_smul_76888 + p1_smul_76889;
  assign p2_add_79534_comb = p2_add_79160_comb + p2_add_79161_comb;
  assign p2_add_79535_comb = p1_smul_76894 + p1_smul_76895;
  assign p2_add_79538_comb = p2_add_79162_comb + p2_add_79163_comb;
  assign p2_add_79539_comb = p1_smul_76900 + p1_smul_76901;
  assign p2_add_79542_comb = p2_add_79164_comb + p2_add_79165_comb;
  assign p2_add_79543_comb = p1_smul_76906 + p1_smul_76907;
  assign p2_add_79546_comb = p2_add_79166_comb + p2_add_79167_comb;
  assign p2_add_79547_comb = p1_smul_76912 + p1_smul_76913;
  assign p2_add_79550_comb = p2_add_79168_comb + p2_add_79169_comb;
  assign p2_add_79551_comb = p1_smul_76918 + p1_smul_76919;
  assign p2_add_79554_comb = p2_add_79170_comb + p2_add_79171_comb;
  assign p2_add_79555_comb = p1_smul_76924 + p1_smul_76925;
  assign p2_add_79558_comb = p2_add_79172_comb + p2_add_79173_comb;
  assign p2_add_79559_comb = p1_smul_76930 + p1_smul_76931;
  assign p2_add_79562_comb = p2_add_79174_comb + p2_add_79175_comb;
  assign p2_add_79563_comb = p1_smul_76936 + p1_smul_76937;
  assign p2_add_79566_comb = p2_add_79176_comb + p2_add_79177_comb;
  assign p2_add_79567_comb = p1_smul_76942 + p1_smul_76943;
  assign p2_add_79570_comb = p2_add_79178_comb + p2_add_79179_comb;
  assign p2_add_79571_comb = p1_smul_76948 + p1_smul_76949;
  assign p2_add_79574_comb = p2_add_79180_comb + p2_add_79181_comb;
  assign p2_add_79575_comb = p1_smul_76954 + p1_smul_76955;
  assign p2_add_79578_comb = p2_add_79182_comb + p2_add_79183_comb;
  assign p2_add_79579_comb = p1_smul_76960 + p1_smul_76961;
  assign p2_add_79582_comb = p2_add_79184_comb + p2_add_79185_comb;
  assign p2_add_79583_comb = p1_smul_76966 + p1_smul_76967;
  assign p2_add_79586_comb = p2_add_79188_comb + p2_add_79189_comb;
  assign p2_add_79587_comb = p2_add_79192_comb + p2_add_79193_comb;
  assign p2_add_79588_comb = p2_add_79196_comb + p2_add_79197_comb;
  assign p2_add_79589_comb = p2_add_79200_comb + p2_add_79201_comb;
  assign p2_add_79590_comb = p2_add_79204_comb + p2_add_79205_comb;
  assign p2_add_79591_comb = p2_add_79208_comb + p2_add_79209_comb;
  assign p2_add_79592_comb = p2_add_79212_comb + p2_add_79213_comb;
  assign p2_add_79593_comb = p2_add_79216_comb + p2_add_79217_comb;
  assign p2_add_79594_comb = p2_add_79220_comb + p2_add_79221_comb;
  assign p2_add_79595_comb = p2_add_79224_comb + p2_add_79225_comb;
  assign p2_add_79596_comb = p2_add_79228_comb + p2_add_79229_comb;
  assign p2_add_79597_comb = p2_add_79232_comb + p2_add_79233_comb;
  assign p2_add_79598_comb = p2_add_79236_comb + p2_add_79237_comb;
  assign p2_add_79599_comb = p2_add_79240_comb + p2_add_79241_comb;
  assign p2_add_79600_comb = p2_add_79244_comb + p2_add_79245_comb;
  assign p2_add_79601_comb = p2_add_79248_comb + p2_add_79249_comb;
  assign p2_add_79602_comb = p2_add_79252_comb + p2_add_79253_comb;
  assign p2_add_79603_comb = p2_add_79256_comb + p2_add_79257_comb;
  assign p2_add_79604_comb = p2_add_79260_comb + p2_add_79261_comb;
  assign p2_add_79605_comb = p2_add_79264_comb + p2_add_79265_comb;
  assign p2_add_79606_comb = p2_add_79268_comb + p2_add_79269_comb;
  assign p2_add_79607_comb = p2_add_79272_comb + p2_add_79273_comb;
  assign p2_add_79608_comb = p2_add_79276_comb + p2_add_79277_comb;
  assign p2_add_79609_comb = p2_add_79280_comb + p2_add_79281_comb;
  assign p2_add_79610_comb = p2_add_79284_comb + p2_add_79285_comb;
  assign p2_add_79611_comb = p2_add_79288_comb + p2_add_79289_comb;
  assign p2_add_79612_comb = p2_add_79292_comb + p2_add_79293_comb;
  assign p2_add_79613_comb = p2_add_79296_comb + p2_add_79297_comb;
  assign p2_add_79614_comb = p2_add_79300_comb + p2_add_79301_comb;
  assign p2_add_79615_comb = p2_add_79304_comb + p2_add_79305_comb;
  assign p2_add_79616_comb = p2_add_79308_comb + p2_add_79309_comb;
  assign p2_add_79617_comb = p2_add_79312_comb + p2_add_79313_comb;
  assign p2_add_79618_comb = p2_add_79316_comb + p2_add_79317_comb;
  assign p2_add_79619_comb = p2_add_79320_comb + p2_add_79321_comb;
  assign p2_add_79620_comb = p2_add_79324_comb + p2_add_79325_comb;
  assign p2_add_79621_comb = p2_add_79328_comb + p2_add_79329_comb;
  assign p2_add_79622_comb = p2_add_79332_comb + p2_add_79333_comb;
  assign p2_add_79623_comb = p2_add_79336_comb + p2_add_79337_comb;
  assign p2_add_79624_comb = p2_add_79340_comb + p2_add_79341_comb;
  assign p2_add_79625_comb = p2_add_79344_comb + p2_add_79345_comb;
  assign p2_add_79626_comb = p2_add_79348_comb + p2_add_79349_comb;
  assign p2_add_79627_comb = p2_add_79352_comb + p2_add_79353_comb;
  assign p2_add_79628_comb = p2_add_79356_comb + p2_add_79357_comb;
  assign p2_add_79629_comb = p2_add_79360_comb + p2_add_79361_comb;
  assign p2_add_79630_comb = p2_add_79364_comb + p2_add_79365_comb;
  assign p2_add_79631_comb = p2_add_79368_comb + p2_add_79369_comb;
  assign p2_add_79632_comb = p2_add_79372_comb + p2_add_79373_comb;
  assign p2_add_79633_comb = p2_add_79376_comb + p2_add_79377_comb;
  assign p2_add_79634_comb = p2_add_79380_comb + p2_add_79381_comb;
  assign p2_add_79635_comb = p2_add_79384_comb + p2_add_79385_comb;
  assign p2_add_79636_comb = p2_add_79388_comb + p2_add_79389_comb;
  assign p2_add_79637_comb = p2_add_79392_comb + p2_add_79393_comb;
  assign p2_add_79638_comb = p2_add_79396_comb + p2_add_79397_comb;
  assign p2_add_79639_comb = p2_add_79400_comb + p2_add_79401_comb;
  assign p2_add_79640_comb = p2_add_79404_comb + p2_add_79405_comb;
  assign p2_add_79641_comb = p2_add_79408_comb + p2_add_79409_comb;
  assign p2_add_79642_comb = p2_add_79412_comb + p2_add_79413_comb;
  assign p2_add_79643_comb = p2_add_79416_comb + p2_add_79417_comb;
  assign p2_add_79644_comb = p2_add_79420_comb + p2_add_79421_comb;
  assign p2_add_79645_comb = p2_add_79424_comb + p2_add_79425_comb;
  assign p2_add_79646_comb = p2_add_79428_comb + p2_add_79429_comb;
  assign p2_add_79647_comb = p2_add_79432_comb + p2_add_79433_comb;
  assign p2_add_79648_comb = p2_add_79436_comb + p2_add_79437_comb;
  assign p2_add_79649_comb = p2_add_79440_comb + p2_add_79441_comb;
  assign p2_add_79650_comb = p2_add_79444_comb + p2_add_79445_comb;
  assign p2_add_79651_comb = p2_add_79448_comb + p2_add_79449_comb;
  assign p2_add_79652_comb = p2_add_79452_comb + p2_add_79453_comb;
  assign p2_add_79653_comb = p2_add_79456_comb + p2_add_79457_comb;
  assign p2_add_79654_comb = p2_add_79460_comb + p2_add_79461_comb;
  assign p2_add_79655_comb = p2_add_79464_comb + p2_add_79465_comb;
  assign p2_add_79656_comb = p2_add_79468_comb + p2_add_79469_comb;
  assign p2_add_79657_comb = p2_add_79472_comb + p2_add_79473_comb;
  assign p2_add_79658_comb = p2_add_79476_comb + p2_add_79477_comb;
  assign p2_add_79659_comb = p2_add_79480_comb + p2_add_79481_comb;
  assign p2_add_79660_comb = p2_add_79484_comb + p2_add_79485_comb;
  assign p2_add_79661_comb = p2_add_79488_comb + p2_add_79489_comb;
  assign p2_add_79662_comb = p2_add_79492_comb + p2_add_79493_comb;
  assign p2_add_79663_comb = p2_add_79496_comb + p2_add_79497_comb;
  assign p2_add_79664_comb = p2_add_79500_comb + p2_add_79501_comb;
  assign p2_add_79665_comb = p2_add_79504_comb + p2_add_79505_comb;
  assign p2_add_79666_comb = p2_add_79508_comb + p2_add_79509_comb;
  assign p2_add_79667_comb = p2_add_79512_comb + p2_add_79513_comb;
  assign p2_add_79668_comb = p2_add_79516_comb + p2_add_79517_comb;
  assign p2_add_79669_comb = p2_add_79520_comb + p2_add_79521_comb;
  assign p2_add_79670_comb = p2_add_79524_comb + p2_add_79525_comb;
  assign p2_add_79671_comb = p2_add_79528_comb + p2_add_79529_comb;
  assign p2_add_79672_comb = p2_add_79532_comb + p2_add_79533_comb;
  assign p2_add_79673_comb = p2_add_79536_comb + p2_add_79537_comb;
  assign p2_add_79674_comb = p2_add_79540_comb + p2_add_79541_comb;
  assign p2_add_79675_comb = p2_add_79544_comb + p2_add_79545_comb;
  assign p2_add_79676_comb = p2_add_79548_comb + p2_add_79549_comb;
  assign p2_add_79677_comb = p2_add_79552_comb + p2_add_79553_comb;
  assign p2_add_79678_comb = p2_add_79556_comb + p2_add_79557_comb;
  assign p2_add_79679_comb = p2_add_79560_comb + p2_add_79561_comb;
  assign p2_add_79680_comb = p2_add_79564_comb + p2_add_79565_comb;
  assign p2_add_79681_comb = p2_add_79568_comb + p2_add_79569_comb;
  assign p2_add_79682_comb = p2_add_79572_comb + p2_add_79573_comb;
  assign p2_add_79683_comb = p2_add_79576_comb + p2_add_79577_comb;
  assign p2_add_79684_comb = p2_add_79580_comb + p2_add_79581_comb;
  assign p2_add_79685_comb = p2_add_79584_comb + p2_add_79585_comb;

  // Registers for pipe stage 2:
  reg [31:0] p2_add_79186;
  reg [31:0] p2_add_79187;
  reg [31:0] p2_add_79190;
  reg [31:0] p2_add_79191;
  reg [31:0] p2_add_79194;
  reg [31:0] p2_add_79195;
  reg [31:0] p2_add_79198;
  reg [31:0] p2_add_79199;
  reg [31:0] p2_add_79202;
  reg [31:0] p2_add_79203;
  reg [31:0] p2_add_79206;
  reg [31:0] p2_add_79207;
  reg [31:0] p2_add_79210;
  reg [31:0] p2_add_79211;
  reg [31:0] p2_add_79214;
  reg [31:0] p2_add_79215;
  reg [31:0] p2_add_79218;
  reg [31:0] p2_add_79219;
  reg [31:0] p2_add_79222;
  reg [31:0] p2_add_79223;
  reg [31:0] p2_add_79226;
  reg [31:0] p2_add_79227;
  reg [31:0] p2_add_79230;
  reg [31:0] p2_add_79231;
  reg [31:0] p2_add_79234;
  reg [31:0] p2_add_79235;
  reg [31:0] p2_add_79238;
  reg [31:0] p2_add_79239;
  reg [31:0] p2_add_79242;
  reg [31:0] p2_add_79243;
  reg [31:0] p2_add_79246;
  reg [31:0] p2_add_79247;
  reg [31:0] p2_add_79250;
  reg [31:0] p2_add_79251;
  reg [31:0] p2_add_79254;
  reg [31:0] p2_add_79255;
  reg [31:0] p2_add_79258;
  reg [31:0] p2_add_79259;
  reg [31:0] p2_add_79262;
  reg [31:0] p2_add_79263;
  reg [31:0] p2_add_79266;
  reg [31:0] p2_add_79267;
  reg [31:0] p2_add_79270;
  reg [31:0] p2_add_79271;
  reg [31:0] p2_add_79274;
  reg [31:0] p2_add_79275;
  reg [31:0] p2_add_79278;
  reg [31:0] p2_add_79279;
  reg [31:0] p2_add_79282;
  reg [31:0] p2_add_79283;
  reg [31:0] p2_add_79286;
  reg [31:0] p2_add_79287;
  reg [31:0] p2_add_79290;
  reg [31:0] p2_add_79291;
  reg [31:0] p2_add_79294;
  reg [31:0] p2_add_79295;
  reg [31:0] p2_add_79298;
  reg [31:0] p2_add_79299;
  reg [31:0] p2_add_79302;
  reg [31:0] p2_add_79303;
  reg [31:0] p2_add_79306;
  reg [31:0] p2_add_79307;
  reg [31:0] p2_add_79310;
  reg [31:0] p2_add_79311;
  reg [31:0] p2_add_79314;
  reg [31:0] p2_add_79315;
  reg [31:0] p2_add_79318;
  reg [31:0] p2_add_79319;
  reg [31:0] p2_add_79322;
  reg [31:0] p2_add_79323;
  reg [31:0] p2_add_79326;
  reg [31:0] p2_add_79327;
  reg [31:0] p2_add_79330;
  reg [31:0] p2_add_79331;
  reg [31:0] p2_add_79334;
  reg [31:0] p2_add_79335;
  reg [31:0] p2_add_79338;
  reg [31:0] p2_add_79339;
  reg [31:0] p2_add_79342;
  reg [31:0] p2_add_79343;
  reg [31:0] p2_add_79346;
  reg [31:0] p2_add_79347;
  reg [31:0] p2_add_79350;
  reg [31:0] p2_add_79351;
  reg [31:0] p2_add_79354;
  reg [31:0] p2_add_79355;
  reg [31:0] p2_add_79358;
  reg [31:0] p2_add_79359;
  reg [31:0] p2_add_79362;
  reg [31:0] p2_add_79363;
  reg [31:0] p2_add_79366;
  reg [31:0] p2_add_79367;
  reg [31:0] p2_add_79370;
  reg [31:0] p2_add_79371;
  reg [31:0] p2_add_79374;
  reg [31:0] p2_add_79375;
  reg [31:0] p2_add_79378;
  reg [31:0] p2_add_79379;
  reg [31:0] p2_add_79382;
  reg [31:0] p2_add_79383;
  reg [31:0] p2_add_79386;
  reg [31:0] p2_add_79387;
  reg [31:0] p2_add_79390;
  reg [31:0] p2_add_79391;
  reg [31:0] p2_add_79394;
  reg [31:0] p2_add_79395;
  reg [31:0] p2_add_79398;
  reg [31:0] p2_add_79399;
  reg [31:0] p2_add_79402;
  reg [31:0] p2_add_79403;
  reg [31:0] p2_add_79406;
  reg [31:0] p2_add_79407;
  reg [31:0] p2_add_79410;
  reg [31:0] p2_add_79411;
  reg [31:0] p2_add_79414;
  reg [31:0] p2_add_79415;
  reg [31:0] p2_add_79418;
  reg [31:0] p2_add_79419;
  reg [31:0] p2_add_79422;
  reg [31:0] p2_add_79423;
  reg [31:0] p2_add_79426;
  reg [31:0] p2_add_79427;
  reg [31:0] p2_add_79430;
  reg [31:0] p2_add_79431;
  reg [31:0] p2_add_79434;
  reg [31:0] p2_add_79435;
  reg [31:0] p2_add_79438;
  reg [31:0] p2_add_79439;
  reg [31:0] p2_add_79442;
  reg [31:0] p2_add_79443;
  reg [31:0] p2_add_79446;
  reg [31:0] p2_add_79447;
  reg [31:0] p2_add_79450;
  reg [31:0] p2_add_79451;
  reg [31:0] p2_add_79454;
  reg [31:0] p2_add_79455;
  reg [31:0] p2_add_79458;
  reg [31:0] p2_add_79459;
  reg [31:0] p2_add_79462;
  reg [31:0] p2_add_79463;
  reg [31:0] p2_add_79466;
  reg [31:0] p2_add_79467;
  reg [31:0] p2_add_79470;
  reg [31:0] p2_add_79471;
  reg [31:0] p2_add_79474;
  reg [31:0] p2_add_79475;
  reg [31:0] p2_add_79478;
  reg [31:0] p2_add_79479;
  reg [31:0] p2_add_79482;
  reg [31:0] p2_add_79483;
  reg [31:0] p2_add_79486;
  reg [31:0] p2_add_79487;
  reg [31:0] p2_add_79490;
  reg [31:0] p2_add_79491;
  reg [31:0] p2_add_79494;
  reg [31:0] p2_add_79495;
  reg [31:0] p2_add_79498;
  reg [31:0] p2_add_79499;
  reg [31:0] p2_add_79502;
  reg [31:0] p2_add_79503;
  reg [31:0] p2_add_79506;
  reg [31:0] p2_add_79507;
  reg [31:0] p2_add_79510;
  reg [31:0] p2_add_79511;
  reg [31:0] p2_add_79514;
  reg [31:0] p2_add_79515;
  reg [31:0] p2_add_79518;
  reg [31:0] p2_add_79519;
  reg [31:0] p2_add_79522;
  reg [31:0] p2_add_79523;
  reg [31:0] p2_add_79526;
  reg [31:0] p2_add_79527;
  reg [31:0] p2_add_79530;
  reg [31:0] p2_add_79531;
  reg [31:0] p2_add_79534;
  reg [31:0] p2_add_79535;
  reg [31:0] p2_add_79538;
  reg [31:0] p2_add_79539;
  reg [31:0] p2_add_79542;
  reg [31:0] p2_add_79543;
  reg [31:0] p2_add_79546;
  reg [31:0] p2_add_79547;
  reg [31:0] p2_add_79550;
  reg [31:0] p2_add_79551;
  reg [31:0] p2_add_79554;
  reg [31:0] p2_add_79555;
  reg [31:0] p2_add_79558;
  reg [31:0] p2_add_79559;
  reg [31:0] p2_add_79562;
  reg [31:0] p2_add_79563;
  reg [31:0] p2_add_79566;
  reg [31:0] p2_add_79567;
  reg [31:0] p2_add_79570;
  reg [31:0] p2_add_79571;
  reg [31:0] p2_add_79574;
  reg [31:0] p2_add_79575;
  reg [31:0] p2_add_79578;
  reg [31:0] p2_add_79579;
  reg [31:0] p2_add_79582;
  reg [31:0] p2_add_79583;
  reg [31:0] p2_add_79586;
  reg [31:0] p2_add_79587;
  reg [31:0] p2_add_79588;
  reg [31:0] p2_add_79589;
  reg [31:0] p2_add_79590;
  reg [31:0] p2_add_79591;
  reg [31:0] p2_add_79592;
  reg [31:0] p2_add_79593;
  reg [31:0] p2_add_79594;
  reg [31:0] p2_add_79595;
  reg [31:0] p2_add_79596;
  reg [31:0] p2_add_79597;
  reg [31:0] p2_add_79598;
  reg [31:0] p2_add_79599;
  reg [31:0] p2_add_79600;
  reg [31:0] p2_add_79601;
  reg [31:0] p2_add_79602;
  reg [31:0] p2_add_79603;
  reg [31:0] p2_add_79604;
  reg [31:0] p2_add_79605;
  reg [31:0] p2_add_79606;
  reg [31:0] p2_add_79607;
  reg [31:0] p2_add_79608;
  reg [31:0] p2_add_79609;
  reg [31:0] p2_add_79610;
  reg [31:0] p2_add_79611;
  reg [31:0] p2_add_79612;
  reg [31:0] p2_add_79613;
  reg [31:0] p2_add_79614;
  reg [31:0] p2_add_79615;
  reg [31:0] p2_add_79616;
  reg [31:0] p2_add_79617;
  reg [31:0] p2_add_79618;
  reg [31:0] p2_add_79619;
  reg [31:0] p2_add_79620;
  reg [31:0] p2_add_79621;
  reg [31:0] p2_add_79622;
  reg [31:0] p2_add_79623;
  reg [31:0] p2_add_79624;
  reg [31:0] p2_add_79625;
  reg [31:0] p2_add_79626;
  reg [31:0] p2_add_79627;
  reg [31:0] p2_add_79628;
  reg [31:0] p2_add_79629;
  reg [31:0] p2_add_79630;
  reg [31:0] p2_add_79631;
  reg [31:0] p2_add_79632;
  reg [31:0] p2_add_79633;
  reg [31:0] p2_add_79634;
  reg [31:0] p2_add_79635;
  reg [31:0] p2_add_79636;
  reg [31:0] p2_add_79637;
  reg [31:0] p2_add_79638;
  reg [31:0] p2_add_79639;
  reg [31:0] p2_add_79640;
  reg [31:0] p2_add_79641;
  reg [31:0] p2_add_79642;
  reg [31:0] p2_add_79643;
  reg [31:0] p2_add_79644;
  reg [31:0] p2_add_79645;
  reg [31:0] p2_add_79646;
  reg [31:0] p2_add_79647;
  reg [31:0] p2_add_79648;
  reg [31:0] p2_add_79649;
  reg [31:0] p2_add_79650;
  reg [31:0] p2_add_79651;
  reg [31:0] p2_add_79652;
  reg [31:0] p2_add_79653;
  reg [31:0] p2_add_79654;
  reg [31:0] p2_add_79655;
  reg [31:0] p2_add_79656;
  reg [31:0] p2_add_79657;
  reg [31:0] p2_add_79658;
  reg [31:0] p2_add_79659;
  reg [31:0] p2_add_79660;
  reg [31:0] p2_add_79661;
  reg [31:0] p2_add_79662;
  reg [31:0] p2_add_79663;
  reg [31:0] p2_add_79664;
  reg [31:0] p2_add_79665;
  reg [31:0] p2_add_79666;
  reg [31:0] p2_add_79667;
  reg [31:0] p2_add_79668;
  reg [31:0] p2_add_79669;
  reg [31:0] p2_add_79670;
  reg [31:0] p2_add_79671;
  reg [31:0] p2_add_79672;
  reg [31:0] p2_add_79673;
  reg [31:0] p2_add_79674;
  reg [31:0] p2_add_79675;
  reg [31:0] p2_add_79676;
  reg [31:0] p2_add_79677;
  reg [31:0] p2_add_79678;
  reg [31:0] p2_add_79679;
  reg [31:0] p2_add_79680;
  reg [31:0] p2_add_79681;
  reg [31:0] p2_add_79682;
  reg [31:0] p2_add_79683;
  reg [31:0] p2_add_79684;
  reg [31:0] p2_add_79685;
  always_ff @ (posedge clk) begin
    p2_add_79186 <= p2_add_79186_comb;
    p2_add_79187 <= p2_add_79187_comb;
    p2_add_79190 <= p2_add_79190_comb;
    p2_add_79191 <= p2_add_79191_comb;
    p2_add_79194 <= p2_add_79194_comb;
    p2_add_79195 <= p2_add_79195_comb;
    p2_add_79198 <= p2_add_79198_comb;
    p2_add_79199 <= p2_add_79199_comb;
    p2_add_79202 <= p2_add_79202_comb;
    p2_add_79203 <= p2_add_79203_comb;
    p2_add_79206 <= p2_add_79206_comb;
    p2_add_79207 <= p2_add_79207_comb;
    p2_add_79210 <= p2_add_79210_comb;
    p2_add_79211 <= p2_add_79211_comb;
    p2_add_79214 <= p2_add_79214_comb;
    p2_add_79215 <= p2_add_79215_comb;
    p2_add_79218 <= p2_add_79218_comb;
    p2_add_79219 <= p2_add_79219_comb;
    p2_add_79222 <= p2_add_79222_comb;
    p2_add_79223 <= p2_add_79223_comb;
    p2_add_79226 <= p2_add_79226_comb;
    p2_add_79227 <= p2_add_79227_comb;
    p2_add_79230 <= p2_add_79230_comb;
    p2_add_79231 <= p2_add_79231_comb;
    p2_add_79234 <= p2_add_79234_comb;
    p2_add_79235 <= p2_add_79235_comb;
    p2_add_79238 <= p2_add_79238_comb;
    p2_add_79239 <= p2_add_79239_comb;
    p2_add_79242 <= p2_add_79242_comb;
    p2_add_79243 <= p2_add_79243_comb;
    p2_add_79246 <= p2_add_79246_comb;
    p2_add_79247 <= p2_add_79247_comb;
    p2_add_79250 <= p2_add_79250_comb;
    p2_add_79251 <= p2_add_79251_comb;
    p2_add_79254 <= p2_add_79254_comb;
    p2_add_79255 <= p2_add_79255_comb;
    p2_add_79258 <= p2_add_79258_comb;
    p2_add_79259 <= p2_add_79259_comb;
    p2_add_79262 <= p2_add_79262_comb;
    p2_add_79263 <= p2_add_79263_comb;
    p2_add_79266 <= p2_add_79266_comb;
    p2_add_79267 <= p2_add_79267_comb;
    p2_add_79270 <= p2_add_79270_comb;
    p2_add_79271 <= p2_add_79271_comb;
    p2_add_79274 <= p2_add_79274_comb;
    p2_add_79275 <= p2_add_79275_comb;
    p2_add_79278 <= p2_add_79278_comb;
    p2_add_79279 <= p2_add_79279_comb;
    p2_add_79282 <= p2_add_79282_comb;
    p2_add_79283 <= p2_add_79283_comb;
    p2_add_79286 <= p2_add_79286_comb;
    p2_add_79287 <= p2_add_79287_comb;
    p2_add_79290 <= p2_add_79290_comb;
    p2_add_79291 <= p2_add_79291_comb;
    p2_add_79294 <= p2_add_79294_comb;
    p2_add_79295 <= p2_add_79295_comb;
    p2_add_79298 <= p2_add_79298_comb;
    p2_add_79299 <= p2_add_79299_comb;
    p2_add_79302 <= p2_add_79302_comb;
    p2_add_79303 <= p2_add_79303_comb;
    p2_add_79306 <= p2_add_79306_comb;
    p2_add_79307 <= p2_add_79307_comb;
    p2_add_79310 <= p2_add_79310_comb;
    p2_add_79311 <= p2_add_79311_comb;
    p2_add_79314 <= p2_add_79314_comb;
    p2_add_79315 <= p2_add_79315_comb;
    p2_add_79318 <= p2_add_79318_comb;
    p2_add_79319 <= p2_add_79319_comb;
    p2_add_79322 <= p2_add_79322_comb;
    p2_add_79323 <= p2_add_79323_comb;
    p2_add_79326 <= p2_add_79326_comb;
    p2_add_79327 <= p2_add_79327_comb;
    p2_add_79330 <= p2_add_79330_comb;
    p2_add_79331 <= p2_add_79331_comb;
    p2_add_79334 <= p2_add_79334_comb;
    p2_add_79335 <= p2_add_79335_comb;
    p2_add_79338 <= p2_add_79338_comb;
    p2_add_79339 <= p2_add_79339_comb;
    p2_add_79342 <= p2_add_79342_comb;
    p2_add_79343 <= p2_add_79343_comb;
    p2_add_79346 <= p2_add_79346_comb;
    p2_add_79347 <= p2_add_79347_comb;
    p2_add_79350 <= p2_add_79350_comb;
    p2_add_79351 <= p2_add_79351_comb;
    p2_add_79354 <= p2_add_79354_comb;
    p2_add_79355 <= p2_add_79355_comb;
    p2_add_79358 <= p2_add_79358_comb;
    p2_add_79359 <= p2_add_79359_comb;
    p2_add_79362 <= p2_add_79362_comb;
    p2_add_79363 <= p2_add_79363_comb;
    p2_add_79366 <= p2_add_79366_comb;
    p2_add_79367 <= p2_add_79367_comb;
    p2_add_79370 <= p2_add_79370_comb;
    p2_add_79371 <= p2_add_79371_comb;
    p2_add_79374 <= p2_add_79374_comb;
    p2_add_79375 <= p2_add_79375_comb;
    p2_add_79378 <= p2_add_79378_comb;
    p2_add_79379 <= p2_add_79379_comb;
    p2_add_79382 <= p2_add_79382_comb;
    p2_add_79383 <= p2_add_79383_comb;
    p2_add_79386 <= p2_add_79386_comb;
    p2_add_79387 <= p2_add_79387_comb;
    p2_add_79390 <= p2_add_79390_comb;
    p2_add_79391 <= p2_add_79391_comb;
    p2_add_79394 <= p2_add_79394_comb;
    p2_add_79395 <= p2_add_79395_comb;
    p2_add_79398 <= p2_add_79398_comb;
    p2_add_79399 <= p2_add_79399_comb;
    p2_add_79402 <= p2_add_79402_comb;
    p2_add_79403 <= p2_add_79403_comb;
    p2_add_79406 <= p2_add_79406_comb;
    p2_add_79407 <= p2_add_79407_comb;
    p2_add_79410 <= p2_add_79410_comb;
    p2_add_79411 <= p2_add_79411_comb;
    p2_add_79414 <= p2_add_79414_comb;
    p2_add_79415 <= p2_add_79415_comb;
    p2_add_79418 <= p2_add_79418_comb;
    p2_add_79419 <= p2_add_79419_comb;
    p2_add_79422 <= p2_add_79422_comb;
    p2_add_79423 <= p2_add_79423_comb;
    p2_add_79426 <= p2_add_79426_comb;
    p2_add_79427 <= p2_add_79427_comb;
    p2_add_79430 <= p2_add_79430_comb;
    p2_add_79431 <= p2_add_79431_comb;
    p2_add_79434 <= p2_add_79434_comb;
    p2_add_79435 <= p2_add_79435_comb;
    p2_add_79438 <= p2_add_79438_comb;
    p2_add_79439 <= p2_add_79439_comb;
    p2_add_79442 <= p2_add_79442_comb;
    p2_add_79443 <= p2_add_79443_comb;
    p2_add_79446 <= p2_add_79446_comb;
    p2_add_79447 <= p2_add_79447_comb;
    p2_add_79450 <= p2_add_79450_comb;
    p2_add_79451 <= p2_add_79451_comb;
    p2_add_79454 <= p2_add_79454_comb;
    p2_add_79455 <= p2_add_79455_comb;
    p2_add_79458 <= p2_add_79458_comb;
    p2_add_79459 <= p2_add_79459_comb;
    p2_add_79462 <= p2_add_79462_comb;
    p2_add_79463 <= p2_add_79463_comb;
    p2_add_79466 <= p2_add_79466_comb;
    p2_add_79467 <= p2_add_79467_comb;
    p2_add_79470 <= p2_add_79470_comb;
    p2_add_79471 <= p2_add_79471_comb;
    p2_add_79474 <= p2_add_79474_comb;
    p2_add_79475 <= p2_add_79475_comb;
    p2_add_79478 <= p2_add_79478_comb;
    p2_add_79479 <= p2_add_79479_comb;
    p2_add_79482 <= p2_add_79482_comb;
    p2_add_79483 <= p2_add_79483_comb;
    p2_add_79486 <= p2_add_79486_comb;
    p2_add_79487 <= p2_add_79487_comb;
    p2_add_79490 <= p2_add_79490_comb;
    p2_add_79491 <= p2_add_79491_comb;
    p2_add_79494 <= p2_add_79494_comb;
    p2_add_79495 <= p2_add_79495_comb;
    p2_add_79498 <= p2_add_79498_comb;
    p2_add_79499 <= p2_add_79499_comb;
    p2_add_79502 <= p2_add_79502_comb;
    p2_add_79503 <= p2_add_79503_comb;
    p2_add_79506 <= p2_add_79506_comb;
    p2_add_79507 <= p2_add_79507_comb;
    p2_add_79510 <= p2_add_79510_comb;
    p2_add_79511 <= p2_add_79511_comb;
    p2_add_79514 <= p2_add_79514_comb;
    p2_add_79515 <= p2_add_79515_comb;
    p2_add_79518 <= p2_add_79518_comb;
    p2_add_79519 <= p2_add_79519_comb;
    p2_add_79522 <= p2_add_79522_comb;
    p2_add_79523 <= p2_add_79523_comb;
    p2_add_79526 <= p2_add_79526_comb;
    p2_add_79527 <= p2_add_79527_comb;
    p2_add_79530 <= p2_add_79530_comb;
    p2_add_79531 <= p2_add_79531_comb;
    p2_add_79534 <= p2_add_79534_comb;
    p2_add_79535 <= p2_add_79535_comb;
    p2_add_79538 <= p2_add_79538_comb;
    p2_add_79539 <= p2_add_79539_comb;
    p2_add_79542 <= p2_add_79542_comb;
    p2_add_79543 <= p2_add_79543_comb;
    p2_add_79546 <= p2_add_79546_comb;
    p2_add_79547 <= p2_add_79547_comb;
    p2_add_79550 <= p2_add_79550_comb;
    p2_add_79551 <= p2_add_79551_comb;
    p2_add_79554 <= p2_add_79554_comb;
    p2_add_79555 <= p2_add_79555_comb;
    p2_add_79558 <= p2_add_79558_comb;
    p2_add_79559 <= p2_add_79559_comb;
    p2_add_79562 <= p2_add_79562_comb;
    p2_add_79563 <= p2_add_79563_comb;
    p2_add_79566 <= p2_add_79566_comb;
    p2_add_79567 <= p2_add_79567_comb;
    p2_add_79570 <= p2_add_79570_comb;
    p2_add_79571 <= p2_add_79571_comb;
    p2_add_79574 <= p2_add_79574_comb;
    p2_add_79575 <= p2_add_79575_comb;
    p2_add_79578 <= p2_add_79578_comb;
    p2_add_79579 <= p2_add_79579_comb;
    p2_add_79582 <= p2_add_79582_comb;
    p2_add_79583 <= p2_add_79583_comb;
    p2_add_79586 <= p2_add_79586_comb;
    p2_add_79587 <= p2_add_79587_comb;
    p2_add_79588 <= p2_add_79588_comb;
    p2_add_79589 <= p2_add_79589_comb;
    p2_add_79590 <= p2_add_79590_comb;
    p2_add_79591 <= p2_add_79591_comb;
    p2_add_79592 <= p2_add_79592_comb;
    p2_add_79593 <= p2_add_79593_comb;
    p2_add_79594 <= p2_add_79594_comb;
    p2_add_79595 <= p2_add_79595_comb;
    p2_add_79596 <= p2_add_79596_comb;
    p2_add_79597 <= p2_add_79597_comb;
    p2_add_79598 <= p2_add_79598_comb;
    p2_add_79599 <= p2_add_79599_comb;
    p2_add_79600 <= p2_add_79600_comb;
    p2_add_79601 <= p2_add_79601_comb;
    p2_add_79602 <= p2_add_79602_comb;
    p2_add_79603 <= p2_add_79603_comb;
    p2_add_79604 <= p2_add_79604_comb;
    p2_add_79605 <= p2_add_79605_comb;
    p2_add_79606 <= p2_add_79606_comb;
    p2_add_79607 <= p2_add_79607_comb;
    p2_add_79608 <= p2_add_79608_comb;
    p2_add_79609 <= p2_add_79609_comb;
    p2_add_79610 <= p2_add_79610_comb;
    p2_add_79611 <= p2_add_79611_comb;
    p2_add_79612 <= p2_add_79612_comb;
    p2_add_79613 <= p2_add_79613_comb;
    p2_add_79614 <= p2_add_79614_comb;
    p2_add_79615 <= p2_add_79615_comb;
    p2_add_79616 <= p2_add_79616_comb;
    p2_add_79617 <= p2_add_79617_comb;
    p2_add_79618 <= p2_add_79618_comb;
    p2_add_79619 <= p2_add_79619_comb;
    p2_add_79620 <= p2_add_79620_comb;
    p2_add_79621 <= p2_add_79621_comb;
    p2_add_79622 <= p2_add_79622_comb;
    p2_add_79623 <= p2_add_79623_comb;
    p2_add_79624 <= p2_add_79624_comb;
    p2_add_79625 <= p2_add_79625_comb;
    p2_add_79626 <= p2_add_79626_comb;
    p2_add_79627 <= p2_add_79627_comb;
    p2_add_79628 <= p2_add_79628_comb;
    p2_add_79629 <= p2_add_79629_comb;
    p2_add_79630 <= p2_add_79630_comb;
    p2_add_79631 <= p2_add_79631_comb;
    p2_add_79632 <= p2_add_79632_comb;
    p2_add_79633 <= p2_add_79633_comb;
    p2_add_79634 <= p2_add_79634_comb;
    p2_add_79635 <= p2_add_79635_comb;
    p2_add_79636 <= p2_add_79636_comb;
    p2_add_79637 <= p2_add_79637_comb;
    p2_add_79638 <= p2_add_79638_comb;
    p2_add_79639 <= p2_add_79639_comb;
    p2_add_79640 <= p2_add_79640_comb;
    p2_add_79641 <= p2_add_79641_comb;
    p2_add_79642 <= p2_add_79642_comb;
    p2_add_79643 <= p2_add_79643_comb;
    p2_add_79644 <= p2_add_79644_comb;
    p2_add_79645 <= p2_add_79645_comb;
    p2_add_79646 <= p2_add_79646_comb;
    p2_add_79647 <= p2_add_79647_comb;
    p2_add_79648 <= p2_add_79648_comb;
    p2_add_79649 <= p2_add_79649_comb;
    p2_add_79650 <= p2_add_79650_comb;
    p2_add_79651 <= p2_add_79651_comb;
    p2_add_79652 <= p2_add_79652_comb;
    p2_add_79653 <= p2_add_79653_comb;
    p2_add_79654 <= p2_add_79654_comb;
    p2_add_79655 <= p2_add_79655_comb;
    p2_add_79656 <= p2_add_79656_comb;
    p2_add_79657 <= p2_add_79657_comb;
    p2_add_79658 <= p2_add_79658_comb;
    p2_add_79659 <= p2_add_79659_comb;
    p2_add_79660 <= p2_add_79660_comb;
    p2_add_79661 <= p2_add_79661_comb;
    p2_add_79662 <= p2_add_79662_comb;
    p2_add_79663 <= p2_add_79663_comb;
    p2_add_79664 <= p2_add_79664_comb;
    p2_add_79665 <= p2_add_79665_comb;
    p2_add_79666 <= p2_add_79666_comb;
    p2_add_79667 <= p2_add_79667_comb;
    p2_add_79668 <= p2_add_79668_comb;
    p2_add_79669 <= p2_add_79669_comb;
    p2_add_79670 <= p2_add_79670_comb;
    p2_add_79671 <= p2_add_79671_comb;
    p2_add_79672 <= p2_add_79672_comb;
    p2_add_79673 <= p2_add_79673_comb;
    p2_add_79674 <= p2_add_79674_comb;
    p2_add_79675 <= p2_add_79675_comb;
    p2_add_79676 <= p2_add_79676_comb;
    p2_add_79677 <= p2_add_79677_comb;
    p2_add_79678 <= p2_add_79678_comb;
    p2_add_79679 <= p2_add_79679_comb;
    p2_add_79680 <= p2_add_79680_comb;
    p2_add_79681 <= p2_add_79681_comb;
    p2_add_79682 <= p2_add_79682_comb;
    p2_add_79683 <= p2_add_79683_comb;
    p2_add_79684 <= p2_add_79684_comb;
    p2_add_79685 <= p2_add_79685_comb;
  end

  // ===== Pipe stage 3:
  wire [31:0] p3_add_80299_comb;
  wire [31:0] p3_add_80300_comb;
  wire [31:0] p3_add_80301_comb;
  wire [31:0] p3_add_80302_comb;
  wire [31:0] p3_add_80303_comb;
  wire [31:0] p3_add_80304_comb;
  wire [31:0] p3_add_80305_comb;
  wire [31:0] p3_add_80306_comb;
  wire [31:0] p3_add_80307_comb;
  wire [31:0] p3_add_80308_comb;
  wire [31:0] p3_add_80309_comb;
  wire [31:0] p3_add_80310_comb;
  wire [31:0] p3_add_80311_comb;
  wire [31:0] p3_add_80312_comb;
  wire [31:0] p3_add_80313_comb;
  wire [31:0] p3_add_80314_comb;
  wire [31:0] p3_add_80315_comb;
  wire [31:0] p3_add_80316_comb;
  wire [31:0] p3_add_80317_comb;
  wire [31:0] p3_add_80318_comb;
  wire [31:0] p3_add_80319_comb;
  wire [31:0] p3_add_80320_comb;
  wire [31:0] p3_add_80321_comb;
  wire [31:0] p3_add_80322_comb;
  wire [31:0] p3_add_80323_comb;
  wire [31:0] p3_add_80324_comb;
  wire [31:0] p3_add_80325_comb;
  wire [31:0] p3_add_80326_comb;
  wire [31:0] p3_add_80327_comb;
  wire [31:0] p3_add_80328_comb;
  wire [31:0] p3_add_80329_comb;
  wire [31:0] p3_add_80330_comb;
  wire [31:0] p3_add_80331_comb;
  wire [31:0] p3_add_80332_comb;
  wire [31:0] p3_add_80333_comb;
  wire [31:0] p3_add_80334_comb;
  wire [31:0] p3_add_80335_comb;
  wire [31:0] p3_add_80336_comb;
  wire [31:0] p3_add_80337_comb;
  wire [31:0] p3_add_80338_comb;
  wire [31:0] p3_add_80339_comb;
  wire [31:0] p3_add_80340_comb;
  wire [31:0] p3_add_80341_comb;
  wire [31:0] p3_add_80342_comb;
  wire [31:0] p3_add_80343_comb;
  wire [31:0] p3_add_80344_comb;
  wire [31:0] p3_add_80345_comb;
  wire [31:0] p3_add_80346_comb;
  wire [31:0] p3_add_80347_comb;
  wire [31:0] p3_add_80348_comb;
  wire [31:0] p3_add_80349_comb;
  wire [31:0] p3_add_80350_comb;
  wire [31:0] p3_add_80351_comb;
  wire [31:0] p3_add_80352_comb;
  wire [31:0] p3_add_80353_comb;
  wire [31:0] p3_add_80354_comb;
  wire [31:0] p3_add_80355_comb;
  wire [31:0] p3_add_80356_comb;
  wire [31:0] p3_add_80357_comb;
  wire [31:0] p3_add_80358_comb;
  wire [31:0] p3_add_80359_comb;
  wire [31:0] p3_add_80360_comb;
  wire [31:0] p3_add_80361_comb;
  wire [31:0] p3_add_80362_comb;
  wire [31:0] p3_add_80363_comb;
  wire [31:0] p3_add_80364_comb;
  wire [31:0] p3_add_80365_comb;
  wire [31:0] p3_add_80366_comb;
  wire [31:0] p3_add_80367_comb;
  wire [31:0] p3_add_80368_comb;
  wire [31:0] p3_add_80369_comb;
  wire [31:0] p3_add_80370_comb;
  wire [31:0] p3_add_80371_comb;
  wire [31:0] p3_add_80372_comb;
  wire [31:0] p3_add_80373_comb;
  wire [31:0] p3_add_80374_comb;
  wire [31:0] p3_add_80375_comb;
  wire [31:0] p3_add_80376_comb;
  wire [31:0] p3_add_80377_comb;
  wire [31:0] p3_add_80378_comb;
  wire [31:0] p3_add_80379_comb;
  wire [31:0] p3_add_80380_comb;
  wire [31:0] p3_add_80381_comb;
  wire [31:0] p3_add_80382_comb;
  wire [31:0] p3_add_80383_comb;
  wire [31:0] p3_add_80384_comb;
  wire [31:0] p3_add_80385_comb;
  wire [31:0] p3_add_80386_comb;
  wire [31:0] p3_add_80387_comb;
  wire [31:0] p3_add_80388_comb;
  wire [31:0] p3_add_80389_comb;
  wire [31:0] p3_add_80390_comb;
  wire [31:0] p3_add_80391_comb;
  wire [31:0] p3_add_80392_comb;
  wire [31:0] p3_add_80393_comb;
  wire [31:0] p3_add_80394_comb;
  wire [31:0] p3_add_80395_comb;
  wire [31:0] p3_add_80396_comb;
  wire [31:0] p3_add_80397_comb;
  wire [31:0] p3_add_80398_comb;
  wire [31:0] p3_add_80399_comb;
  wire [31:0] p3_add_80400_comb;
  wire [31:0] p3_add_80401_comb;
  wire [31:0] p3_add_80402_comb;
  wire [31:0] p3_add_80403_comb;
  wire [31:0] p3_add_80404_comb;
  wire [31:0] p3_add_80405_comb;
  wire [31:0] p3_add_80406_comb;
  wire [31:0] p3_add_80407_comb;
  wire [31:0] p3_add_80408_comb;
  wire [31:0] p3_add_80409_comb;
  wire [31:0] p3_add_80410_comb;
  wire [31:0] p3_add_80411_comb;
  wire [31:0] p3_add_80412_comb;
  wire [31:0] p3_add_80413_comb;
  wire [31:0] p3_add_80414_comb;
  wire [31:0] p3_add_80415_comb;
  wire [31:0] p3_add_80416_comb;
  wire [31:0] p3_add_80417_comb;
  wire [31:0] p3_add_80418_comb;
  wire [31:0] p3_add_80419_comb;
  wire [31:0] p3_add_80420_comb;
  wire [31:0] p3_add_80421_comb;
  wire [31:0] p3_add_80422_comb;
  wire [31:0] p3_add_80423_comb;
  wire [31:0] p3_add_80424_comb;
  wire [31:0] p3_add_80425_comb;
  wire [31:0] p3_add_80426_comb;
  wire [31:0] p3_add_80427_comb;
  wire [31:0] p3_add_80428_comb;
  wire [31:0] p3_add_80429_comb;
  wire [31:0] p3_add_80430_comb;
  wire [31:0] p3_add_80431_comb;
  wire [31:0] p3_add_80432_comb;
  wire [31:0] p3_add_80433_comb;
  wire [31:0] p3_add_80434_comb;
  wire [31:0] p3_add_80435_comb;
  wire [31:0] p3_add_80436_comb;
  wire [31:0] p3_add_80437_comb;
  wire [31:0] p3_add_80438_comb;
  wire [31:0] p3_add_80439_comb;
  wire [31:0] p3_add_80440_comb;
  wire [31:0] p3_add_80441_comb;
  wire [31:0] p3_add_80442_comb;
  wire [31:0] p3_add_80443_comb;
  wire [31:0] p3_add_80444_comb;
  wire [31:0] p3_add_80445_comb;
  wire [31:0] p3_add_80446_comb;
  wire [31:0] p3_add_80447_comb;
  wire [31:0] p3_add_80448_comb;
  wire [31:0] p3_add_80449_comb;
  wire [31:0] p3_add_80450_comb;
  wire [31:0] p3_add_80451_comb;
  wire [31:0] p3_add_80452_comb;
  wire [31:0] p3_add_80453_comb;
  wire [31:0] p3_add_80454_comb;
  wire [31:0] p3_add_80455_comb;
  wire [31:0] p3_add_80456_comb;
  wire [31:0] p3_add_80457_comb;
  wire [31:0] p3_add_80458_comb;
  wire [31:0] p3_add_80459_comb;
  wire [31:0] p3_add_80460_comb;
  wire [31:0] p3_add_80461_comb;
  wire [31:0] p3_add_80462_comb;
  wire [31:0] p3_add_80463_comb;
  wire [31:0] p3_add_80464_comb;
  wire [31:0] p3_add_80465_comb;
  wire [31:0] p3_add_80466_comb;
  wire [31:0] p3_add_80467_comb;
  wire [31:0] p3_add_80468_comb;
  wire [31:0] p3_add_80469_comb;
  wire [31:0] p3_add_80470_comb;
  wire [31:0] p3_add_80471_comb;
  wire [31:0] p3_add_80472_comb;
  wire [31:0] p3_add_80473_comb;
  wire [31:0] p3_add_80474_comb;
  wire [31:0] p3_add_80475_comb;
  wire [31:0] p3_add_80476_comb;
  wire [31:0] p3_add_80477_comb;
  wire [31:0] p3_add_80478_comb;
  wire [31:0] p3_add_80479_comb;
  wire [31:0] p3_add_80480_comb;
  wire [31:0] p3_add_80481_comb;
  wire [31:0] p3_add_80482_comb;
  wire [31:0] p3_add_80483_comb;
  wire [31:0] p3_add_80484_comb;
  wire [31:0] p3_add_80485_comb;
  wire [31:0] p3_add_80486_comb;
  wire [31:0] p3_add_80487_comb;
  wire [31:0] p3_add_80488_comb;
  wire [31:0] p3_add_80489_comb;
  wire [31:0] p3_add_80490_comb;
  wire [31:0] p3_add_80491_comb;
  wire [31:0] p3_add_80492_comb;
  wire [31:0] p3_add_80493_comb;
  wire [31:0] p3_add_80494_comb;
  wire [31:0] p3_add_80495_comb;
  wire [31:0] p3_add_80496_comb;
  wire [31:0] p3_add_80497_comb;
  wire [31:0] p3_add_80498_comb;
  assign p3_add_80299_comb = p2_add_79186 + p2_add_79187;
  assign p3_add_80300_comb = p2_add_79190 + p2_add_79191;
  assign p3_add_80301_comb = p2_add_79194 + p2_add_79195;
  assign p3_add_80302_comb = p2_add_79198 + p2_add_79199;
  assign p3_add_80303_comb = p2_add_79202 + p2_add_79203;
  assign p3_add_80304_comb = p2_add_79206 + p2_add_79207;
  assign p3_add_80305_comb = p2_add_79210 + p2_add_79211;
  assign p3_add_80306_comb = p2_add_79214 + p2_add_79215;
  assign p3_add_80307_comb = p2_add_79218 + p2_add_79219;
  assign p3_add_80308_comb = p2_add_79222 + p2_add_79223;
  assign p3_add_80309_comb = p2_add_79226 + p2_add_79227;
  assign p3_add_80310_comb = p2_add_79230 + p2_add_79231;
  assign p3_add_80311_comb = p2_add_79234 + p2_add_79235;
  assign p3_add_80312_comb = p2_add_79238 + p2_add_79239;
  assign p3_add_80313_comb = p2_add_79242 + p2_add_79243;
  assign p3_add_80314_comb = p2_add_79246 + p2_add_79247;
  assign p3_add_80315_comb = p2_add_79250 + p2_add_79251;
  assign p3_add_80316_comb = p2_add_79254 + p2_add_79255;
  assign p3_add_80317_comb = p2_add_79258 + p2_add_79259;
  assign p3_add_80318_comb = p2_add_79262 + p2_add_79263;
  assign p3_add_80319_comb = p2_add_79266 + p2_add_79267;
  assign p3_add_80320_comb = p2_add_79270 + p2_add_79271;
  assign p3_add_80321_comb = p2_add_79274 + p2_add_79275;
  assign p3_add_80322_comb = p2_add_79278 + p2_add_79279;
  assign p3_add_80323_comb = p2_add_79282 + p2_add_79283;
  assign p3_add_80324_comb = p2_add_79286 + p2_add_79287;
  assign p3_add_80325_comb = p2_add_79290 + p2_add_79291;
  assign p3_add_80326_comb = p2_add_79294 + p2_add_79295;
  assign p3_add_80327_comb = p2_add_79298 + p2_add_79299;
  assign p3_add_80328_comb = p2_add_79302 + p2_add_79303;
  assign p3_add_80329_comb = p2_add_79306 + p2_add_79307;
  assign p3_add_80330_comb = p2_add_79310 + p2_add_79311;
  assign p3_add_80331_comb = p2_add_79314 + p2_add_79315;
  assign p3_add_80332_comb = p2_add_79318 + p2_add_79319;
  assign p3_add_80333_comb = p2_add_79322 + p2_add_79323;
  assign p3_add_80334_comb = p2_add_79326 + p2_add_79327;
  assign p3_add_80335_comb = p2_add_79330 + p2_add_79331;
  assign p3_add_80336_comb = p2_add_79334 + p2_add_79335;
  assign p3_add_80337_comb = p2_add_79338 + p2_add_79339;
  assign p3_add_80338_comb = p2_add_79342 + p2_add_79343;
  assign p3_add_80339_comb = p2_add_79346 + p2_add_79347;
  assign p3_add_80340_comb = p2_add_79350 + p2_add_79351;
  assign p3_add_80341_comb = p2_add_79354 + p2_add_79355;
  assign p3_add_80342_comb = p2_add_79358 + p2_add_79359;
  assign p3_add_80343_comb = p2_add_79362 + p2_add_79363;
  assign p3_add_80344_comb = p2_add_79366 + p2_add_79367;
  assign p3_add_80345_comb = p2_add_79370 + p2_add_79371;
  assign p3_add_80346_comb = p2_add_79374 + p2_add_79375;
  assign p3_add_80347_comb = p2_add_79378 + p2_add_79379;
  assign p3_add_80348_comb = p2_add_79382 + p2_add_79383;
  assign p3_add_80349_comb = p2_add_79386 + p2_add_79387;
  assign p3_add_80350_comb = p2_add_79390 + p2_add_79391;
  assign p3_add_80351_comb = p2_add_79394 + p2_add_79395;
  assign p3_add_80352_comb = p2_add_79398 + p2_add_79399;
  assign p3_add_80353_comb = p2_add_79402 + p2_add_79403;
  assign p3_add_80354_comb = p2_add_79406 + p2_add_79407;
  assign p3_add_80355_comb = p2_add_79410 + p2_add_79411;
  assign p3_add_80356_comb = p2_add_79414 + p2_add_79415;
  assign p3_add_80357_comb = p2_add_79418 + p2_add_79419;
  assign p3_add_80358_comb = p2_add_79422 + p2_add_79423;
  assign p3_add_80359_comb = p2_add_79426 + p2_add_79427;
  assign p3_add_80360_comb = p2_add_79430 + p2_add_79431;
  assign p3_add_80361_comb = p2_add_79434 + p2_add_79435;
  assign p3_add_80362_comb = p2_add_79438 + p2_add_79439;
  assign p3_add_80363_comb = p2_add_79442 + p2_add_79443;
  assign p3_add_80364_comb = p2_add_79446 + p2_add_79447;
  assign p3_add_80365_comb = p2_add_79450 + p2_add_79451;
  assign p3_add_80366_comb = p2_add_79454 + p2_add_79455;
  assign p3_add_80367_comb = p2_add_79458 + p2_add_79459;
  assign p3_add_80368_comb = p2_add_79462 + p2_add_79463;
  assign p3_add_80369_comb = p2_add_79466 + p2_add_79467;
  assign p3_add_80370_comb = p2_add_79470 + p2_add_79471;
  assign p3_add_80371_comb = p2_add_79474 + p2_add_79475;
  assign p3_add_80372_comb = p2_add_79478 + p2_add_79479;
  assign p3_add_80373_comb = p2_add_79482 + p2_add_79483;
  assign p3_add_80374_comb = p2_add_79486 + p2_add_79487;
  assign p3_add_80375_comb = p2_add_79490 + p2_add_79491;
  assign p3_add_80376_comb = p2_add_79494 + p2_add_79495;
  assign p3_add_80377_comb = p2_add_79498 + p2_add_79499;
  assign p3_add_80378_comb = p2_add_79502 + p2_add_79503;
  assign p3_add_80379_comb = p2_add_79506 + p2_add_79507;
  assign p3_add_80380_comb = p2_add_79510 + p2_add_79511;
  assign p3_add_80381_comb = p2_add_79514 + p2_add_79515;
  assign p3_add_80382_comb = p2_add_79518 + p2_add_79519;
  assign p3_add_80383_comb = p2_add_79522 + p2_add_79523;
  assign p3_add_80384_comb = p2_add_79526 + p2_add_79527;
  assign p3_add_80385_comb = p2_add_79530 + p2_add_79531;
  assign p3_add_80386_comb = p2_add_79534 + p2_add_79535;
  assign p3_add_80387_comb = p2_add_79538 + p2_add_79539;
  assign p3_add_80388_comb = p2_add_79542 + p2_add_79543;
  assign p3_add_80389_comb = p2_add_79546 + p2_add_79547;
  assign p3_add_80390_comb = p2_add_79550 + p2_add_79551;
  assign p3_add_80391_comb = p2_add_79554 + p2_add_79555;
  assign p3_add_80392_comb = p2_add_79558 + p2_add_79559;
  assign p3_add_80393_comb = p2_add_79562 + p2_add_79563;
  assign p3_add_80394_comb = p2_add_79566 + p2_add_79567;
  assign p3_add_80395_comb = p2_add_79570 + p2_add_79571;
  assign p3_add_80396_comb = p2_add_79574 + p2_add_79575;
  assign p3_add_80397_comb = p2_add_79578 + p2_add_79579;
  assign p3_add_80398_comb = p2_add_79582 + p2_add_79583;
  assign p3_add_80399_comb = p3_add_80299_comb + p2_add_79586;
  assign p3_add_80400_comb = p3_add_80300_comb + p2_add_79587;
  assign p3_add_80401_comb = p3_add_80301_comb + p2_add_79588;
  assign p3_add_80402_comb = p3_add_80302_comb + p2_add_79589;
  assign p3_add_80403_comb = p3_add_80303_comb + p2_add_79590;
  assign p3_add_80404_comb = p3_add_80304_comb + p2_add_79591;
  assign p3_add_80405_comb = p3_add_80305_comb + p2_add_79592;
  assign p3_add_80406_comb = p3_add_80306_comb + p2_add_79593;
  assign p3_add_80407_comb = p3_add_80307_comb + p2_add_79594;
  assign p3_add_80408_comb = p3_add_80308_comb + p2_add_79595;
  assign p3_add_80409_comb = p3_add_80309_comb + p2_add_79596;
  assign p3_add_80410_comb = p3_add_80310_comb + p2_add_79597;
  assign p3_add_80411_comb = p3_add_80311_comb + p2_add_79598;
  assign p3_add_80412_comb = p3_add_80312_comb + p2_add_79599;
  assign p3_add_80413_comb = p3_add_80313_comb + p2_add_79600;
  assign p3_add_80414_comb = p3_add_80314_comb + p2_add_79601;
  assign p3_add_80415_comb = p3_add_80315_comb + p2_add_79602;
  assign p3_add_80416_comb = p3_add_80316_comb + p2_add_79603;
  assign p3_add_80417_comb = p3_add_80317_comb + p2_add_79604;
  assign p3_add_80418_comb = p3_add_80318_comb + p2_add_79605;
  assign p3_add_80419_comb = p3_add_80319_comb + p2_add_79606;
  assign p3_add_80420_comb = p3_add_80320_comb + p2_add_79607;
  assign p3_add_80421_comb = p3_add_80321_comb + p2_add_79608;
  assign p3_add_80422_comb = p3_add_80322_comb + p2_add_79609;
  assign p3_add_80423_comb = p3_add_80323_comb + p2_add_79610;
  assign p3_add_80424_comb = p3_add_80324_comb + p2_add_79611;
  assign p3_add_80425_comb = p3_add_80325_comb + p2_add_79612;
  assign p3_add_80426_comb = p3_add_80326_comb + p2_add_79613;
  assign p3_add_80427_comb = p3_add_80327_comb + p2_add_79614;
  assign p3_add_80428_comb = p3_add_80328_comb + p2_add_79615;
  assign p3_add_80429_comb = p3_add_80329_comb + p2_add_79616;
  assign p3_add_80430_comb = p3_add_80330_comb + p2_add_79617;
  assign p3_add_80431_comb = p3_add_80331_comb + p2_add_79618;
  assign p3_add_80432_comb = p3_add_80332_comb + p2_add_79619;
  assign p3_add_80433_comb = p3_add_80333_comb + p2_add_79620;
  assign p3_add_80434_comb = p3_add_80334_comb + p2_add_79621;
  assign p3_add_80435_comb = p3_add_80335_comb + p2_add_79622;
  assign p3_add_80436_comb = p3_add_80336_comb + p2_add_79623;
  assign p3_add_80437_comb = p3_add_80337_comb + p2_add_79624;
  assign p3_add_80438_comb = p3_add_80338_comb + p2_add_79625;
  assign p3_add_80439_comb = p3_add_80339_comb + p2_add_79626;
  assign p3_add_80440_comb = p3_add_80340_comb + p2_add_79627;
  assign p3_add_80441_comb = p3_add_80341_comb + p2_add_79628;
  assign p3_add_80442_comb = p3_add_80342_comb + p2_add_79629;
  assign p3_add_80443_comb = p3_add_80343_comb + p2_add_79630;
  assign p3_add_80444_comb = p3_add_80344_comb + p2_add_79631;
  assign p3_add_80445_comb = p3_add_80345_comb + p2_add_79632;
  assign p3_add_80446_comb = p3_add_80346_comb + p2_add_79633;
  assign p3_add_80447_comb = p3_add_80347_comb + p2_add_79634;
  assign p3_add_80448_comb = p3_add_80348_comb + p2_add_79635;
  assign p3_add_80449_comb = p3_add_80349_comb + p2_add_79636;
  assign p3_add_80450_comb = p3_add_80350_comb + p2_add_79637;
  assign p3_add_80451_comb = p3_add_80351_comb + p2_add_79638;
  assign p3_add_80452_comb = p3_add_80352_comb + p2_add_79639;
  assign p3_add_80453_comb = p3_add_80353_comb + p2_add_79640;
  assign p3_add_80454_comb = p3_add_80354_comb + p2_add_79641;
  assign p3_add_80455_comb = p3_add_80355_comb + p2_add_79642;
  assign p3_add_80456_comb = p3_add_80356_comb + p2_add_79643;
  assign p3_add_80457_comb = p3_add_80357_comb + p2_add_79644;
  assign p3_add_80458_comb = p3_add_80358_comb + p2_add_79645;
  assign p3_add_80459_comb = p3_add_80359_comb + p2_add_79646;
  assign p3_add_80460_comb = p3_add_80360_comb + p2_add_79647;
  assign p3_add_80461_comb = p3_add_80361_comb + p2_add_79648;
  assign p3_add_80462_comb = p3_add_80362_comb + p2_add_79649;
  assign p3_add_80463_comb = p3_add_80363_comb + p2_add_79650;
  assign p3_add_80464_comb = p3_add_80364_comb + p2_add_79651;
  assign p3_add_80465_comb = p3_add_80365_comb + p2_add_79652;
  assign p3_add_80466_comb = p3_add_80366_comb + p2_add_79653;
  assign p3_add_80467_comb = p3_add_80367_comb + p2_add_79654;
  assign p3_add_80468_comb = p3_add_80368_comb + p2_add_79655;
  assign p3_add_80469_comb = p3_add_80369_comb + p2_add_79656;
  assign p3_add_80470_comb = p3_add_80370_comb + p2_add_79657;
  assign p3_add_80471_comb = p3_add_80371_comb + p2_add_79658;
  assign p3_add_80472_comb = p3_add_80372_comb + p2_add_79659;
  assign p3_add_80473_comb = p3_add_80373_comb + p2_add_79660;
  assign p3_add_80474_comb = p3_add_80374_comb + p2_add_79661;
  assign p3_add_80475_comb = p3_add_80375_comb + p2_add_79662;
  assign p3_add_80476_comb = p3_add_80376_comb + p2_add_79663;
  assign p3_add_80477_comb = p3_add_80377_comb + p2_add_79664;
  assign p3_add_80478_comb = p3_add_80378_comb + p2_add_79665;
  assign p3_add_80479_comb = p3_add_80379_comb + p2_add_79666;
  assign p3_add_80480_comb = p3_add_80380_comb + p2_add_79667;
  assign p3_add_80481_comb = p3_add_80381_comb + p2_add_79668;
  assign p3_add_80482_comb = p3_add_80382_comb + p2_add_79669;
  assign p3_add_80483_comb = p3_add_80383_comb + p2_add_79670;
  assign p3_add_80484_comb = p3_add_80384_comb + p2_add_79671;
  assign p3_add_80485_comb = p3_add_80385_comb + p2_add_79672;
  assign p3_add_80486_comb = p3_add_80386_comb + p2_add_79673;
  assign p3_add_80487_comb = p3_add_80387_comb + p2_add_79674;
  assign p3_add_80488_comb = p3_add_80388_comb + p2_add_79675;
  assign p3_add_80489_comb = p3_add_80389_comb + p2_add_79676;
  assign p3_add_80490_comb = p3_add_80390_comb + p2_add_79677;
  assign p3_add_80491_comb = p3_add_80391_comb + p2_add_79678;
  assign p3_add_80492_comb = p3_add_80392_comb + p2_add_79679;
  assign p3_add_80493_comb = p3_add_80393_comb + p2_add_79680;
  assign p3_add_80494_comb = p3_add_80394_comb + p2_add_79681;
  assign p3_add_80495_comb = p3_add_80395_comb + p2_add_79682;
  assign p3_add_80496_comb = p3_add_80396_comb + p2_add_79683;
  assign p3_add_80497_comb = p3_add_80397_comb + p2_add_79684;
  assign p3_add_80498_comb = p3_add_80398_comb + p2_add_79685;

  // Registers for pipe stage 3:
  reg [31:0] p3_add_80399;
  reg [31:0] p3_add_80400;
  reg [31:0] p3_add_80401;
  reg [31:0] p3_add_80402;
  reg [31:0] p3_add_80403;
  reg [31:0] p3_add_80404;
  reg [31:0] p3_add_80405;
  reg [31:0] p3_add_80406;
  reg [31:0] p3_add_80407;
  reg [31:0] p3_add_80408;
  reg [31:0] p3_add_80409;
  reg [31:0] p3_add_80410;
  reg [31:0] p3_add_80411;
  reg [31:0] p3_add_80412;
  reg [31:0] p3_add_80413;
  reg [31:0] p3_add_80414;
  reg [31:0] p3_add_80415;
  reg [31:0] p3_add_80416;
  reg [31:0] p3_add_80417;
  reg [31:0] p3_add_80418;
  reg [31:0] p3_add_80419;
  reg [31:0] p3_add_80420;
  reg [31:0] p3_add_80421;
  reg [31:0] p3_add_80422;
  reg [31:0] p3_add_80423;
  reg [31:0] p3_add_80424;
  reg [31:0] p3_add_80425;
  reg [31:0] p3_add_80426;
  reg [31:0] p3_add_80427;
  reg [31:0] p3_add_80428;
  reg [31:0] p3_add_80429;
  reg [31:0] p3_add_80430;
  reg [31:0] p3_add_80431;
  reg [31:0] p3_add_80432;
  reg [31:0] p3_add_80433;
  reg [31:0] p3_add_80434;
  reg [31:0] p3_add_80435;
  reg [31:0] p3_add_80436;
  reg [31:0] p3_add_80437;
  reg [31:0] p3_add_80438;
  reg [31:0] p3_add_80439;
  reg [31:0] p3_add_80440;
  reg [31:0] p3_add_80441;
  reg [31:0] p3_add_80442;
  reg [31:0] p3_add_80443;
  reg [31:0] p3_add_80444;
  reg [31:0] p3_add_80445;
  reg [31:0] p3_add_80446;
  reg [31:0] p3_add_80447;
  reg [31:0] p3_add_80448;
  reg [31:0] p3_add_80449;
  reg [31:0] p3_add_80450;
  reg [31:0] p3_add_80451;
  reg [31:0] p3_add_80452;
  reg [31:0] p3_add_80453;
  reg [31:0] p3_add_80454;
  reg [31:0] p3_add_80455;
  reg [31:0] p3_add_80456;
  reg [31:0] p3_add_80457;
  reg [31:0] p3_add_80458;
  reg [31:0] p3_add_80459;
  reg [31:0] p3_add_80460;
  reg [31:0] p3_add_80461;
  reg [31:0] p3_add_80462;
  reg [31:0] p3_add_80463;
  reg [31:0] p3_add_80464;
  reg [31:0] p3_add_80465;
  reg [31:0] p3_add_80466;
  reg [31:0] p3_add_80467;
  reg [31:0] p3_add_80468;
  reg [31:0] p3_add_80469;
  reg [31:0] p3_add_80470;
  reg [31:0] p3_add_80471;
  reg [31:0] p3_add_80472;
  reg [31:0] p3_add_80473;
  reg [31:0] p3_add_80474;
  reg [31:0] p3_add_80475;
  reg [31:0] p3_add_80476;
  reg [31:0] p3_add_80477;
  reg [31:0] p3_add_80478;
  reg [31:0] p3_add_80479;
  reg [31:0] p3_add_80480;
  reg [31:0] p3_add_80481;
  reg [31:0] p3_add_80482;
  reg [31:0] p3_add_80483;
  reg [31:0] p3_add_80484;
  reg [31:0] p3_add_80485;
  reg [31:0] p3_add_80486;
  reg [31:0] p3_add_80487;
  reg [31:0] p3_add_80488;
  reg [31:0] p3_add_80489;
  reg [31:0] p3_add_80490;
  reg [31:0] p3_add_80491;
  reg [31:0] p3_add_80492;
  reg [31:0] p3_add_80493;
  reg [31:0] p3_add_80494;
  reg [31:0] p3_add_80495;
  reg [31:0] p3_add_80496;
  reg [31:0] p3_add_80497;
  reg [31:0] p3_add_80498;
  always_ff @ (posedge clk) begin
    p3_add_80399 <= p3_add_80399_comb;
    p3_add_80400 <= p3_add_80400_comb;
    p3_add_80401 <= p3_add_80401_comb;
    p3_add_80402 <= p3_add_80402_comb;
    p3_add_80403 <= p3_add_80403_comb;
    p3_add_80404 <= p3_add_80404_comb;
    p3_add_80405 <= p3_add_80405_comb;
    p3_add_80406 <= p3_add_80406_comb;
    p3_add_80407 <= p3_add_80407_comb;
    p3_add_80408 <= p3_add_80408_comb;
    p3_add_80409 <= p3_add_80409_comb;
    p3_add_80410 <= p3_add_80410_comb;
    p3_add_80411 <= p3_add_80411_comb;
    p3_add_80412 <= p3_add_80412_comb;
    p3_add_80413 <= p3_add_80413_comb;
    p3_add_80414 <= p3_add_80414_comb;
    p3_add_80415 <= p3_add_80415_comb;
    p3_add_80416 <= p3_add_80416_comb;
    p3_add_80417 <= p3_add_80417_comb;
    p3_add_80418 <= p3_add_80418_comb;
    p3_add_80419 <= p3_add_80419_comb;
    p3_add_80420 <= p3_add_80420_comb;
    p3_add_80421 <= p3_add_80421_comb;
    p3_add_80422 <= p3_add_80422_comb;
    p3_add_80423 <= p3_add_80423_comb;
    p3_add_80424 <= p3_add_80424_comb;
    p3_add_80425 <= p3_add_80425_comb;
    p3_add_80426 <= p3_add_80426_comb;
    p3_add_80427 <= p3_add_80427_comb;
    p3_add_80428 <= p3_add_80428_comb;
    p3_add_80429 <= p3_add_80429_comb;
    p3_add_80430 <= p3_add_80430_comb;
    p3_add_80431 <= p3_add_80431_comb;
    p3_add_80432 <= p3_add_80432_comb;
    p3_add_80433 <= p3_add_80433_comb;
    p3_add_80434 <= p3_add_80434_comb;
    p3_add_80435 <= p3_add_80435_comb;
    p3_add_80436 <= p3_add_80436_comb;
    p3_add_80437 <= p3_add_80437_comb;
    p3_add_80438 <= p3_add_80438_comb;
    p3_add_80439 <= p3_add_80439_comb;
    p3_add_80440 <= p3_add_80440_comb;
    p3_add_80441 <= p3_add_80441_comb;
    p3_add_80442 <= p3_add_80442_comb;
    p3_add_80443 <= p3_add_80443_comb;
    p3_add_80444 <= p3_add_80444_comb;
    p3_add_80445 <= p3_add_80445_comb;
    p3_add_80446 <= p3_add_80446_comb;
    p3_add_80447 <= p3_add_80447_comb;
    p3_add_80448 <= p3_add_80448_comb;
    p3_add_80449 <= p3_add_80449_comb;
    p3_add_80450 <= p3_add_80450_comb;
    p3_add_80451 <= p3_add_80451_comb;
    p3_add_80452 <= p3_add_80452_comb;
    p3_add_80453 <= p3_add_80453_comb;
    p3_add_80454 <= p3_add_80454_comb;
    p3_add_80455 <= p3_add_80455_comb;
    p3_add_80456 <= p3_add_80456_comb;
    p3_add_80457 <= p3_add_80457_comb;
    p3_add_80458 <= p3_add_80458_comb;
    p3_add_80459 <= p3_add_80459_comb;
    p3_add_80460 <= p3_add_80460_comb;
    p3_add_80461 <= p3_add_80461_comb;
    p3_add_80462 <= p3_add_80462_comb;
    p3_add_80463 <= p3_add_80463_comb;
    p3_add_80464 <= p3_add_80464_comb;
    p3_add_80465 <= p3_add_80465_comb;
    p3_add_80466 <= p3_add_80466_comb;
    p3_add_80467 <= p3_add_80467_comb;
    p3_add_80468 <= p3_add_80468_comb;
    p3_add_80469 <= p3_add_80469_comb;
    p3_add_80470 <= p3_add_80470_comb;
    p3_add_80471 <= p3_add_80471_comb;
    p3_add_80472 <= p3_add_80472_comb;
    p3_add_80473 <= p3_add_80473_comb;
    p3_add_80474 <= p3_add_80474_comb;
    p3_add_80475 <= p3_add_80475_comb;
    p3_add_80476 <= p3_add_80476_comb;
    p3_add_80477 <= p3_add_80477_comb;
    p3_add_80478 <= p3_add_80478_comb;
    p3_add_80479 <= p3_add_80479_comb;
    p3_add_80480 <= p3_add_80480_comb;
    p3_add_80481 <= p3_add_80481_comb;
    p3_add_80482 <= p3_add_80482_comb;
    p3_add_80483 <= p3_add_80483_comb;
    p3_add_80484 <= p3_add_80484_comb;
    p3_add_80485 <= p3_add_80485_comb;
    p3_add_80486 <= p3_add_80486_comb;
    p3_add_80487 <= p3_add_80487_comb;
    p3_add_80488 <= p3_add_80488_comb;
    p3_add_80489 <= p3_add_80489_comb;
    p3_add_80490 <= p3_add_80490_comb;
    p3_add_80491 <= p3_add_80491_comb;
    p3_add_80492 <= p3_add_80492_comb;
    p3_add_80493 <= p3_add_80493_comb;
    p3_add_80494 <= p3_add_80494_comb;
    p3_add_80495 <= p3_add_80495_comb;
    p3_add_80496 <= p3_add_80496_comb;
    p3_add_80497 <= p3_add_80497_comb;
    p3_add_80498 <= p3_add_80498_comb;
  end

  // ===== Pipe stage 4:

  // Registers for pipe stage 4:
  reg [31:0] p4_add_80399;
  reg [31:0] p4_add_80400;
  reg [31:0] p4_add_80401;
  reg [31:0] p4_add_80402;
  reg [31:0] p4_add_80403;
  reg [31:0] p4_add_80404;
  reg [31:0] p4_add_80405;
  reg [31:0] p4_add_80406;
  reg [31:0] p4_add_80407;
  reg [31:0] p4_add_80408;
  reg [31:0] p4_add_80409;
  reg [31:0] p4_add_80410;
  reg [31:0] p4_add_80411;
  reg [31:0] p4_add_80412;
  reg [31:0] p4_add_80413;
  reg [31:0] p4_add_80414;
  reg [31:0] p4_add_80415;
  reg [31:0] p4_add_80416;
  reg [31:0] p4_add_80417;
  reg [31:0] p4_add_80418;
  reg [31:0] p4_add_80419;
  reg [31:0] p4_add_80420;
  reg [31:0] p4_add_80421;
  reg [31:0] p4_add_80422;
  reg [31:0] p4_add_80423;
  reg [31:0] p4_add_80424;
  reg [31:0] p4_add_80425;
  reg [31:0] p4_add_80426;
  reg [31:0] p4_add_80427;
  reg [31:0] p4_add_80428;
  reg [31:0] p4_add_80429;
  reg [31:0] p4_add_80430;
  reg [31:0] p4_add_80431;
  reg [31:0] p4_add_80432;
  reg [31:0] p4_add_80433;
  reg [31:0] p4_add_80434;
  reg [31:0] p4_add_80435;
  reg [31:0] p4_add_80436;
  reg [31:0] p4_add_80437;
  reg [31:0] p4_add_80438;
  reg [31:0] p4_add_80439;
  reg [31:0] p4_add_80440;
  reg [31:0] p4_add_80441;
  reg [31:0] p4_add_80442;
  reg [31:0] p4_add_80443;
  reg [31:0] p4_add_80444;
  reg [31:0] p4_add_80445;
  reg [31:0] p4_add_80446;
  reg [31:0] p4_add_80447;
  reg [31:0] p4_add_80448;
  reg [31:0] p4_add_80449;
  reg [31:0] p4_add_80450;
  reg [31:0] p4_add_80451;
  reg [31:0] p4_add_80452;
  reg [31:0] p4_add_80453;
  reg [31:0] p4_add_80454;
  reg [31:0] p4_add_80455;
  reg [31:0] p4_add_80456;
  reg [31:0] p4_add_80457;
  reg [31:0] p4_add_80458;
  reg [31:0] p4_add_80459;
  reg [31:0] p4_add_80460;
  reg [31:0] p4_add_80461;
  reg [31:0] p4_add_80462;
  reg [31:0] p4_add_80463;
  reg [31:0] p4_add_80464;
  reg [31:0] p4_add_80465;
  reg [31:0] p4_add_80466;
  reg [31:0] p4_add_80467;
  reg [31:0] p4_add_80468;
  reg [31:0] p4_add_80469;
  reg [31:0] p4_add_80470;
  reg [31:0] p4_add_80471;
  reg [31:0] p4_add_80472;
  reg [31:0] p4_add_80473;
  reg [31:0] p4_add_80474;
  reg [31:0] p4_add_80475;
  reg [31:0] p4_add_80476;
  reg [31:0] p4_add_80477;
  reg [31:0] p4_add_80478;
  reg [31:0] p4_add_80479;
  reg [31:0] p4_add_80480;
  reg [31:0] p4_add_80481;
  reg [31:0] p4_add_80482;
  reg [31:0] p4_add_80483;
  reg [31:0] p4_add_80484;
  reg [31:0] p4_add_80485;
  reg [31:0] p4_add_80486;
  reg [31:0] p4_add_80487;
  reg [31:0] p4_add_80488;
  reg [31:0] p4_add_80489;
  reg [31:0] p4_add_80490;
  reg [31:0] p4_add_80491;
  reg [31:0] p4_add_80492;
  reg [31:0] p4_add_80493;
  reg [31:0] p4_add_80494;
  reg [31:0] p4_add_80495;
  reg [31:0] p4_add_80496;
  reg [31:0] p4_add_80497;
  reg [31:0] p4_add_80498;
  always_ff @ (posedge clk) begin
    p4_add_80399 <= p3_add_80399;
    p4_add_80400 <= p3_add_80400;
    p4_add_80401 <= p3_add_80401;
    p4_add_80402 <= p3_add_80402;
    p4_add_80403 <= p3_add_80403;
    p4_add_80404 <= p3_add_80404;
    p4_add_80405 <= p3_add_80405;
    p4_add_80406 <= p3_add_80406;
    p4_add_80407 <= p3_add_80407;
    p4_add_80408 <= p3_add_80408;
    p4_add_80409 <= p3_add_80409;
    p4_add_80410 <= p3_add_80410;
    p4_add_80411 <= p3_add_80411;
    p4_add_80412 <= p3_add_80412;
    p4_add_80413 <= p3_add_80413;
    p4_add_80414 <= p3_add_80414;
    p4_add_80415 <= p3_add_80415;
    p4_add_80416 <= p3_add_80416;
    p4_add_80417 <= p3_add_80417;
    p4_add_80418 <= p3_add_80418;
    p4_add_80419 <= p3_add_80419;
    p4_add_80420 <= p3_add_80420;
    p4_add_80421 <= p3_add_80421;
    p4_add_80422 <= p3_add_80422;
    p4_add_80423 <= p3_add_80423;
    p4_add_80424 <= p3_add_80424;
    p4_add_80425 <= p3_add_80425;
    p4_add_80426 <= p3_add_80426;
    p4_add_80427 <= p3_add_80427;
    p4_add_80428 <= p3_add_80428;
    p4_add_80429 <= p3_add_80429;
    p4_add_80430 <= p3_add_80430;
    p4_add_80431 <= p3_add_80431;
    p4_add_80432 <= p3_add_80432;
    p4_add_80433 <= p3_add_80433;
    p4_add_80434 <= p3_add_80434;
    p4_add_80435 <= p3_add_80435;
    p4_add_80436 <= p3_add_80436;
    p4_add_80437 <= p3_add_80437;
    p4_add_80438 <= p3_add_80438;
    p4_add_80439 <= p3_add_80439;
    p4_add_80440 <= p3_add_80440;
    p4_add_80441 <= p3_add_80441;
    p4_add_80442 <= p3_add_80442;
    p4_add_80443 <= p3_add_80443;
    p4_add_80444 <= p3_add_80444;
    p4_add_80445 <= p3_add_80445;
    p4_add_80446 <= p3_add_80446;
    p4_add_80447 <= p3_add_80447;
    p4_add_80448 <= p3_add_80448;
    p4_add_80449 <= p3_add_80449;
    p4_add_80450 <= p3_add_80450;
    p4_add_80451 <= p3_add_80451;
    p4_add_80452 <= p3_add_80452;
    p4_add_80453 <= p3_add_80453;
    p4_add_80454 <= p3_add_80454;
    p4_add_80455 <= p3_add_80455;
    p4_add_80456 <= p3_add_80456;
    p4_add_80457 <= p3_add_80457;
    p4_add_80458 <= p3_add_80458;
    p4_add_80459 <= p3_add_80459;
    p4_add_80460 <= p3_add_80460;
    p4_add_80461 <= p3_add_80461;
    p4_add_80462 <= p3_add_80462;
    p4_add_80463 <= p3_add_80463;
    p4_add_80464 <= p3_add_80464;
    p4_add_80465 <= p3_add_80465;
    p4_add_80466 <= p3_add_80466;
    p4_add_80467 <= p3_add_80467;
    p4_add_80468 <= p3_add_80468;
    p4_add_80469 <= p3_add_80469;
    p4_add_80470 <= p3_add_80470;
    p4_add_80471 <= p3_add_80471;
    p4_add_80472 <= p3_add_80472;
    p4_add_80473 <= p3_add_80473;
    p4_add_80474 <= p3_add_80474;
    p4_add_80475 <= p3_add_80475;
    p4_add_80476 <= p3_add_80476;
    p4_add_80477 <= p3_add_80477;
    p4_add_80478 <= p3_add_80478;
    p4_add_80479 <= p3_add_80479;
    p4_add_80480 <= p3_add_80480;
    p4_add_80481 <= p3_add_80481;
    p4_add_80482 <= p3_add_80482;
    p4_add_80483 <= p3_add_80483;
    p4_add_80484 <= p3_add_80484;
    p4_add_80485 <= p3_add_80485;
    p4_add_80486 <= p3_add_80486;
    p4_add_80487 <= p3_add_80487;
    p4_add_80488 <= p3_add_80488;
    p4_add_80489 <= p3_add_80489;
    p4_add_80490 <= p3_add_80490;
    p4_add_80491 <= p3_add_80491;
    p4_add_80492 <= p3_add_80492;
    p4_add_80493 <= p3_add_80493;
    p4_add_80494 <= p3_add_80494;
    p4_add_80495 <= p3_add_80495;
    p4_add_80496 <= p3_add_80496;
    p4_add_80497 <= p3_add_80497;
    p4_add_80498 <= p3_add_80498;
  end

  // ===== Pipe stage 5:
  wire [3499:0] p5_tuple_81325_comb;
  wire p5_tuple_index_81329_comb;
  wire p5_tuple_index_81332_comb;
  wire p5_tuple_index_81335_comb;
  wire p5_tuple_index_81338_comb;
  wire p5_tuple_index_81341_comb;
  wire p5_tuple_index_81344_comb;
  wire p5_tuple_index_81347_comb;
  wire p5_tuple_index_81350_comb;
  wire p5_tuple_index_81353_comb;
  wire p5_tuple_index_81356_comb;
  wire p5_tuple_index_81359_comb;
  wire p5_tuple_index_81362_comb;
  wire p5_tuple_index_81365_comb;
  wire p5_tuple_index_81368_comb;
  wire p5_tuple_index_81371_comb;
  wire p5_tuple_index_81374_comb;
  wire p5_tuple_index_81377_comb;
  wire p5_tuple_index_81380_comb;
  wire p5_tuple_index_81383_comb;
  wire p5_tuple_index_81386_comb;
  wire p5_tuple_index_81389_comb;
  wire p5_tuple_index_81392_comb;
  wire p5_tuple_index_81395_comb;
  wire p5_tuple_index_81398_comb;
  wire p5_tuple_index_81401_comb;
  wire p5_tuple_index_81404_comb;
  wire p5_tuple_index_81407_comb;
  wire p5_tuple_index_81410_comb;
  wire p5_tuple_index_81413_comb;
  wire p5_tuple_index_81416_comb;
  wire p5_tuple_index_81419_comb;
  wire p5_tuple_index_81422_comb;
  wire p5_tuple_index_81425_comb;
  wire p5_tuple_index_81428_comb;
  wire p5_tuple_index_81431_comb;
  wire p5_tuple_index_81434_comb;
  wire p5_tuple_index_81437_comb;
  wire p5_tuple_index_81440_comb;
  wire p5_tuple_index_81443_comb;
  wire p5_tuple_index_81446_comb;
  wire p5_tuple_index_81449_comb;
  wire p5_tuple_index_81452_comb;
  wire p5_tuple_index_81455_comb;
  wire p5_tuple_index_81458_comb;
  wire p5_tuple_index_81461_comb;
  wire p5_tuple_index_81464_comb;
  wire p5_tuple_index_81467_comb;
  wire p5_tuple_index_81470_comb;
  wire p5_tuple_index_81473_comb;
  wire p5_tuple_index_81476_comb;
  wire p5_tuple_index_81479_comb;
  wire p5_tuple_index_81482_comb;
  wire p5_tuple_index_81485_comb;
  wire p5_tuple_index_81488_comb;
  wire p5_tuple_index_81491_comb;
  wire p5_tuple_index_81494_comb;
  wire p5_tuple_index_81497_comb;
  wire p5_tuple_index_81500_comb;
  wire p5_tuple_index_81503_comb;
  wire p5_tuple_index_81506_comb;
  wire p5_tuple_index_81509_comb;
  wire p5_tuple_index_81512_comb;
  wire p5_tuple_index_81515_comb;
  wire p5_tuple_index_81518_comb;
  wire p5_tuple_index_81521_comb;
  wire p5_tuple_index_81524_comb;
  wire p5_tuple_index_81527_comb;
  wire p5_tuple_index_81530_comb;
  wire p5_tuple_index_81533_comb;
  wire p5_tuple_index_81536_comb;
  wire p5_tuple_index_81539_comb;
  wire p5_tuple_index_81542_comb;
  wire p5_tuple_index_81545_comb;
  wire p5_tuple_index_81548_comb;
  wire p5_tuple_index_81551_comb;
  wire p5_tuple_index_81554_comb;
  wire p5_tuple_index_81557_comb;
  wire p5_tuple_index_81560_comb;
  wire p5_tuple_index_81563_comb;
  wire p5_tuple_index_81566_comb;
  wire p5_tuple_index_81569_comb;
  wire p5_tuple_index_81572_comb;
  wire p5_tuple_index_81575_comb;
  wire p5_tuple_index_81578_comb;
  wire p5_tuple_index_81581_comb;
  wire p5_tuple_index_81584_comb;
  wire p5_tuple_index_81587_comb;
  wire p5_tuple_index_81590_comb;
  wire p5_tuple_index_81593_comb;
  wire p5_tuple_index_81596_comb;
  wire p5_tuple_index_81599_comb;
  wire p5_tuple_index_81602_comb;
  wire p5_tuple_index_81605_comb;
  wire p5_tuple_index_81608_comb;
  wire p5_tuple_index_81611_comb;
  wire p5_tuple_index_81614_comb;
  wire p5_tuple_index_81617_comb;
  wire p5_tuple_index_81620_comb;
  wire p5_tuple_index_81623_comb;
  wire p5_tuple_index_81626_comb;
  wire p5_tuple_index_81629_comb;
  wire p5_tuple_index_81632_comb;
  wire p5_tuple_index_81635_comb;
  wire p5_tuple_index_81638_comb;
  wire p5_tuple_index_81641_comb;
  wire p5_tuple_index_81644_comb;
  wire p5_tuple_index_81647_comb;
  wire p5_tuple_index_81650_comb;
  wire p5_tuple_index_81653_comb;
  wire p5_tuple_index_81656_comb;
  wire p5_tuple_index_81659_comb;
  wire p5_tuple_index_81662_comb;
  wire p5_tuple_index_81665_comb;
  wire p5_tuple_index_81668_comb;
  wire p5_tuple_index_81671_comb;
  wire p5_tuple_index_81674_comb;
  wire p5_tuple_index_81677_comb;
  wire p5_tuple_index_81680_comb;
  wire p5_tuple_index_81683_comb;
  wire p5_tuple_index_81686_comb;
  wire p5_tuple_index_81689_comb;
  wire p5_tuple_index_81692_comb;
  wire p5_tuple_index_81695_comb;
  wire p5_tuple_index_81698_comb;
  wire p5_tuple_index_81701_comb;
  wire p5_tuple_index_81704_comb;
  wire p5_tuple_index_81707_comb;
  wire p5_tuple_index_81710_comb;
  wire p5_tuple_index_81713_comb;
  wire p5_tuple_index_81716_comb;
  wire p5_tuple_index_81719_comb;
  wire p5_tuple_index_81722_comb;
  wire p5_tuple_index_81725_comb;
  wire p5_tuple_index_81728_comb;
  wire p5_tuple_index_81731_comb;
  wire p5_tuple_index_81734_comb;
  wire p5_tuple_index_81737_comb;
  wire p5_tuple_index_81740_comb;
  wire p5_tuple_index_81743_comb;
  wire p5_tuple_index_81746_comb;
  wire p5_tuple_index_81749_comb;
  wire p5_tuple_index_81752_comb;
  wire p5_tuple_index_81755_comb;
  wire p5_tuple_index_81758_comb;
  wire p5_tuple_index_81761_comb;
  wire p5_tuple_index_81764_comb;
  wire p5_tuple_index_81767_comb;
  wire p5_tuple_index_81770_comb;
  wire p5_tuple_index_81773_comb;
  wire p5_tuple_index_81776_comb;
  wire p5_tuple_index_81779_comb;
  wire p5_tuple_index_81782_comb;
  wire p5_tuple_index_81785_comb;
  wire p5_tuple_index_81788_comb;
  wire p5_tuple_index_81791_comb;
  wire p5_tuple_index_81794_comb;
  wire p5_tuple_index_81797_comb;
  wire p5_tuple_index_81800_comb;
  wire p5_tuple_index_81803_comb;
  wire p5_tuple_index_81806_comb;
  wire p5_tuple_index_81809_comb;
  wire p5_tuple_index_81812_comb;
  wire p5_tuple_index_81815_comb;
  wire p5_tuple_index_81818_comb;
  wire p5_tuple_index_81821_comb;
  wire p5_tuple_index_81824_comb;
  wire p5_tuple_index_81827_comb;
  wire p5_tuple_index_81830_comb;
  wire p5_tuple_index_81833_comb;
  wire p5_tuple_index_81836_comb;
  wire p5_tuple_index_81839_comb;
  wire p5_tuple_index_81842_comb;
  wire p5_tuple_index_81845_comb;
  wire p5_tuple_index_81848_comb;
  wire p5_tuple_index_81851_comb;
  wire p5_tuple_index_81854_comb;
  wire p5_tuple_index_81857_comb;
  wire p5_tuple_index_81860_comb;
  wire p5_tuple_index_81863_comb;
  wire p5_tuple_index_81866_comb;
  wire p5_tuple_index_81869_comb;
  wire p5_tuple_index_81872_comb;
  wire p5_tuple_index_81875_comb;
  wire p5_tuple_index_81878_comb;
  wire p5_tuple_index_81881_comb;
  wire p5_tuple_index_81884_comb;
  wire p5_tuple_index_81887_comb;
  wire p5_tuple_index_81890_comb;
  wire p5_tuple_index_81893_comb;
  wire p5_tuple_index_81896_comb;
  wire p5_tuple_index_81899_comb;
  wire p5_tuple_index_81902_comb;
  wire p5_tuple_index_81905_comb;
  wire p5_tuple_index_81908_comb;
  wire p5_tuple_index_81911_comb;
  wire p5_tuple_index_81914_comb;
  wire p5_tuple_index_81917_comb;
  wire p5_tuple_index_81920_comb;
  wire p5_tuple_index_81923_comb;
  wire p5_tuple_index_81926_comb;
  wire [32:0] p5_tuple_index_81929_comb;
  wire [32:0] p5_tuple_index_81932_comb;
  wire [32:0] p5_tuple_index_81935_comb;
  wire [32:0] p5_tuple_index_81938_comb;
  wire [32:0] p5_tuple_index_81941_comb;
  wire [32:0] p5_tuple_index_81944_comb;
  wire [32:0] p5_tuple_index_81947_comb;
  wire [32:0] p5_tuple_index_81950_comb;
  wire [32:0] p5_tuple_index_81953_comb;
  wire [32:0] p5_tuple_index_81956_comb;
  wire [32:0] p5_tuple_index_81959_comb;
  wire [32:0] p5_tuple_index_81962_comb;
  wire [32:0] p5_tuple_index_81965_comb;
  wire [32:0] p5_tuple_index_81968_comb;
  wire [32:0] p5_tuple_index_81971_comb;
  wire [32:0] p5_tuple_index_81974_comb;
  wire [32:0] p5_tuple_index_81977_comb;
  wire [32:0] p5_tuple_index_81980_comb;
  wire [32:0] p5_tuple_index_81983_comb;
  wire [32:0] p5_tuple_index_81986_comb;
  wire [32:0] p5_tuple_index_81989_comb;
  wire [32:0] p5_tuple_index_81992_comb;
  wire [32:0] p5_tuple_index_81995_comb;
  wire [32:0] p5_tuple_index_81998_comb;
  wire [32:0] p5_tuple_index_82001_comb;
  wire [32:0] p5_tuple_index_82004_comb;
  wire [32:0] p5_tuple_index_82007_comb;
  wire [32:0] p5_tuple_index_82010_comb;
  wire [32:0] p5_tuple_index_82013_comb;
  wire [32:0] p5_tuple_index_82016_comb;
  wire [32:0] p5_tuple_index_82019_comb;
  wire [32:0] p5_tuple_index_82022_comb;
  wire [32:0] p5_tuple_index_82025_comb;
  wire [32:0] p5_tuple_index_82028_comb;
  wire [32:0] p5_tuple_index_82031_comb;
  wire [32:0] p5_tuple_index_82034_comb;
  wire [32:0] p5_tuple_index_82037_comb;
  wire [32:0] p5_tuple_index_82040_comb;
  wire [32:0] p5_tuple_index_82043_comb;
  wire [32:0] p5_tuple_index_82046_comb;
  wire [32:0] p5_tuple_index_82049_comb;
  wire [32:0] p5_tuple_index_82052_comb;
  wire [32:0] p5_tuple_index_82055_comb;
  wire [32:0] p5_tuple_index_82058_comb;
  wire [32:0] p5_tuple_index_82061_comb;
  wire [32:0] p5_tuple_index_82064_comb;
  wire [32:0] p5_tuple_index_82067_comb;
  wire [32:0] p5_tuple_index_82070_comb;
  wire [32:0] p5_tuple_index_82073_comb;
  wire [32:0] p5_tuple_index_82076_comb;
  wire [32:0] p5_tuple_index_82079_comb;
  wire [32:0] p5_tuple_index_82082_comb;
  wire [32:0] p5_tuple_index_82085_comb;
  wire [32:0] p5_tuple_index_82088_comb;
  wire [32:0] p5_tuple_index_82091_comb;
  wire [32:0] p5_tuple_index_82094_comb;
  wire [32:0] p5_tuple_index_82097_comb;
  wire [32:0] p5_tuple_index_82100_comb;
  wire [32:0] p5_tuple_index_82103_comb;
  wire [32:0] p5_tuple_index_82106_comb;
  wire [32:0] p5_tuple_index_82109_comb;
  wire [32:0] p5_tuple_index_82112_comb;
  wire [32:0] p5_tuple_index_82115_comb;
  wire [32:0] p5_tuple_index_82118_comb;
  wire [32:0] p5_tuple_index_82121_comb;
  wire [32:0] p5_tuple_index_82124_comb;
  wire [32:0] p5_tuple_index_82127_comb;
  wire [32:0] p5_tuple_index_82130_comb;
  wire [32:0] p5_tuple_index_82133_comb;
  wire [32:0] p5_tuple_index_82136_comb;
  wire [32:0] p5_tuple_index_82139_comb;
  wire [32:0] p5_tuple_index_82142_comb;
  wire [32:0] p5_tuple_index_82145_comb;
  wire [32:0] p5_tuple_index_82148_comb;
  wire [32:0] p5_tuple_index_82151_comb;
  wire [32:0] p5_tuple_index_82154_comb;
  wire [32:0] p5_tuple_index_82157_comb;
  wire [32:0] p5_tuple_index_82160_comb;
  wire [32:0] p5_tuple_index_82163_comb;
  wire [32:0] p5_tuple_index_82166_comb;
  wire [32:0] p5_tuple_index_82169_comb;
  wire [32:0] p5_tuple_index_82172_comb;
  wire [32:0] p5_tuple_index_82175_comb;
  wire [32:0] p5_tuple_index_82178_comb;
  wire [32:0] p5_tuple_index_82181_comb;
  wire [32:0] p5_tuple_index_82184_comb;
  wire [32:0] p5_tuple_index_82187_comb;
  wire [32:0] p5_tuple_index_82190_comb;
  wire [32:0] p5_tuple_index_82193_comb;
  wire [32:0] p5_tuple_index_82196_comb;
  wire [32:0] p5_tuple_index_82199_comb;
  wire [32:0] p5_tuple_index_82202_comb;
  wire [32:0] p5_tuple_index_82205_comb;
  wire [32:0] p5_tuple_index_82208_comb;
  wire [32:0] p5_tuple_index_82211_comb;
  wire [32:0] p5_tuple_index_82214_comb;
  wire [32:0] p5_tuple_index_82217_comb;
  wire [32:0] p5_tuple_index_82220_comb;
  wire [32:0] p5_tuple_index_82223_comb;
  wire [32:0] p5_tuple_index_82226_comb;
  assign p5_tuple_81325_comb = {1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, 1'h1, {p4_add_80399, 1'h1}, {p4_add_80400, 1'h1}, {p4_add_80401, 1'h1}, {p4_add_80402, 1'h1}, {p4_add_80403, 1'h1}, {p4_add_80404, 1'h1}, {p4_add_80405, 1'h1}, {p4_add_80406, 1'h1}, {p4_add_80407, 1'h1}, {p4_add_80408, 1'h1}, {p4_add_80409, 1'h1}, {p4_add_80410, 1'h1}, {p4_add_80411, 1'h1}, {p4_add_80412, 1'h1}, {p4_add_80413, 1'h1}, {p4_add_80414, 1'h1}, {p4_add_80415, 1'h1}, {p4_add_80416, 1'h1}, {p4_add_80417, 1'h1}, {p4_add_80418, 1'h1}, {p4_add_80419, 1'h1}, {p4_add_80420, 1'h1}, {p4_add_80421, 1'h1}, {p4_add_80422, 1'h1}, {p4_add_80423, 1'h1}, {p4_add_80424, 1'h1}, {p4_add_80425, 1'h1}, {p4_add_80426, 1'h1}, {p4_add_80427, 1'h1}, {p4_add_80428, 1'h1}, {p4_add_80429, 1'h1}, {p4_add_80430, 1'h1}, {p4_add_80431, 1'h1}, {p4_add_80432, 1'h1}, {p4_add_80433, 1'h1}, {p4_add_80434, 1'h1}, {p4_add_80435, 1'h1}, {p4_add_80436, 1'h1}, {p4_add_80437, 1'h1}, {p4_add_80438, 1'h1}, {p4_add_80439, 1'h1}, {p4_add_80440, 1'h1}, {p4_add_80441, 1'h1}, {p4_add_80442, 1'h1}, {p4_add_80443, 1'h1}, {p4_add_80444, 1'h1}, {p4_add_80445, 1'h1}, {p4_add_80446, 1'h1}, {p4_add_80447, 1'h1}, {p4_add_80448, 1'h1}, {p4_add_80449, 1'h1}, {p4_add_80450, 1'h1}, {p4_add_80451, 1'h1}, {p4_add_80452, 1'h1}, {p4_add_80453, 1'h1}, {p4_add_80454, 1'h1}, {p4_add_80455, 1'h1}, {p4_add_80456, 1'h1}, {p4_add_80457, 1'h1}, {p4_add_80458, 1'h1}, {p4_add_80459, 1'h1}, {p4_add_80460, 1'h1}, {p4_add_80461, 1'h1}, {p4_add_80462, 1'h1}, {p4_add_80463, 1'h1}, {p4_add_80464, 1'h1}, {p4_add_80465, 1'h1}, {p4_add_80466, 1'h1}, {p4_add_80467, 1'h1}, {p4_add_80468, 1'h1}, {p4_add_80469, 1'h1}, {p4_add_80470, 1'h1}, {p4_add_80471, 1'h1}, {p4_add_80472, 1'h1}, {p4_add_80473, 1'h1}, {p4_add_80474, 1'h1}, {p4_add_80475, 1'h1}, {p4_add_80476, 1'h1}, {p4_add_80477, 1'h1}, {p4_add_80478, 1'h1}, {p4_add_80479, 1'h1}, {p4_add_80480, 1'h1}, {p4_add_80481, 1'h1}, {p4_add_80482, 1'h1}, {p4_add_80483, 1'h1}, {p4_add_80484, 1'h1}, {p4_add_80485, 1'h1}, {p4_add_80486, 1'h1}, {p4_add_80487, 1'h1}, {p4_add_80488, 1'h1}, {p4_add_80489, 1'h1}, {p4_add_80490, 1'h1}, {p4_add_80491, 1'h1}, {p4_add_80492, 1'h1}, {p4_add_80493, 1'h1}, {p4_add_80494, 1'h1}, {p4_add_80495, 1'h1}, {p4_add_80496, 1'h1}, {p4_add_80497, 1'h1}, {p4_add_80498, 1'h1}};
  assign p5_tuple_index_81329_comb = p5_tuple_81325_comb[3499:3499];
  assign p5_tuple_index_81332_comb = p5_tuple_81325_comb[3498:3498];
  assign p5_tuple_index_81335_comb = p5_tuple_81325_comb[3497:3497];
  assign p5_tuple_index_81338_comb = p5_tuple_81325_comb[3496:3496];
  assign p5_tuple_index_81341_comb = p5_tuple_81325_comb[3495:3495];
  assign p5_tuple_index_81344_comb = p5_tuple_81325_comb[3494:3494];
  assign p5_tuple_index_81347_comb = p5_tuple_81325_comb[3493:3493];
  assign p5_tuple_index_81350_comb = p5_tuple_81325_comb[3492:3492];
  assign p5_tuple_index_81353_comb = p5_tuple_81325_comb[3491:3491];
  assign p5_tuple_index_81356_comb = p5_tuple_81325_comb[3490:3490];
  assign p5_tuple_index_81359_comb = p5_tuple_81325_comb[3489:3489];
  assign p5_tuple_index_81362_comb = p5_tuple_81325_comb[3488:3488];
  assign p5_tuple_index_81365_comb = p5_tuple_81325_comb[3487:3487];
  assign p5_tuple_index_81368_comb = p5_tuple_81325_comb[3486:3486];
  assign p5_tuple_index_81371_comb = p5_tuple_81325_comb[3485:3485];
  assign p5_tuple_index_81374_comb = p5_tuple_81325_comb[3484:3484];
  assign p5_tuple_index_81377_comb = p5_tuple_81325_comb[3483:3483];
  assign p5_tuple_index_81380_comb = p5_tuple_81325_comb[3482:3482];
  assign p5_tuple_index_81383_comb = p5_tuple_81325_comb[3481:3481];
  assign p5_tuple_index_81386_comb = p5_tuple_81325_comb[3480:3480];
  assign p5_tuple_index_81389_comb = p5_tuple_81325_comb[3479:3479];
  assign p5_tuple_index_81392_comb = p5_tuple_81325_comb[3478:3478];
  assign p5_tuple_index_81395_comb = p5_tuple_81325_comb[3477:3477];
  assign p5_tuple_index_81398_comb = p5_tuple_81325_comb[3476:3476];
  assign p5_tuple_index_81401_comb = p5_tuple_81325_comb[3475:3475];
  assign p5_tuple_index_81404_comb = p5_tuple_81325_comb[3474:3474];
  assign p5_tuple_index_81407_comb = p5_tuple_81325_comb[3473:3473];
  assign p5_tuple_index_81410_comb = p5_tuple_81325_comb[3472:3472];
  assign p5_tuple_index_81413_comb = p5_tuple_81325_comb[3471:3471];
  assign p5_tuple_index_81416_comb = p5_tuple_81325_comb[3470:3470];
  assign p5_tuple_index_81419_comb = p5_tuple_81325_comb[3469:3469];
  assign p5_tuple_index_81422_comb = p5_tuple_81325_comb[3468:3468];
  assign p5_tuple_index_81425_comb = p5_tuple_81325_comb[3467:3467];
  assign p5_tuple_index_81428_comb = p5_tuple_81325_comb[3466:3466];
  assign p5_tuple_index_81431_comb = p5_tuple_81325_comb[3465:3465];
  assign p5_tuple_index_81434_comb = p5_tuple_81325_comb[3464:3464];
  assign p5_tuple_index_81437_comb = p5_tuple_81325_comb[3463:3463];
  assign p5_tuple_index_81440_comb = p5_tuple_81325_comb[3462:3462];
  assign p5_tuple_index_81443_comb = p5_tuple_81325_comb[3461:3461];
  assign p5_tuple_index_81446_comb = p5_tuple_81325_comb[3460:3460];
  assign p5_tuple_index_81449_comb = p5_tuple_81325_comb[3459:3459];
  assign p5_tuple_index_81452_comb = p5_tuple_81325_comb[3458:3458];
  assign p5_tuple_index_81455_comb = p5_tuple_81325_comb[3457:3457];
  assign p5_tuple_index_81458_comb = p5_tuple_81325_comb[3456:3456];
  assign p5_tuple_index_81461_comb = p5_tuple_81325_comb[3455:3455];
  assign p5_tuple_index_81464_comb = p5_tuple_81325_comb[3454:3454];
  assign p5_tuple_index_81467_comb = p5_tuple_81325_comb[3453:3453];
  assign p5_tuple_index_81470_comb = p5_tuple_81325_comb[3452:3452];
  assign p5_tuple_index_81473_comb = p5_tuple_81325_comb[3451:3451];
  assign p5_tuple_index_81476_comb = p5_tuple_81325_comb[3450:3450];
  assign p5_tuple_index_81479_comb = p5_tuple_81325_comb[3449:3449];
  assign p5_tuple_index_81482_comb = p5_tuple_81325_comb[3448:3448];
  assign p5_tuple_index_81485_comb = p5_tuple_81325_comb[3447:3447];
  assign p5_tuple_index_81488_comb = p5_tuple_81325_comb[3446:3446];
  assign p5_tuple_index_81491_comb = p5_tuple_81325_comb[3445:3445];
  assign p5_tuple_index_81494_comb = p5_tuple_81325_comb[3444:3444];
  assign p5_tuple_index_81497_comb = p5_tuple_81325_comb[3443:3443];
  assign p5_tuple_index_81500_comb = p5_tuple_81325_comb[3442:3442];
  assign p5_tuple_index_81503_comb = p5_tuple_81325_comb[3441:3441];
  assign p5_tuple_index_81506_comb = p5_tuple_81325_comb[3440:3440];
  assign p5_tuple_index_81509_comb = p5_tuple_81325_comb[3439:3439];
  assign p5_tuple_index_81512_comb = p5_tuple_81325_comb[3438:3438];
  assign p5_tuple_index_81515_comb = p5_tuple_81325_comb[3437:3437];
  assign p5_tuple_index_81518_comb = p5_tuple_81325_comb[3436:3436];
  assign p5_tuple_index_81521_comb = p5_tuple_81325_comb[3435:3435];
  assign p5_tuple_index_81524_comb = p5_tuple_81325_comb[3434:3434];
  assign p5_tuple_index_81527_comb = p5_tuple_81325_comb[3433:3433];
  assign p5_tuple_index_81530_comb = p5_tuple_81325_comb[3432:3432];
  assign p5_tuple_index_81533_comb = p5_tuple_81325_comb[3431:3431];
  assign p5_tuple_index_81536_comb = p5_tuple_81325_comb[3430:3430];
  assign p5_tuple_index_81539_comb = p5_tuple_81325_comb[3429:3429];
  assign p5_tuple_index_81542_comb = p5_tuple_81325_comb[3428:3428];
  assign p5_tuple_index_81545_comb = p5_tuple_81325_comb[3427:3427];
  assign p5_tuple_index_81548_comb = p5_tuple_81325_comb[3426:3426];
  assign p5_tuple_index_81551_comb = p5_tuple_81325_comb[3425:3425];
  assign p5_tuple_index_81554_comb = p5_tuple_81325_comb[3424:3424];
  assign p5_tuple_index_81557_comb = p5_tuple_81325_comb[3423:3423];
  assign p5_tuple_index_81560_comb = p5_tuple_81325_comb[3422:3422];
  assign p5_tuple_index_81563_comb = p5_tuple_81325_comb[3421:3421];
  assign p5_tuple_index_81566_comb = p5_tuple_81325_comb[3420:3420];
  assign p5_tuple_index_81569_comb = p5_tuple_81325_comb[3419:3419];
  assign p5_tuple_index_81572_comb = p5_tuple_81325_comb[3418:3418];
  assign p5_tuple_index_81575_comb = p5_tuple_81325_comb[3417:3417];
  assign p5_tuple_index_81578_comb = p5_tuple_81325_comb[3416:3416];
  assign p5_tuple_index_81581_comb = p5_tuple_81325_comb[3415:3415];
  assign p5_tuple_index_81584_comb = p5_tuple_81325_comb[3414:3414];
  assign p5_tuple_index_81587_comb = p5_tuple_81325_comb[3413:3413];
  assign p5_tuple_index_81590_comb = p5_tuple_81325_comb[3412:3412];
  assign p5_tuple_index_81593_comb = p5_tuple_81325_comb[3411:3411];
  assign p5_tuple_index_81596_comb = p5_tuple_81325_comb[3410:3410];
  assign p5_tuple_index_81599_comb = p5_tuple_81325_comb[3409:3409];
  assign p5_tuple_index_81602_comb = p5_tuple_81325_comb[3408:3408];
  assign p5_tuple_index_81605_comb = p5_tuple_81325_comb[3407:3407];
  assign p5_tuple_index_81608_comb = p5_tuple_81325_comb[3406:3406];
  assign p5_tuple_index_81611_comb = p5_tuple_81325_comb[3405:3405];
  assign p5_tuple_index_81614_comb = p5_tuple_81325_comb[3404:3404];
  assign p5_tuple_index_81617_comb = p5_tuple_81325_comb[3403:3403];
  assign p5_tuple_index_81620_comb = p5_tuple_81325_comb[3402:3402];
  assign p5_tuple_index_81623_comb = p5_tuple_81325_comb[3401:3401];
  assign p5_tuple_index_81626_comb = p5_tuple_81325_comb[3400:3400];
  assign p5_tuple_index_81629_comb = p5_tuple_81325_comb[3399:3399];
  assign p5_tuple_index_81632_comb = p5_tuple_81325_comb[3398:3398];
  assign p5_tuple_index_81635_comb = p5_tuple_81325_comb[3397:3397];
  assign p5_tuple_index_81638_comb = p5_tuple_81325_comb[3396:3396];
  assign p5_tuple_index_81641_comb = p5_tuple_81325_comb[3395:3395];
  assign p5_tuple_index_81644_comb = p5_tuple_81325_comb[3394:3394];
  assign p5_tuple_index_81647_comb = p5_tuple_81325_comb[3393:3393];
  assign p5_tuple_index_81650_comb = p5_tuple_81325_comb[3392:3392];
  assign p5_tuple_index_81653_comb = p5_tuple_81325_comb[3391:3391];
  assign p5_tuple_index_81656_comb = p5_tuple_81325_comb[3390:3390];
  assign p5_tuple_index_81659_comb = p5_tuple_81325_comb[3389:3389];
  assign p5_tuple_index_81662_comb = p5_tuple_81325_comb[3388:3388];
  assign p5_tuple_index_81665_comb = p5_tuple_81325_comb[3387:3387];
  assign p5_tuple_index_81668_comb = p5_tuple_81325_comb[3386:3386];
  assign p5_tuple_index_81671_comb = p5_tuple_81325_comb[3385:3385];
  assign p5_tuple_index_81674_comb = p5_tuple_81325_comb[3384:3384];
  assign p5_tuple_index_81677_comb = p5_tuple_81325_comb[3383:3383];
  assign p5_tuple_index_81680_comb = p5_tuple_81325_comb[3382:3382];
  assign p5_tuple_index_81683_comb = p5_tuple_81325_comb[3381:3381];
  assign p5_tuple_index_81686_comb = p5_tuple_81325_comb[3380:3380];
  assign p5_tuple_index_81689_comb = p5_tuple_81325_comb[3379:3379];
  assign p5_tuple_index_81692_comb = p5_tuple_81325_comb[3378:3378];
  assign p5_tuple_index_81695_comb = p5_tuple_81325_comb[3377:3377];
  assign p5_tuple_index_81698_comb = p5_tuple_81325_comb[3376:3376];
  assign p5_tuple_index_81701_comb = p5_tuple_81325_comb[3375:3375];
  assign p5_tuple_index_81704_comb = p5_tuple_81325_comb[3374:3374];
  assign p5_tuple_index_81707_comb = p5_tuple_81325_comb[3373:3373];
  assign p5_tuple_index_81710_comb = p5_tuple_81325_comb[3372:3372];
  assign p5_tuple_index_81713_comb = p5_tuple_81325_comb[3371:3371];
  assign p5_tuple_index_81716_comb = p5_tuple_81325_comb[3370:3370];
  assign p5_tuple_index_81719_comb = p5_tuple_81325_comb[3369:3369];
  assign p5_tuple_index_81722_comb = p5_tuple_81325_comb[3368:3368];
  assign p5_tuple_index_81725_comb = p5_tuple_81325_comb[3367:3367];
  assign p5_tuple_index_81728_comb = p5_tuple_81325_comb[3366:3366];
  assign p5_tuple_index_81731_comb = p5_tuple_81325_comb[3365:3365];
  assign p5_tuple_index_81734_comb = p5_tuple_81325_comb[3364:3364];
  assign p5_tuple_index_81737_comb = p5_tuple_81325_comb[3363:3363];
  assign p5_tuple_index_81740_comb = p5_tuple_81325_comb[3362:3362];
  assign p5_tuple_index_81743_comb = p5_tuple_81325_comb[3361:3361];
  assign p5_tuple_index_81746_comb = p5_tuple_81325_comb[3360:3360];
  assign p5_tuple_index_81749_comb = p5_tuple_81325_comb[3359:3359];
  assign p5_tuple_index_81752_comb = p5_tuple_81325_comb[3358:3358];
  assign p5_tuple_index_81755_comb = p5_tuple_81325_comb[3357:3357];
  assign p5_tuple_index_81758_comb = p5_tuple_81325_comb[3356:3356];
  assign p5_tuple_index_81761_comb = p5_tuple_81325_comb[3355:3355];
  assign p5_tuple_index_81764_comb = p5_tuple_81325_comb[3354:3354];
  assign p5_tuple_index_81767_comb = p5_tuple_81325_comb[3353:3353];
  assign p5_tuple_index_81770_comb = p5_tuple_81325_comb[3352:3352];
  assign p5_tuple_index_81773_comb = p5_tuple_81325_comb[3351:3351];
  assign p5_tuple_index_81776_comb = p5_tuple_81325_comb[3350:3350];
  assign p5_tuple_index_81779_comb = p5_tuple_81325_comb[3349:3349];
  assign p5_tuple_index_81782_comb = p5_tuple_81325_comb[3348:3348];
  assign p5_tuple_index_81785_comb = p5_tuple_81325_comb[3347:3347];
  assign p5_tuple_index_81788_comb = p5_tuple_81325_comb[3346:3346];
  assign p5_tuple_index_81791_comb = p5_tuple_81325_comb[3345:3345];
  assign p5_tuple_index_81794_comb = p5_tuple_81325_comb[3344:3344];
  assign p5_tuple_index_81797_comb = p5_tuple_81325_comb[3343:3343];
  assign p5_tuple_index_81800_comb = p5_tuple_81325_comb[3342:3342];
  assign p5_tuple_index_81803_comb = p5_tuple_81325_comb[3341:3341];
  assign p5_tuple_index_81806_comb = p5_tuple_81325_comb[3340:3340];
  assign p5_tuple_index_81809_comb = p5_tuple_81325_comb[3339:3339];
  assign p5_tuple_index_81812_comb = p5_tuple_81325_comb[3338:3338];
  assign p5_tuple_index_81815_comb = p5_tuple_81325_comb[3337:3337];
  assign p5_tuple_index_81818_comb = p5_tuple_81325_comb[3336:3336];
  assign p5_tuple_index_81821_comb = p5_tuple_81325_comb[3335:3335];
  assign p5_tuple_index_81824_comb = p5_tuple_81325_comb[3334:3334];
  assign p5_tuple_index_81827_comb = p5_tuple_81325_comb[3333:3333];
  assign p5_tuple_index_81830_comb = p5_tuple_81325_comb[3332:3332];
  assign p5_tuple_index_81833_comb = p5_tuple_81325_comb[3331:3331];
  assign p5_tuple_index_81836_comb = p5_tuple_81325_comb[3330:3330];
  assign p5_tuple_index_81839_comb = p5_tuple_81325_comb[3329:3329];
  assign p5_tuple_index_81842_comb = p5_tuple_81325_comb[3328:3328];
  assign p5_tuple_index_81845_comb = p5_tuple_81325_comb[3327:3327];
  assign p5_tuple_index_81848_comb = p5_tuple_81325_comb[3326:3326];
  assign p5_tuple_index_81851_comb = p5_tuple_81325_comb[3325:3325];
  assign p5_tuple_index_81854_comb = p5_tuple_81325_comb[3324:3324];
  assign p5_tuple_index_81857_comb = p5_tuple_81325_comb[3323:3323];
  assign p5_tuple_index_81860_comb = p5_tuple_81325_comb[3322:3322];
  assign p5_tuple_index_81863_comb = p5_tuple_81325_comb[3321:3321];
  assign p5_tuple_index_81866_comb = p5_tuple_81325_comb[3320:3320];
  assign p5_tuple_index_81869_comb = p5_tuple_81325_comb[3319:3319];
  assign p5_tuple_index_81872_comb = p5_tuple_81325_comb[3318:3318];
  assign p5_tuple_index_81875_comb = p5_tuple_81325_comb[3317:3317];
  assign p5_tuple_index_81878_comb = p5_tuple_81325_comb[3316:3316];
  assign p5_tuple_index_81881_comb = p5_tuple_81325_comb[3315:3315];
  assign p5_tuple_index_81884_comb = p5_tuple_81325_comb[3314:3314];
  assign p5_tuple_index_81887_comb = p5_tuple_81325_comb[3313:3313];
  assign p5_tuple_index_81890_comb = p5_tuple_81325_comb[3312:3312];
  assign p5_tuple_index_81893_comb = p5_tuple_81325_comb[3311:3311];
  assign p5_tuple_index_81896_comb = p5_tuple_81325_comb[3310:3310];
  assign p5_tuple_index_81899_comb = p5_tuple_81325_comb[3309:3309];
  assign p5_tuple_index_81902_comb = p5_tuple_81325_comb[3308:3308];
  assign p5_tuple_index_81905_comb = p5_tuple_81325_comb[3307:3307];
  assign p5_tuple_index_81908_comb = p5_tuple_81325_comb[3306:3306];
  assign p5_tuple_index_81911_comb = p5_tuple_81325_comb[3305:3305];
  assign p5_tuple_index_81914_comb = p5_tuple_81325_comb[3304:3304];
  assign p5_tuple_index_81917_comb = p5_tuple_81325_comb[3303:3303];
  assign p5_tuple_index_81920_comb = p5_tuple_81325_comb[3302:3302];
  assign p5_tuple_index_81923_comb = p5_tuple_81325_comb[3301:3301];
  assign p5_tuple_index_81926_comb = p5_tuple_81325_comb[3300:3300];
  assign p5_tuple_index_81929_comb = p5_tuple_81325_comb[3299:3267];
  assign p5_tuple_index_81932_comb = p5_tuple_81325_comb[3266:3234];
  assign p5_tuple_index_81935_comb = p5_tuple_81325_comb[3233:3201];
  assign p5_tuple_index_81938_comb = p5_tuple_81325_comb[3200:3168];
  assign p5_tuple_index_81941_comb = p5_tuple_81325_comb[3167:3135];
  assign p5_tuple_index_81944_comb = p5_tuple_81325_comb[3134:3102];
  assign p5_tuple_index_81947_comb = p5_tuple_81325_comb[3101:3069];
  assign p5_tuple_index_81950_comb = p5_tuple_81325_comb[3068:3036];
  assign p5_tuple_index_81953_comb = p5_tuple_81325_comb[3035:3003];
  assign p5_tuple_index_81956_comb = p5_tuple_81325_comb[3002:2970];
  assign p5_tuple_index_81959_comb = p5_tuple_81325_comb[2969:2937];
  assign p5_tuple_index_81962_comb = p5_tuple_81325_comb[2936:2904];
  assign p5_tuple_index_81965_comb = p5_tuple_81325_comb[2903:2871];
  assign p5_tuple_index_81968_comb = p5_tuple_81325_comb[2870:2838];
  assign p5_tuple_index_81971_comb = p5_tuple_81325_comb[2837:2805];
  assign p5_tuple_index_81974_comb = p5_tuple_81325_comb[2804:2772];
  assign p5_tuple_index_81977_comb = p5_tuple_81325_comb[2771:2739];
  assign p5_tuple_index_81980_comb = p5_tuple_81325_comb[2738:2706];
  assign p5_tuple_index_81983_comb = p5_tuple_81325_comb[2705:2673];
  assign p5_tuple_index_81986_comb = p5_tuple_81325_comb[2672:2640];
  assign p5_tuple_index_81989_comb = p5_tuple_81325_comb[2639:2607];
  assign p5_tuple_index_81992_comb = p5_tuple_81325_comb[2606:2574];
  assign p5_tuple_index_81995_comb = p5_tuple_81325_comb[2573:2541];
  assign p5_tuple_index_81998_comb = p5_tuple_81325_comb[2540:2508];
  assign p5_tuple_index_82001_comb = p5_tuple_81325_comb[2507:2475];
  assign p5_tuple_index_82004_comb = p5_tuple_81325_comb[2474:2442];
  assign p5_tuple_index_82007_comb = p5_tuple_81325_comb[2441:2409];
  assign p5_tuple_index_82010_comb = p5_tuple_81325_comb[2408:2376];
  assign p5_tuple_index_82013_comb = p5_tuple_81325_comb[2375:2343];
  assign p5_tuple_index_82016_comb = p5_tuple_81325_comb[2342:2310];
  assign p5_tuple_index_82019_comb = p5_tuple_81325_comb[2309:2277];
  assign p5_tuple_index_82022_comb = p5_tuple_81325_comb[2276:2244];
  assign p5_tuple_index_82025_comb = p5_tuple_81325_comb[2243:2211];
  assign p5_tuple_index_82028_comb = p5_tuple_81325_comb[2210:2178];
  assign p5_tuple_index_82031_comb = p5_tuple_81325_comb[2177:2145];
  assign p5_tuple_index_82034_comb = p5_tuple_81325_comb[2144:2112];
  assign p5_tuple_index_82037_comb = p5_tuple_81325_comb[2111:2079];
  assign p5_tuple_index_82040_comb = p5_tuple_81325_comb[2078:2046];
  assign p5_tuple_index_82043_comb = p5_tuple_81325_comb[2045:2013];
  assign p5_tuple_index_82046_comb = p5_tuple_81325_comb[2012:1980];
  assign p5_tuple_index_82049_comb = p5_tuple_81325_comb[1979:1947];
  assign p5_tuple_index_82052_comb = p5_tuple_81325_comb[1946:1914];
  assign p5_tuple_index_82055_comb = p5_tuple_81325_comb[1913:1881];
  assign p5_tuple_index_82058_comb = p5_tuple_81325_comb[1880:1848];
  assign p5_tuple_index_82061_comb = p5_tuple_81325_comb[1847:1815];
  assign p5_tuple_index_82064_comb = p5_tuple_81325_comb[1814:1782];
  assign p5_tuple_index_82067_comb = p5_tuple_81325_comb[1781:1749];
  assign p5_tuple_index_82070_comb = p5_tuple_81325_comb[1748:1716];
  assign p5_tuple_index_82073_comb = p5_tuple_81325_comb[1715:1683];
  assign p5_tuple_index_82076_comb = p5_tuple_81325_comb[1682:1650];
  assign p5_tuple_index_82079_comb = p5_tuple_81325_comb[1649:1617];
  assign p5_tuple_index_82082_comb = p5_tuple_81325_comb[1616:1584];
  assign p5_tuple_index_82085_comb = p5_tuple_81325_comb[1583:1551];
  assign p5_tuple_index_82088_comb = p5_tuple_81325_comb[1550:1518];
  assign p5_tuple_index_82091_comb = p5_tuple_81325_comb[1517:1485];
  assign p5_tuple_index_82094_comb = p5_tuple_81325_comb[1484:1452];
  assign p5_tuple_index_82097_comb = p5_tuple_81325_comb[1451:1419];
  assign p5_tuple_index_82100_comb = p5_tuple_81325_comb[1418:1386];
  assign p5_tuple_index_82103_comb = p5_tuple_81325_comb[1385:1353];
  assign p5_tuple_index_82106_comb = p5_tuple_81325_comb[1352:1320];
  assign p5_tuple_index_82109_comb = p5_tuple_81325_comb[1319:1287];
  assign p5_tuple_index_82112_comb = p5_tuple_81325_comb[1286:1254];
  assign p5_tuple_index_82115_comb = p5_tuple_81325_comb[1253:1221];
  assign p5_tuple_index_82118_comb = p5_tuple_81325_comb[1220:1188];
  assign p5_tuple_index_82121_comb = p5_tuple_81325_comb[1187:1155];
  assign p5_tuple_index_82124_comb = p5_tuple_81325_comb[1154:1122];
  assign p5_tuple_index_82127_comb = p5_tuple_81325_comb[1121:1089];
  assign p5_tuple_index_82130_comb = p5_tuple_81325_comb[1088:1056];
  assign p5_tuple_index_82133_comb = p5_tuple_81325_comb[1055:1023];
  assign p5_tuple_index_82136_comb = p5_tuple_81325_comb[1022:990];
  assign p5_tuple_index_82139_comb = p5_tuple_81325_comb[989:957];
  assign p5_tuple_index_82142_comb = p5_tuple_81325_comb[956:924];
  assign p5_tuple_index_82145_comb = p5_tuple_81325_comb[923:891];
  assign p5_tuple_index_82148_comb = p5_tuple_81325_comb[890:858];
  assign p5_tuple_index_82151_comb = p5_tuple_81325_comb[857:825];
  assign p5_tuple_index_82154_comb = p5_tuple_81325_comb[824:792];
  assign p5_tuple_index_82157_comb = p5_tuple_81325_comb[791:759];
  assign p5_tuple_index_82160_comb = p5_tuple_81325_comb[758:726];
  assign p5_tuple_index_82163_comb = p5_tuple_81325_comb[725:693];
  assign p5_tuple_index_82166_comb = p5_tuple_81325_comb[692:660];
  assign p5_tuple_index_82169_comb = p5_tuple_81325_comb[659:627];
  assign p5_tuple_index_82172_comb = p5_tuple_81325_comb[626:594];
  assign p5_tuple_index_82175_comb = p5_tuple_81325_comb[593:561];
  assign p5_tuple_index_82178_comb = p5_tuple_81325_comb[560:528];
  assign p5_tuple_index_82181_comb = p5_tuple_81325_comb[527:495];
  assign p5_tuple_index_82184_comb = p5_tuple_81325_comb[494:462];
  assign p5_tuple_index_82187_comb = p5_tuple_81325_comb[461:429];
  assign p5_tuple_index_82190_comb = p5_tuple_81325_comb[428:396];
  assign p5_tuple_index_82193_comb = p5_tuple_81325_comb[395:363];
  assign p5_tuple_index_82196_comb = p5_tuple_81325_comb[362:330];
  assign p5_tuple_index_82199_comb = p5_tuple_81325_comb[329:297];
  assign p5_tuple_index_82202_comb = p5_tuple_81325_comb[296:264];
  assign p5_tuple_index_82205_comb = p5_tuple_81325_comb[263:231];
  assign p5_tuple_index_82208_comb = p5_tuple_81325_comb[230:198];
  assign p5_tuple_index_82211_comb = p5_tuple_81325_comb[197:165];
  assign p5_tuple_index_82214_comb = p5_tuple_81325_comb[164:132];
  assign p5_tuple_index_82217_comb = p5_tuple_81325_comb[131:99];
  assign p5_tuple_index_82220_comb = p5_tuple_81325_comb[98:66];
  assign p5_tuple_index_82223_comb = p5_tuple_81325_comb[65:33];
  assign p5_tuple_index_82226_comb = p5_tuple_81325_comb[32:0];

  // Registers for pipe stage 5:
  reg p5_tuple_81325_index1;
  reg p5_tuple_81325_index2;
  reg p5_tuple_81325_index3;
  reg p5_tuple_81325_index4;
  reg p5_tuple_81325_index5;
  reg p5_tuple_81325_index6;
  reg p5_tuple_81325_index7;
  reg p5_tuple_81325_index8;
  reg p5_tuple_81325_index9;
  reg p5_tuple_81325_index10;
  reg p5_tuple_81325_index11;
  reg p5_tuple_81325_index12;
  reg p5_tuple_81325_index13;
  reg p5_tuple_81325_index14;
  reg p5_tuple_81325_index15;
  reg p5_tuple_81325_index16;
  reg p5_tuple_81325_index17;
  reg p5_tuple_81325_index18;
  reg p5_tuple_81325_index19;
  reg p5_tuple_81325_index20;
  reg p5_tuple_81325_index21;
  reg p5_tuple_81325_index22;
  reg p5_tuple_81325_index23;
  reg p5_tuple_81325_index24;
  reg p5_tuple_81325_index25;
  reg p5_tuple_81325_index26;
  reg p5_tuple_81325_index27;
  reg p5_tuple_81325_index28;
  reg p5_tuple_81325_index29;
  reg p5_tuple_81325_index30;
  reg p5_tuple_81325_index31;
  reg p5_tuple_81325_index32;
  reg p5_tuple_81325_index33;
  reg p5_tuple_81325_index34;
  reg p5_tuple_81325_index35;
  reg p5_tuple_81325_index36;
  reg p5_tuple_81325_index37;
  reg p5_tuple_81325_index38;
  reg p5_tuple_81325_index39;
  reg p5_tuple_81325_index40;
  reg p5_tuple_81325_index41;
  reg p5_tuple_81325_index42;
  reg p5_tuple_81325_index43;
  reg p5_tuple_81325_index44;
  reg p5_tuple_81325_index45;
  reg p5_tuple_81325_index46;
  reg p5_tuple_81325_index47;
  reg p5_tuple_81325_index48;
  reg p5_tuple_81325_index49;
  reg p5_tuple_81325_index50;
  reg p5_tuple_81325_index51;
  reg p5_tuple_81325_index52;
  reg p5_tuple_81325_index53;
  reg p5_tuple_81325_index54;
  reg p5_tuple_81325_index55;
  reg p5_tuple_81325_index56;
  reg p5_tuple_81325_index57;
  reg p5_tuple_81325_index58;
  reg p5_tuple_81325_index59;
  reg p5_tuple_81325_index60;
  reg p5_tuple_81325_index61;
  reg p5_tuple_81325_index62;
  reg p5_tuple_81325_index63;
  reg p5_tuple_81325_index64;
  reg p5_tuple_81325_index65;
  reg p5_tuple_81325_index66;
  reg p5_tuple_81325_index67;
  reg p5_tuple_81325_index68;
  reg p5_tuple_81325_index69;
  reg p5_tuple_81325_index70;
  reg p5_tuple_81325_index71;
  reg p5_tuple_81325_index72;
  reg p5_tuple_81325_index73;
  reg p5_tuple_81325_index74;
  reg p5_tuple_81325_index75;
  reg p5_tuple_81325_index76;
  reg p5_tuple_81325_index77;
  reg p5_tuple_81325_index78;
  reg p5_tuple_81325_index79;
  reg p5_tuple_81325_index80;
  reg p5_tuple_81325_index81;
  reg p5_tuple_81325_index82;
  reg p5_tuple_81325_index83;
  reg p5_tuple_81325_index84;
  reg p5_tuple_81325_index85;
  reg p5_tuple_81325_index86;
  reg p5_tuple_81325_index87;
  reg p5_tuple_81325_index88;
  reg p5_tuple_81325_index89;
  reg p5_tuple_81325_index90;
  reg p5_tuple_81325_index91;
  reg p5_tuple_81325_index92;
  reg p5_tuple_81325_index93;
  reg p5_tuple_81325_index94;
  reg p5_tuple_81325_index95;
  reg p5_tuple_81325_index96;
  reg p5_tuple_81325_index97;
  reg p5_tuple_81325_index98;
  reg p5_tuple_81325_index99;
  reg p5_tuple_81325_index100;
  reg p5_tuple_81325_index101;
  reg p5_tuple_81325_index102;
  reg p5_tuple_81325_index103;
  reg p5_tuple_81325_index104;
  reg p5_tuple_81325_index105;
  reg p5_tuple_81325_index106;
  reg p5_tuple_81325_index107;
  reg p5_tuple_81325_index108;
  reg p5_tuple_81325_index109;
  reg p5_tuple_81325_index110;
  reg p5_tuple_81325_index111;
  reg p5_tuple_81325_index112;
  reg p5_tuple_81325_index113;
  reg p5_tuple_81325_index114;
  reg p5_tuple_81325_index115;
  reg p5_tuple_81325_index116;
  reg p5_tuple_81325_index117;
  reg p5_tuple_81325_index118;
  reg p5_tuple_81325_index119;
  reg p5_tuple_81325_index120;
  reg p5_tuple_81325_index121;
  reg p5_tuple_81325_index122;
  reg p5_tuple_81325_index123;
  reg p5_tuple_81325_index124;
  reg p5_tuple_81325_index125;
  reg p5_tuple_81325_index126;
  reg p5_tuple_81325_index127;
  reg p5_tuple_81325_index128;
  reg p5_tuple_81325_index129;
  reg p5_tuple_81325_index130;
  reg p5_tuple_81325_index131;
  reg p5_tuple_81325_index132;
  reg p5_tuple_81325_index133;
  reg p5_tuple_81325_index134;
  reg p5_tuple_81325_index135;
  reg p5_tuple_81325_index136;
  reg p5_tuple_81325_index137;
  reg p5_tuple_81325_index138;
  reg p5_tuple_81325_index139;
  reg p5_tuple_81325_index140;
  reg p5_tuple_81325_index141;
  reg p5_tuple_81325_index142;
  reg p5_tuple_81325_index143;
  reg p5_tuple_81325_index144;
  reg p5_tuple_81325_index145;
  reg p5_tuple_81325_index146;
  reg p5_tuple_81325_index147;
  reg p5_tuple_81325_index148;
  reg p5_tuple_81325_index149;
  reg p5_tuple_81325_index150;
  reg p5_tuple_81325_index151;
  reg p5_tuple_81325_index152;
  reg p5_tuple_81325_index153;
  reg p5_tuple_81325_index154;
  reg p5_tuple_81325_index155;
  reg p5_tuple_81325_index156;
  reg p5_tuple_81325_index157;
  reg p5_tuple_81325_index158;
  reg p5_tuple_81325_index159;
  reg p5_tuple_81325_index160;
  reg p5_tuple_81325_index161;
  reg p5_tuple_81325_index162;
  reg p5_tuple_81325_index163;
  reg p5_tuple_81325_index164;
  reg p5_tuple_81325_index165;
  reg p5_tuple_81325_index166;
  reg p5_tuple_81325_index167;
  reg p5_tuple_81325_index168;
  reg p5_tuple_81325_index169;
  reg p5_tuple_81325_index170;
  reg p5_tuple_81325_index171;
  reg p5_tuple_81325_index172;
  reg p5_tuple_81325_index173;
  reg p5_tuple_81325_index174;
  reg p5_tuple_81325_index175;
  reg p5_tuple_81325_index176;
  reg p5_tuple_81325_index177;
  reg p5_tuple_81325_index178;
  reg p5_tuple_81325_index179;
  reg p5_tuple_81325_index180;
  reg p5_tuple_81325_index181;
  reg p5_tuple_81325_index182;
  reg p5_tuple_81325_index183;
  reg p5_tuple_81325_index184;
  reg p5_tuple_81325_index185;
  reg p5_tuple_81325_index186;
  reg p5_tuple_81325_index187;
  reg p5_tuple_81325_index188;
  reg p5_tuple_81325_index189;
  reg p5_tuple_81325_index190;
  reg p5_tuple_81325_index191;
  reg p5_tuple_81325_index192;
  reg p5_tuple_81325_index193;
  reg p5_tuple_81325_index194;
  reg p5_tuple_81325_index195;
  reg p5_tuple_81325_index196;
  reg p5_tuple_81325_index197;
  reg p5_tuple_81325_index198;
  reg p5_tuple_81325_index199;
  reg p5_tuple_81325_index200;
  reg [32:0] p5_tuple_81325_index201;
  reg [32:0] p5_tuple_81325_index202;
  reg [32:0] p5_tuple_81325_index203;
  reg [32:0] p5_tuple_81325_index204;
  reg [32:0] p5_tuple_81325_index205;
  reg [32:0] p5_tuple_81325_index206;
  reg [32:0] p5_tuple_81325_index207;
  reg [32:0] p5_tuple_81325_index208;
  reg [32:0] p5_tuple_81325_index209;
  reg [32:0] p5_tuple_81325_index210;
  reg [32:0] p5_tuple_81325_index211;
  reg [32:0] p5_tuple_81325_index212;
  reg [32:0] p5_tuple_81325_index213;
  reg [32:0] p5_tuple_81325_index214;
  reg [32:0] p5_tuple_81325_index215;
  reg [32:0] p5_tuple_81325_index216;
  reg [32:0] p5_tuple_81325_index217;
  reg [32:0] p5_tuple_81325_index218;
  reg [32:0] p5_tuple_81325_index219;
  reg [32:0] p5_tuple_81325_index220;
  reg [32:0] p5_tuple_81325_index221;
  reg [32:0] p5_tuple_81325_index222;
  reg [32:0] p5_tuple_81325_index223;
  reg [32:0] p5_tuple_81325_index224;
  reg [32:0] p5_tuple_81325_index225;
  reg [32:0] p5_tuple_81325_index226;
  reg [32:0] p5_tuple_81325_index227;
  reg [32:0] p5_tuple_81325_index228;
  reg [32:0] p5_tuple_81325_index229;
  reg [32:0] p5_tuple_81325_index230;
  reg [32:0] p5_tuple_81325_index231;
  reg [32:0] p5_tuple_81325_index232;
  reg [32:0] p5_tuple_81325_index233;
  reg [32:0] p5_tuple_81325_index234;
  reg [32:0] p5_tuple_81325_index235;
  reg [32:0] p5_tuple_81325_index236;
  reg [32:0] p5_tuple_81325_index237;
  reg [32:0] p5_tuple_81325_index238;
  reg [32:0] p5_tuple_81325_index239;
  reg [32:0] p5_tuple_81325_index240;
  reg [32:0] p5_tuple_81325_index241;
  reg [32:0] p5_tuple_81325_index242;
  reg [32:0] p5_tuple_81325_index243;
  reg [32:0] p5_tuple_81325_index244;
  reg [32:0] p5_tuple_81325_index245;
  reg [32:0] p5_tuple_81325_index246;
  reg [32:0] p5_tuple_81325_index247;
  reg [32:0] p5_tuple_81325_index248;
  reg [32:0] p5_tuple_81325_index249;
  reg [32:0] p5_tuple_81325_index250;
  reg [32:0] p5_tuple_81325_index251;
  reg [32:0] p5_tuple_81325_index252;
  reg [32:0] p5_tuple_81325_index253;
  reg [32:0] p5_tuple_81325_index254;
  reg [32:0] p5_tuple_81325_index255;
  reg [32:0] p5_tuple_81325_index256;
  reg [32:0] p5_tuple_81325_index257;
  reg [32:0] p5_tuple_81325_index258;
  reg [32:0] p5_tuple_81325_index259;
  reg [32:0] p5_tuple_81325_index260;
  reg [32:0] p5_tuple_81325_index261;
  reg [32:0] p5_tuple_81325_index262;
  reg [32:0] p5_tuple_81325_index263;
  reg [32:0] p5_tuple_81325_index264;
  reg [32:0] p5_tuple_81325_index265;
  reg [32:0] p5_tuple_81325_index266;
  reg [32:0] p5_tuple_81325_index267;
  reg [32:0] p5_tuple_81325_index268;
  reg [32:0] p5_tuple_81325_index269;
  reg [32:0] p5_tuple_81325_index270;
  reg [32:0] p5_tuple_81325_index271;
  reg [32:0] p5_tuple_81325_index272;
  reg [32:0] p5_tuple_81325_index273;
  reg [32:0] p5_tuple_81325_index274;
  reg [32:0] p5_tuple_81325_index275;
  reg [32:0] p5_tuple_81325_index276;
  reg [32:0] p5_tuple_81325_index277;
  reg [32:0] p5_tuple_81325_index278;
  reg [32:0] p5_tuple_81325_index279;
  reg [32:0] p5_tuple_81325_index280;
  reg [32:0] p5_tuple_81325_index281;
  reg [32:0] p5_tuple_81325_index282;
  reg [32:0] p5_tuple_81325_index283;
  reg [32:0] p5_tuple_81325_index284;
  reg [32:0] p5_tuple_81325_index285;
  reg [32:0] p5_tuple_81325_index286;
  reg [32:0] p5_tuple_81325_index287;
  reg [32:0] p5_tuple_81325_index288;
  reg [32:0] p5_tuple_81325_index289;
  reg [32:0] p5_tuple_81325_index290;
  reg [32:0] p5_tuple_81325_index291;
  reg [32:0] p5_tuple_81325_index292;
  reg [32:0] p5_tuple_81325_index293;
  reg [32:0] p5_tuple_81325_index294;
  reg [32:0] p5_tuple_81325_index295;
  reg [32:0] p5_tuple_81325_index296;
  reg [32:0] p5_tuple_81325_index297;
  reg [32:0] p5_tuple_81325_index298;
  reg [32:0] p5_tuple_81325_index299;
  reg [32:0] p5_tuple_81325_index300;
  always_ff @ (posedge clk) begin
    p5_tuple_81325_index1 <= p5_tuple_index_81329_comb;
    p5_tuple_81325_index2 <= p5_tuple_index_81332_comb;
    p5_tuple_81325_index3 <= p5_tuple_index_81335_comb;
    p5_tuple_81325_index4 <= p5_tuple_index_81338_comb;
    p5_tuple_81325_index5 <= p5_tuple_index_81341_comb;
    p5_tuple_81325_index6 <= p5_tuple_index_81344_comb;
    p5_tuple_81325_index7 <= p5_tuple_index_81347_comb;
    p5_tuple_81325_index8 <= p5_tuple_index_81350_comb;
    p5_tuple_81325_index9 <= p5_tuple_index_81353_comb;
    p5_tuple_81325_index10 <= p5_tuple_index_81356_comb;
    p5_tuple_81325_index11 <= p5_tuple_index_81359_comb;
    p5_tuple_81325_index12 <= p5_tuple_index_81362_comb;
    p5_tuple_81325_index13 <= p5_tuple_index_81365_comb;
    p5_tuple_81325_index14 <= p5_tuple_index_81368_comb;
    p5_tuple_81325_index15 <= p5_tuple_index_81371_comb;
    p5_tuple_81325_index16 <= p5_tuple_index_81374_comb;
    p5_tuple_81325_index17 <= p5_tuple_index_81377_comb;
    p5_tuple_81325_index18 <= p5_tuple_index_81380_comb;
    p5_tuple_81325_index19 <= p5_tuple_index_81383_comb;
    p5_tuple_81325_index20 <= p5_tuple_index_81386_comb;
    p5_tuple_81325_index21 <= p5_tuple_index_81389_comb;
    p5_tuple_81325_index22 <= p5_tuple_index_81392_comb;
    p5_tuple_81325_index23 <= p5_tuple_index_81395_comb;
    p5_tuple_81325_index24 <= p5_tuple_index_81398_comb;
    p5_tuple_81325_index25 <= p5_tuple_index_81401_comb;
    p5_tuple_81325_index26 <= p5_tuple_index_81404_comb;
    p5_tuple_81325_index27 <= p5_tuple_index_81407_comb;
    p5_tuple_81325_index28 <= p5_tuple_index_81410_comb;
    p5_tuple_81325_index29 <= p5_tuple_index_81413_comb;
    p5_tuple_81325_index30 <= p5_tuple_index_81416_comb;
    p5_tuple_81325_index31 <= p5_tuple_index_81419_comb;
    p5_tuple_81325_index32 <= p5_tuple_index_81422_comb;
    p5_tuple_81325_index33 <= p5_tuple_index_81425_comb;
    p5_tuple_81325_index34 <= p5_tuple_index_81428_comb;
    p5_tuple_81325_index35 <= p5_tuple_index_81431_comb;
    p5_tuple_81325_index36 <= p5_tuple_index_81434_comb;
    p5_tuple_81325_index37 <= p5_tuple_index_81437_comb;
    p5_tuple_81325_index38 <= p5_tuple_index_81440_comb;
    p5_tuple_81325_index39 <= p5_tuple_index_81443_comb;
    p5_tuple_81325_index40 <= p5_tuple_index_81446_comb;
    p5_tuple_81325_index41 <= p5_tuple_index_81449_comb;
    p5_tuple_81325_index42 <= p5_tuple_index_81452_comb;
    p5_tuple_81325_index43 <= p5_tuple_index_81455_comb;
    p5_tuple_81325_index44 <= p5_tuple_index_81458_comb;
    p5_tuple_81325_index45 <= p5_tuple_index_81461_comb;
    p5_tuple_81325_index46 <= p5_tuple_index_81464_comb;
    p5_tuple_81325_index47 <= p5_tuple_index_81467_comb;
    p5_tuple_81325_index48 <= p5_tuple_index_81470_comb;
    p5_tuple_81325_index49 <= p5_tuple_index_81473_comb;
    p5_tuple_81325_index50 <= p5_tuple_index_81476_comb;
    p5_tuple_81325_index51 <= p5_tuple_index_81479_comb;
    p5_tuple_81325_index52 <= p5_tuple_index_81482_comb;
    p5_tuple_81325_index53 <= p5_tuple_index_81485_comb;
    p5_tuple_81325_index54 <= p5_tuple_index_81488_comb;
    p5_tuple_81325_index55 <= p5_tuple_index_81491_comb;
    p5_tuple_81325_index56 <= p5_tuple_index_81494_comb;
    p5_tuple_81325_index57 <= p5_tuple_index_81497_comb;
    p5_tuple_81325_index58 <= p5_tuple_index_81500_comb;
    p5_tuple_81325_index59 <= p5_tuple_index_81503_comb;
    p5_tuple_81325_index60 <= p5_tuple_index_81506_comb;
    p5_tuple_81325_index61 <= p5_tuple_index_81509_comb;
    p5_tuple_81325_index62 <= p5_tuple_index_81512_comb;
    p5_tuple_81325_index63 <= p5_tuple_index_81515_comb;
    p5_tuple_81325_index64 <= p5_tuple_index_81518_comb;
    p5_tuple_81325_index65 <= p5_tuple_index_81521_comb;
    p5_tuple_81325_index66 <= p5_tuple_index_81524_comb;
    p5_tuple_81325_index67 <= p5_tuple_index_81527_comb;
    p5_tuple_81325_index68 <= p5_tuple_index_81530_comb;
    p5_tuple_81325_index69 <= p5_tuple_index_81533_comb;
    p5_tuple_81325_index70 <= p5_tuple_index_81536_comb;
    p5_tuple_81325_index71 <= p5_tuple_index_81539_comb;
    p5_tuple_81325_index72 <= p5_tuple_index_81542_comb;
    p5_tuple_81325_index73 <= p5_tuple_index_81545_comb;
    p5_tuple_81325_index74 <= p5_tuple_index_81548_comb;
    p5_tuple_81325_index75 <= p5_tuple_index_81551_comb;
    p5_tuple_81325_index76 <= p5_tuple_index_81554_comb;
    p5_tuple_81325_index77 <= p5_tuple_index_81557_comb;
    p5_tuple_81325_index78 <= p5_tuple_index_81560_comb;
    p5_tuple_81325_index79 <= p5_tuple_index_81563_comb;
    p5_tuple_81325_index80 <= p5_tuple_index_81566_comb;
    p5_tuple_81325_index81 <= p5_tuple_index_81569_comb;
    p5_tuple_81325_index82 <= p5_tuple_index_81572_comb;
    p5_tuple_81325_index83 <= p5_tuple_index_81575_comb;
    p5_tuple_81325_index84 <= p5_tuple_index_81578_comb;
    p5_tuple_81325_index85 <= p5_tuple_index_81581_comb;
    p5_tuple_81325_index86 <= p5_tuple_index_81584_comb;
    p5_tuple_81325_index87 <= p5_tuple_index_81587_comb;
    p5_tuple_81325_index88 <= p5_tuple_index_81590_comb;
    p5_tuple_81325_index89 <= p5_tuple_index_81593_comb;
    p5_tuple_81325_index90 <= p5_tuple_index_81596_comb;
    p5_tuple_81325_index91 <= p5_tuple_index_81599_comb;
    p5_tuple_81325_index92 <= p5_tuple_index_81602_comb;
    p5_tuple_81325_index93 <= p5_tuple_index_81605_comb;
    p5_tuple_81325_index94 <= p5_tuple_index_81608_comb;
    p5_tuple_81325_index95 <= p5_tuple_index_81611_comb;
    p5_tuple_81325_index96 <= p5_tuple_index_81614_comb;
    p5_tuple_81325_index97 <= p5_tuple_index_81617_comb;
    p5_tuple_81325_index98 <= p5_tuple_index_81620_comb;
    p5_tuple_81325_index99 <= p5_tuple_index_81623_comb;
    p5_tuple_81325_index100 <= p5_tuple_index_81626_comb;
    p5_tuple_81325_index101 <= p5_tuple_index_81629_comb;
    p5_tuple_81325_index102 <= p5_tuple_index_81632_comb;
    p5_tuple_81325_index103 <= p5_tuple_index_81635_comb;
    p5_tuple_81325_index104 <= p5_tuple_index_81638_comb;
    p5_tuple_81325_index105 <= p5_tuple_index_81641_comb;
    p5_tuple_81325_index106 <= p5_tuple_index_81644_comb;
    p5_tuple_81325_index107 <= p5_tuple_index_81647_comb;
    p5_tuple_81325_index108 <= p5_tuple_index_81650_comb;
    p5_tuple_81325_index109 <= p5_tuple_index_81653_comb;
    p5_tuple_81325_index110 <= p5_tuple_index_81656_comb;
    p5_tuple_81325_index111 <= p5_tuple_index_81659_comb;
    p5_tuple_81325_index112 <= p5_tuple_index_81662_comb;
    p5_tuple_81325_index113 <= p5_tuple_index_81665_comb;
    p5_tuple_81325_index114 <= p5_tuple_index_81668_comb;
    p5_tuple_81325_index115 <= p5_tuple_index_81671_comb;
    p5_tuple_81325_index116 <= p5_tuple_index_81674_comb;
    p5_tuple_81325_index117 <= p5_tuple_index_81677_comb;
    p5_tuple_81325_index118 <= p5_tuple_index_81680_comb;
    p5_tuple_81325_index119 <= p5_tuple_index_81683_comb;
    p5_tuple_81325_index120 <= p5_tuple_index_81686_comb;
    p5_tuple_81325_index121 <= p5_tuple_index_81689_comb;
    p5_tuple_81325_index122 <= p5_tuple_index_81692_comb;
    p5_tuple_81325_index123 <= p5_tuple_index_81695_comb;
    p5_tuple_81325_index124 <= p5_tuple_index_81698_comb;
    p5_tuple_81325_index125 <= p5_tuple_index_81701_comb;
    p5_tuple_81325_index126 <= p5_tuple_index_81704_comb;
    p5_tuple_81325_index127 <= p5_tuple_index_81707_comb;
    p5_tuple_81325_index128 <= p5_tuple_index_81710_comb;
    p5_tuple_81325_index129 <= p5_tuple_index_81713_comb;
    p5_tuple_81325_index130 <= p5_tuple_index_81716_comb;
    p5_tuple_81325_index131 <= p5_tuple_index_81719_comb;
    p5_tuple_81325_index132 <= p5_tuple_index_81722_comb;
    p5_tuple_81325_index133 <= p5_tuple_index_81725_comb;
    p5_tuple_81325_index134 <= p5_tuple_index_81728_comb;
    p5_tuple_81325_index135 <= p5_tuple_index_81731_comb;
    p5_tuple_81325_index136 <= p5_tuple_index_81734_comb;
    p5_tuple_81325_index137 <= p5_tuple_index_81737_comb;
    p5_tuple_81325_index138 <= p5_tuple_index_81740_comb;
    p5_tuple_81325_index139 <= p5_tuple_index_81743_comb;
    p5_tuple_81325_index140 <= p5_tuple_index_81746_comb;
    p5_tuple_81325_index141 <= p5_tuple_index_81749_comb;
    p5_tuple_81325_index142 <= p5_tuple_index_81752_comb;
    p5_tuple_81325_index143 <= p5_tuple_index_81755_comb;
    p5_tuple_81325_index144 <= p5_tuple_index_81758_comb;
    p5_tuple_81325_index145 <= p5_tuple_index_81761_comb;
    p5_tuple_81325_index146 <= p5_tuple_index_81764_comb;
    p5_tuple_81325_index147 <= p5_tuple_index_81767_comb;
    p5_tuple_81325_index148 <= p5_tuple_index_81770_comb;
    p5_tuple_81325_index149 <= p5_tuple_index_81773_comb;
    p5_tuple_81325_index150 <= p5_tuple_index_81776_comb;
    p5_tuple_81325_index151 <= p5_tuple_index_81779_comb;
    p5_tuple_81325_index152 <= p5_tuple_index_81782_comb;
    p5_tuple_81325_index153 <= p5_tuple_index_81785_comb;
    p5_tuple_81325_index154 <= p5_tuple_index_81788_comb;
    p5_tuple_81325_index155 <= p5_tuple_index_81791_comb;
    p5_tuple_81325_index156 <= p5_tuple_index_81794_comb;
    p5_tuple_81325_index157 <= p5_tuple_index_81797_comb;
    p5_tuple_81325_index158 <= p5_tuple_index_81800_comb;
    p5_tuple_81325_index159 <= p5_tuple_index_81803_comb;
    p5_tuple_81325_index160 <= p5_tuple_index_81806_comb;
    p5_tuple_81325_index161 <= p5_tuple_index_81809_comb;
    p5_tuple_81325_index162 <= p5_tuple_index_81812_comb;
    p5_tuple_81325_index163 <= p5_tuple_index_81815_comb;
    p5_tuple_81325_index164 <= p5_tuple_index_81818_comb;
    p5_tuple_81325_index165 <= p5_tuple_index_81821_comb;
    p5_tuple_81325_index166 <= p5_tuple_index_81824_comb;
    p5_tuple_81325_index167 <= p5_tuple_index_81827_comb;
    p5_tuple_81325_index168 <= p5_tuple_index_81830_comb;
    p5_tuple_81325_index169 <= p5_tuple_index_81833_comb;
    p5_tuple_81325_index170 <= p5_tuple_index_81836_comb;
    p5_tuple_81325_index171 <= p5_tuple_index_81839_comb;
    p5_tuple_81325_index172 <= p5_tuple_index_81842_comb;
    p5_tuple_81325_index173 <= p5_tuple_index_81845_comb;
    p5_tuple_81325_index174 <= p5_tuple_index_81848_comb;
    p5_tuple_81325_index175 <= p5_tuple_index_81851_comb;
    p5_tuple_81325_index176 <= p5_tuple_index_81854_comb;
    p5_tuple_81325_index177 <= p5_tuple_index_81857_comb;
    p5_tuple_81325_index178 <= p5_tuple_index_81860_comb;
    p5_tuple_81325_index179 <= p5_tuple_index_81863_comb;
    p5_tuple_81325_index180 <= p5_tuple_index_81866_comb;
    p5_tuple_81325_index181 <= p5_tuple_index_81869_comb;
    p5_tuple_81325_index182 <= p5_tuple_index_81872_comb;
    p5_tuple_81325_index183 <= p5_tuple_index_81875_comb;
    p5_tuple_81325_index184 <= p5_tuple_index_81878_comb;
    p5_tuple_81325_index185 <= p5_tuple_index_81881_comb;
    p5_tuple_81325_index186 <= p5_tuple_index_81884_comb;
    p5_tuple_81325_index187 <= p5_tuple_index_81887_comb;
    p5_tuple_81325_index188 <= p5_tuple_index_81890_comb;
    p5_tuple_81325_index189 <= p5_tuple_index_81893_comb;
    p5_tuple_81325_index190 <= p5_tuple_index_81896_comb;
    p5_tuple_81325_index191 <= p5_tuple_index_81899_comb;
    p5_tuple_81325_index192 <= p5_tuple_index_81902_comb;
    p5_tuple_81325_index193 <= p5_tuple_index_81905_comb;
    p5_tuple_81325_index194 <= p5_tuple_index_81908_comb;
    p5_tuple_81325_index195 <= p5_tuple_index_81911_comb;
    p5_tuple_81325_index196 <= p5_tuple_index_81914_comb;
    p5_tuple_81325_index197 <= p5_tuple_index_81917_comb;
    p5_tuple_81325_index198 <= p5_tuple_index_81920_comb;
    p5_tuple_81325_index199 <= p5_tuple_index_81923_comb;
    p5_tuple_81325_index200 <= p5_tuple_index_81926_comb;
    p5_tuple_81325_index201 <= p5_tuple_index_81929_comb;
    p5_tuple_81325_index202 <= p5_tuple_index_81932_comb;
    p5_tuple_81325_index203 <= p5_tuple_index_81935_comb;
    p5_tuple_81325_index204 <= p5_tuple_index_81938_comb;
    p5_tuple_81325_index205 <= p5_tuple_index_81941_comb;
    p5_tuple_81325_index206 <= p5_tuple_index_81944_comb;
    p5_tuple_81325_index207 <= p5_tuple_index_81947_comb;
    p5_tuple_81325_index208 <= p5_tuple_index_81950_comb;
    p5_tuple_81325_index209 <= p5_tuple_index_81953_comb;
    p5_tuple_81325_index210 <= p5_tuple_index_81956_comb;
    p5_tuple_81325_index211 <= p5_tuple_index_81959_comb;
    p5_tuple_81325_index212 <= p5_tuple_index_81962_comb;
    p5_tuple_81325_index213 <= p5_tuple_index_81965_comb;
    p5_tuple_81325_index214 <= p5_tuple_index_81968_comb;
    p5_tuple_81325_index215 <= p5_tuple_index_81971_comb;
    p5_tuple_81325_index216 <= p5_tuple_index_81974_comb;
    p5_tuple_81325_index217 <= p5_tuple_index_81977_comb;
    p5_tuple_81325_index218 <= p5_tuple_index_81980_comb;
    p5_tuple_81325_index219 <= p5_tuple_index_81983_comb;
    p5_tuple_81325_index220 <= p5_tuple_index_81986_comb;
    p5_tuple_81325_index221 <= p5_tuple_index_81989_comb;
    p5_tuple_81325_index222 <= p5_tuple_index_81992_comb;
    p5_tuple_81325_index223 <= p5_tuple_index_81995_comb;
    p5_tuple_81325_index224 <= p5_tuple_index_81998_comb;
    p5_tuple_81325_index225 <= p5_tuple_index_82001_comb;
    p5_tuple_81325_index226 <= p5_tuple_index_82004_comb;
    p5_tuple_81325_index227 <= p5_tuple_index_82007_comb;
    p5_tuple_81325_index228 <= p5_tuple_index_82010_comb;
    p5_tuple_81325_index229 <= p5_tuple_index_82013_comb;
    p5_tuple_81325_index230 <= p5_tuple_index_82016_comb;
    p5_tuple_81325_index231 <= p5_tuple_index_82019_comb;
    p5_tuple_81325_index232 <= p5_tuple_index_82022_comb;
    p5_tuple_81325_index233 <= p5_tuple_index_82025_comb;
    p5_tuple_81325_index234 <= p5_tuple_index_82028_comb;
    p5_tuple_81325_index235 <= p5_tuple_index_82031_comb;
    p5_tuple_81325_index236 <= p5_tuple_index_82034_comb;
    p5_tuple_81325_index237 <= p5_tuple_index_82037_comb;
    p5_tuple_81325_index238 <= p5_tuple_index_82040_comb;
    p5_tuple_81325_index239 <= p5_tuple_index_82043_comb;
    p5_tuple_81325_index240 <= p5_tuple_index_82046_comb;
    p5_tuple_81325_index241 <= p5_tuple_index_82049_comb;
    p5_tuple_81325_index242 <= p5_tuple_index_82052_comb;
    p5_tuple_81325_index243 <= p5_tuple_index_82055_comb;
    p5_tuple_81325_index244 <= p5_tuple_index_82058_comb;
    p5_tuple_81325_index245 <= p5_tuple_index_82061_comb;
    p5_tuple_81325_index246 <= p5_tuple_index_82064_comb;
    p5_tuple_81325_index247 <= p5_tuple_index_82067_comb;
    p5_tuple_81325_index248 <= p5_tuple_index_82070_comb;
    p5_tuple_81325_index249 <= p5_tuple_index_82073_comb;
    p5_tuple_81325_index250 <= p5_tuple_index_82076_comb;
    p5_tuple_81325_index251 <= p5_tuple_index_82079_comb;
    p5_tuple_81325_index252 <= p5_tuple_index_82082_comb;
    p5_tuple_81325_index253 <= p5_tuple_index_82085_comb;
    p5_tuple_81325_index254 <= p5_tuple_index_82088_comb;
    p5_tuple_81325_index255 <= p5_tuple_index_82091_comb;
    p5_tuple_81325_index256 <= p5_tuple_index_82094_comb;
    p5_tuple_81325_index257 <= p5_tuple_index_82097_comb;
    p5_tuple_81325_index258 <= p5_tuple_index_82100_comb;
    p5_tuple_81325_index259 <= p5_tuple_index_82103_comb;
    p5_tuple_81325_index260 <= p5_tuple_index_82106_comb;
    p5_tuple_81325_index261 <= p5_tuple_index_82109_comb;
    p5_tuple_81325_index262 <= p5_tuple_index_82112_comb;
    p5_tuple_81325_index263 <= p5_tuple_index_82115_comb;
    p5_tuple_81325_index264 <= p5_tuple_index_82118_comb;
    p5_tuple_81325_index265 <= p5_tuple_index_82121_comb;
    p5_tuple_81325_index266 <= p5_tuple_index_82124_comb;
    p5_tuple_81325_index267 <= p5_tuple_index_82127_comb;
    p5_tuple_81325_index268 <= p5_tuple_index_82130_comb;
    p5_tuple_81325_index269 <= p5_tuple_index_82133_comb;
    p5_tuple_81325_index270 <= p5_tuple_index_82136_comb;
    p5_tuple_81325_index271 <= p5_tuple_index_82139_comb;
    p5_tuple_81325_index272 <= p5_tuple_index_82142_comb;
    p5_tuple_81325_index273 <= p5_tuple_index_82145_comb;
    p5_tuple_81325_index274 <= p5_tuple_index_82148_comb;
    p5_tuple_81325_index275 <= p5_tuple_index_82151_comb;
    p5_tuple_81325_index276 <= p5_tuple_index_82154_comb;
    p5_tuple_81325_index277 <= p5_tuple_index_82157_comb;
    p5_tuple_81325_index278 <= p5_tuple_index_82160_comb;
    p5_tuple_81325_index279 <= p5_tuple_index_82163_comb;
    p5_tuple_81325_index280 <= p5_tuple_index_82166_comb;
    p5_tuple_81325_index281 <= p5_tuple_index_82169_comb;
    p5_tuple_81325_index282 <= p5_tuple_index_82172_comb;
    p5_tuple_81325_index283 <= p5_tuple_index_82175_comb;
    p5_tuple_81325_index284 <= p5_tuple_index_82178_comb;
    p5_tuple_81325_index285 <= p5_tuple_index_82181_comb;
    p5_tuple_81325_index286 <= p5_tuple_index_82184_comb;
    p5_tuple_81325_index287 <= p5_tuple_index_82187_comb;
    p5_tuple_81325_index288 <= p5_tuple_index_82190_comb;
    p5_tuple_81325_index289 <= p5_tuple_index_82193_comb;
    p5_tuple_81325_index290 <= p5_tuple_index_82196_comb;
    p5_tuple_81325_index291 <= p5_tuple_index_82199_comb;
    p5_tuple_81325_index292 <= p5_tuple_index_82202_comb;
    p5_tuple_81325_index293 <= p5_tuple_index_82205_comb;
    p5_tuple_81325_index294 <= p5_tuple_index_82208_comb;
    p5_tuple_81325_index295 <= p5_tuple_index_82211_comb;
    p5_tuple_81325_index296 <= p5_tuple_index_82214_comb;
    p5_tuple_81325_index297 <= p5_tuple_index_82217_comb;
    p5_tuple_81325_index298 <= p5_tuple_index_82220_comb;
    p5_tuple_81325_index299 <= p5_tuple_index_82223_comb;
    p5_tuple_81325_index300 <= p5_tuple_index_82226_comb;
  end

  // ===== Pipe stage 6:
  assign out = {p5_tuple_81325_index1, p5_tuple_81325_index2, p5_tuple_81325_index3, p5_tuple_81325_index4, p5_tuple_81325_index5, p5_tuple_81325_index6, p5_tuple_81325_index7, p5_tuple_81325_index8, p5_tuple_81325_index9, p5_tuple_81325_index10, p5_tuple_81325_index11, p5_tuple_81325_index12, p5_tuple_81325_index13, p5_tuple_81325_index14, p5_tuple_81325_index15, p5_tuple_81325_index16, p5_tuple_81325_index17, p5_tuple_81325_index18, p5_tuple_81325_index19, p5_tuple_81325_index20, p5_tuple_81325_index21, p5_tuple_81325_index22, p5_tuple_81325_index23, p5_tuple_81325_index24, p5_tuple_81325_index25, p5_tuple_81325_index26, p5_tuple_81325_index27, p5_tuple_81325_index28, p5_tuple_81325_index29, p5_tuple_81325_index30, p5_tuple_81325_index31, p5_tuple_81325_index32, p5_tuple_81325_index33, p5_tuple_81325_index34, p5_tuple_81325_index35, p5_tuple_81325_index36, p5_tuple_81325_index37, p5_tuple_81325_index38, p5_tuple_81325_index39, p5_tuple_81325_index40, p5_tuple_81325_index41, p5_tuple_81325_index42, p5_tuple_81325_index43, p5_tuple_81325_index44, p5_tuple_81325_index45, p5_tuple_81325_index46, p5_tuple_81325_index47, p5_tuple_81325_index48, p5_tuple_81325_index49, p5_tuple_81325_index50, p5_tuple_81325_index51, p5_tuple_81325_index52, p5_tuple_81325_index53, p5_tuple_81325_index54, p5_tuple_81325_index55, p5_tuple_81325_index56, p5_tuple_81325_index57, p5_tuple_81325_index58, p5_tuple_81325_index59, p5_tuple_81325_index60, p5_tuple_81325_index61, p5_tuple_81325_index62, p5_tuple_81325_index63, p5_tuple_81325_index64, p5_tuple_81325_index65, p5_tuple_81325_index66, p5_tuple_81325_index67, p5_tuple_81325_index68, p5_tuple_81325_index69, p5_tuple_81325_index70, p5_tuple_81325_index71, p5_tuple_81325_index72, p5_tuple_81325_index73, p5_tuple_81325_index74, p5_tuple_81325_index75, p5_tuple_81325_index76, p5_tuple_81325_index77, p5_tuple_81325_index78, p5_tuple_81325_index79, p5_tuple_81325_index80, p5_tuple_81325_index81, p5_tuple_81325_index82, p5_tuple_81325_index83, p5_tuple_81325_index84, p5_tuple_81325_index85, p5_tuple_81325_index86, p5_tuple_81325_index87, p5_tuple_81325_index88, p5_tuple_81325_index89, p5_tuple_81325_index90, p5_tuple_81325_index91, p5_tuple_81325_index92, p5_tuple_81325_index93, p5_tuple_81325_index94, p5_tuple_81325_index95, p5_tuple_81325_index96, p5_tuple_81325_index97, p5_tuple_81325_index98, p5_tuple_81325_index99, p5_tuple_81325_index100, p5_tuple_81325_index101, p5_tuple_81325_index102, p5_tuple_81325_index103, p5_tuple_81325_index104, p5_tuple_81325_index105, p5_tuple_81325_index106, p5_tuple_81325_index107, p5_tuple_81325_index108, p5_tuple_81325_index109, p5_tuple_81325_index110, p5_tuple_81325_index111, p5_tuple_81325_index112, p5_tuple_81325_index113, p5_tuple_81325_index114, p5_tuple_81325_index115, p5_tuple_81325_index116, p5_tuple_81325_index117, p5_tuple_81325_index118, p5_tuple_81325_index119, p5_tuple_81325_index120, p5_tuple_81325_index121, p5_tuple_81325_index122, p5_tuple_81325_index123, p5_tuple_81325_index124, p5_tuple_81325_index125, p5_tuple_81325_index126, p5_tuple_81325_index127, p5_tuple_81325_index128, p5_tuple_81325_index129, p5_tuple_81325_index130, p5_tuple_81325_index131, p5_tuple_81325_index132, p5_tuple_81325_index133, p5_tuple_81325_index134, p5_tuple_81325_index135, p5_tuple_81325_index136, p5_tuple_81325_index137, p5_tuple_81325_index138, p5_tuple_81325_index139, p5_tuple_81325_index140, p5_tuple_81325_index141, p5_tuple_81325_index142, p5_tuple_81325_index143, p5_tuple_81325_index144, p5_tuple_81325_index145, p5_tuple_81325_index146, p5_tuple_81325_index147, p5_tuple_81325_index148, p5_tuple_81325_index149, p5_tuple_81325_index150, p5_tuple_81325_index151, p5_tuple_81325_index152, p5_tuple_81325_index153, p5_tuple_81325_index154, p5_tuple_81325_index155, p5_tuple_81325_index156, p5_tuple_81325_index157, p5_tuple_81325_index158, p5_tuple_81325_index159, p5_tuple_81325_index160, p5_tuple_81325_index161, p5_tuple_81325_index162, p5_tuple_81325_index163, p5_tuple_81325_index164, p5_tuple_81325_index165, p5_tuple_81325_index166, p5_tuple_81325_index167, p5_tuple_81325_index168, p5_tuple_81325_index169, p5_tuple_81325_index170, p5_tuple_81325_index171, p5_tuple_81325_index172, p5_tuple_81325_index173, p5_tuple_81325_index174, p5_tuple_81325_index175, p5_tuple_81325_index176, p5_tuple_81325_index177, p5_tuple_81325_index178, p5_tuple_81325_index179, p5_tuple_81325_index180, p5_tuple_81325_index181, p5_tuple_81325_index182, p5_tuple_81325_index183, p5_tuple_81325_index184, p5_tuple_81325_index185, p5_tuple_81325_index186, p5_tuple_81325_index187, p5_tuple_81325_index188, p5_tuple_81325_index189, p5_tuple_81325_index190, p5_tuple_81325_index191, p5_tuple_81325_index192, p5_tuple_81325_index193, p5_tuple_81325_index194, p5_tuple_81325_index195, p5_tuple_81325_index196, p5_tuple_81325_index197, p5_tuple_81325_index198, p5_tuple_81325_index199, p5_tuple_81325_index200, p5_tuple_81325_index201, p5_tuple_81325_index202, p5_tuple_81325_index203, p5_tuple_81325_index204, p5_tuple_81325_index205, p5_tuple_81325_index206, p5_tuple_81325_index207, p5_tuple_81325_index208, p5_tuple_81325_index209, p5_tuple_81325_index210, p5_tuple_81325_index211, p5_tuple_81325_index212, p5_tuple_81325_index213, p5_tuple_81325_index214, p5_tuple_81325_index215, p5_tuple_81325_index216, p5_tuple_81325_index217, p5_tuple_81325_index218, p5_tuple_81325_index219, p5_tuple_81325_index220, p5_tuple_81325_index221, p5_tuple_81325_index222, p5_tuple_81325_index223, p5_tuple_81325_index224, p5_tuple_81325_index225, p5_tuple_81325_index226, p5_tuple_81325_index227, p5_tuple_81325_index228, p5_tuple_81325_index229, p5_tuple_81325_index230, p5_tuple_81325_index231, p5_tuple_81325_index232, p5_tuple_81325_index233, p5_tuple_81325_index234, p5_tuple_81325_index235, p5_tuple_81325_index236, p5_tuple_81325_index237, p5_tuple_81325_index238, p5_tuple_81325_index239, p5_tuple_81325_index240, p5_tuple_81325_index241, p5_tuple_81325_index242, p5_tuple_81325_index243, p5_tuple_81325_index244, p5_tuple_81325_index245, p5_tuple_81325_index246, p5_tuple_81325_index247, p5_tuple_81325_index248, p5_tuple_81325_index249, p5_tuple_81325_index250, p5_tuple_81325_index251, p5_tuple_81325_index252, p5_tuple_81325_index253, p5_tuple_81325_index254, p5_tuple_81325_index255, p5_tuple_81325_index256, p5_tuple_81325_index257, p5_tuple_81325_index258, p5_tuple_81325_index259, p5_tuple_81325_index260, p5_tuple_81325_index261, p5_tuple_81325_index262, p5_tuple_81325_index263, p5_tuple_81325_index264, p5_tuple_81325_index265, p5_tuple_81325_index266, p5_tuple_81325_index267, p5_tuple_81325_index268, p5_tuple_81325_index269, p5_tuple_81325_index270, p5_tuple_81325_index271, p5_tuple_81325_index272, p5_tuple_81325_index273, p5_tuple_81325_index274, p5_tuple_81325_index275, p5_tuple_81325_index276, p5_tuple_81325_index277, p5_tuple_81325_index278, p5_tuple_81325_index279, p5_tuple_81325_index280, p5_tuple_81325_index281, p5_tuple_81325_index282, p5_tuple_81325_index283, p5_tuple_81325_index284, p5_tuple_81325_index285, p5_tuple_81325_index286, p5_tuple_81325_index287, p5_tuple_81325_index288, p5_tuple_81325_index289, p5_tuple_81325_index290, p5_tuple_81325_index291, p5_tuple_81325_index292, p5_tuple_81325_index293, p5_tuple_81325_index294, p5_tuple_81325_index295, p5_tuple_81325_index296, p5_tuple_81325_index297, p5_tuple_81325_index298, p5_tuple_81325_index299, p5_tuple_81325_index300};
endmodule
