module matrix_mul_10_comb(
  input wire [31:0] TestBlock__A_op0,
  input wire [31:0] TestBlock__A_op1,
  input wire [31:0] TestBlock__A_op2,
  input wire [31:0] TestBlock__A_op3,
  input wire [31:0] TestBlock__A_op4,
  input wire [31:0] TestBlock__A_op5,
  input wire [31:0] TestBlock__A_op6,
  input wire [31:0] TestBlock__A_op7,
  input wire [31:0] TestBlock__A_op8,
  input wire [31:0] TestBlock__A_op9,
  input wire [31:0] TestBlock__A_op10,
  input wire [31:0] TestBlock__A_op11,
  input wire [31:0] TestBlock__A_op12,
  input wire [31:0] TestBlock__A_op13,
  input wire [31:0] TestBlock__A_op14,
  input wire [31:0] TestBlock__A_op15,
  input wire [31:0] TestBlock__A_op16,
  input wire [31:0] TestBlock__A_op17,
  input wire [31:0] TestBlock__A_op18,
  input wire [31:0] TestBlock__A_op19,
  input wire [31:0] TestBlock__A_op20,
  input wire [31:0] TestBlock__A_op21,
  input wire [31:0] TestBlock__A_op22,
  input wire [31:0] TestBlock__A_op23,
  input wire [31:0] TestBlock__A_op24,
  input wire [31:0] TestBlock__A_op25,
  input wire [31:0] TestBlock__A_op26,
  input wire [31:0] TestBlock__A_op27,
  input wire [31:0] TestBlock__A_op28,
  input wire [31:0] TestBlock__A_op29,
  input wire [31:0] TestBlock__A_op30,
  input wire [31:0] TestBlock__A_op31,
  input wire [31:0] TestBlock__A_op32,
  input wire [31:0] TestBlock__A_op33,
  input wire [31:0] TestBlock__A_op34,
  input wire [31:0] TestBlock__A_op35,
  input wire [31:0] TestBlock__A_op36,
  input wire [31:0] TestBlock__A_op37,
  input wire [31:0] TestBlock__A_op38,
  input wire [31:0] TestBlock__A_op39,
  input wire [31:0] TestBlock__A_op40,
  input wire [31:0] TestBlock__A_op41,
  input wire [31:0] TestBlock__A_op42,
  input wire [31:0] TestBlock__A_op43,
  input wire [31:0] TestBlock__A_op44,
  input wire [31:0] TestBlock__A_op45,
  input wire [31:0] TestBlock__A_op46,
  input wire [31:0] TestBlock__A_op47,
  input wire [31:0] TestBlock__A_op48,
  input wire [31:0] TestBlock__A_op49,
  input wire [31:0] TestBlock__A_op50,
  input wire [31:0] TestBlock__A_op51,
  input wire [31:0] TestBlock__A_op52,
  input wire [31:0] TestBlock__A_op53,
  input wire [31:0] TestBlock__A_op54,
  input wire [31:0] TestBlock__A_op55,
  input wire [31:0] TestBlock__A_op56,
  input wire [31:0] TestBlock__A_op57,
  input wire [31:0] TestBlock__A_op58,
  input wire [31:0] TestBlock__A_op59,
  input wire [31:0] TestBlock__A_op60,
  input wire [31:0] TestBlock__A_op61,
  input wire [31:0] TestBlock__A_op62,
  input wire [31:0] TestBlock__A_op63,
  input wire [31:0] TestBlock__A_op64,
  input wire [31:0] TestBlock__A_op65,
  input wire [31:0] TestBlock__A_op66,
  input wire [31:0] TestBlock__A_op67,
  input wire [31:0] TestBlock__A_op68,
  input wire [31:0] TestBlock__A_op69,
  input wire [31:0] TestBlock__A_op70,
  input wire [31:0] TestBlock__A_op71,
  input wire [31:0] TestBlock__A_op72,
  input wire [31:0] TestBlock__A_op73,
  input wire [31:0] TestBlock__A_op74,
  input wire [31:0] TestBlock__A_op75,
  input wire [31:0] TestBlock__A_op76,
  input wire [31:0] TestBlock__A_op77,
  input wire [31:0] TestBlock__A_op78,
  input wire [31:0] TestBlock__A_op79,
  input wire [31:0] TestBlock__A_op80,
  input wire [31:0] TestBlock__A_op81,
  input wire [31:0] TestBlock__A_op82,
  input wire [31:0] TestBlock__A_op83,
  input wire [31:0] TestBlock__A_op84,
  input wire [31:0] TestBlock__A_op85,
  input wire [31:0] TestBlock__A_op86,
  input wire [31:0] TestBlock__A_op87,
  input wire [31:0] TestBlock__A_op88,
  input wire [31:0] TestBlock__A_op89,
  input wire [31:0] TestBlock__A_op90,
  input wire [31:0] TestBlock__A_op91,
  input wire [31:0] TestBlock__A_op92,
  input wire [31:0] TestBlock__A_op93,
  input wire [31:0] TestBlock__A_op94,
  input wire [31:0] TestBlock__A_op95,
  input wire [31:0] TestBlock__A_op96,
  input wire [31:0] TestBlock__A_op97,
  input wire [31:0] TestBlock__A_op98,
  input wire [31:0] TestBlock__A_op99,
  input wire [31:0] TestBlock__B_op0,
  input wire [31:0] TestBlock__B_op1,
  input wire [31:0] TestBlock__B_op2,
  input wire [31:0] TestBlock__B_op3,
  input wire [31:0] TestBlock__B_op4,
  input wire [31:0] TestBlock__B_op5,
  input wire [31:0] TestBlock__B_op6,
  input wire [31:0] TestBlock__B_op7,
  input wire [31:0] TestBlock__B_op8,
  input wire [31:0] TestBlock__B_op9,
  input wire [31:0] TestBlock__B_op10,
  input wire [31:0] TestBlock__B_op11,
  input wire [31:0] TestBlock__B_op12,
  input wire [31:0] TestBlock__B_op13,
  input wire [31:0] TestBlock__B_op14,
  input wire [31:0] TestBlock__B_op15,
  input wire [31:0] TestBlock__B_op16,
  input wire [31:0] TestBlock__B_op17,
  input wire [31:0] TestBlock__B_op18,
  input wire [31:0] TestBlock__B_op19,
  input wire [31:0] TestBlock__B_op20,
  input wire [31:0] TestBlock__B_op21,
  input wire [31:0] TestBlock__B_op22,
  input wire [31:0] TestBlock__B_op23,
  input wire [31:0] TestBlock__B_op24,
  input wire [31:0] TestBlock__B_op25,
  input wire [31:0] TestBlock__B_op26,
  input wire [31:0] TestBlock__B_op27,
  input wire [31:0] TestBlock__B_op28,
  input wire [31:0] TestBlock__B_op29,
  input wire [31:0] TestBlock__B_op30,
  input wire [31:0] TestBlock__B_op31,
  input wire [31:0] TestBlock__B_op32,
  input wire [31:0] TestBlock__B_op33,
  input wire [31:0] TestBlock__B_op34,
  input wire [31:0] TestBlock__B_op35,
  input wire [31:0] TestBlock__B_op36,
  input wire [31:0] TestBlock__B_op37,
  input wire [31:0] TestBlock__B_op38,
  input wire [31:0] TestBlock__B_op39,
  input wire [31:0] TestBlock__B_op40,
  input wire [31:0] TestBlock__B_op41,
  input wire [31:0] TestBlock__B_op42,
  input wire [31:0] TestBlock__B_op43,
  input wire [31:0] TestBlock__B_op44,
  input wire [31:0] TestBlock__B_op45,
  input wire [31:0] TestBlock__B_op46,
  input wire [31:0] TestBlock__B_op47,
  input wire [31:0] TestBlock__B_op48,
  input wire [31:0] TestBlock__B_op49,
  input wire [31:0] TestBlock__B_op50,
  input wire [31:0] TestBlock__B_op51,
  input wire [31:0] TestBlock__B_op52,
  input wire [31:0] TestBlock__B_op53,
  input wire [31:0] TestBlock__B_op54,
  input wire [31:0] TestBlock__B_op55,
  input wire [31:0] TestBlock__B_op56,
  input wire [31:0] TestBlock__B_op57,
  input wire [31:0] TestBlock__B_op58,
  input wire [31:0] TestBlock__B_op59,
  input wire [31:0] TestBlock__B_op60,
  input wire [31:0] TestBlock__B_op61,
  input wire [31:0] TestBlock__B_op62,
  input wire [31:0] TestBlock__B_op63,
  input wire [31:0] TestBlock__B_op64,
  input wire [31:0] TestBlock__B_op65,
  input wire [31:0] TestBlock__B_op66,
  input wire [31:0] TestBlock__B_op67,
  input wire [31:0] TestBlock__B_op68,
  input wire [31:0] TestBlock__B_op69,
  input wire [31:0] TestBlock__B_op70,
  input wire [31:0] TestBlock__B_op71,
  input wire [31:0] TestBlock__B_op72,
  input wire [31:0] TestBlock__B_op73,
  input wire [31:0] TestBlock__B_op74,
  input wire [31:0] TestBlock__B_op75,
  input wire [31:0] TestBlock__B_op76,
  input wire [31:0] TestBlock__B_op77,
  input wire [31:0] TestBlock__B_op78,
  input wire [31:0] TestBlock__B_op79,
  input wire [31:0] TestBlock__B_op80,
  input wire [31:0] TestBlock__B_op81,
  input wire [31:0] TestBlock__B_op82,
  input wire [31:0] TestBlock__B_op83,
  input wire [31:0] TestBlock__B_op84,
  input wire [31:0] TestBlock__B_op85,
  input wire [31:0] TestBlock__B_op86,
  input wire [31:0] TestBlock__B_op87,
  input wire [31:0] TestBlock__B_op88,
  input wire [31:0] TestBlock__B_op89,
  input wire [31:0] TestBlock__B_op90,
  input wire [31:0] TestBlock__B_op91,
  input wire [31:0] TestBlock__B_op92,
  input wire [31:0] TestBlock__B_op93,
  input wire [31:0] TestBlock__B_op94,
  input wire [31:0] TestBlock__B_op95,
  input wire [31:0] TestBlock__B_op96,
  input wire [31:0] TestBlock__B_op97,
  input wire [31:0] TestBlock__B_op98,
  input wire [31:0] TestBlock__B_op99,
  output wire [3499:0] out
);
  // lint_off SIGNED_TYPE
  // lint_off MULTIPLY
  function automatic [31:0] smul32b_32b_x_32b (input reg [31:0] lhs, input reg [31:0] rhs);
    reg signed [31:0] signed_lhs;
    reg signed [31:0] signed_rhs;
    reg signed [31:0] signed_result;
    begin
      signed_lhs = $signed(lhs);
      signed_rhs = $signed(rhs);
      signed_result = signed_lhs * signed_rhs;
      smul32b_32b_x_32b = $unsigned(signed_result);
    end
  endfunction
  // lint_on MULTIPLY
  // lint_on SIGNED_TYPE
  wire [31:0] smul_75273;
  wire [31:0] smul_75274;
  wire [31:0] smul_75275;
  wire [31:0] smul_75276;
  wire [31:0] smul_75277;
  wire [31:0] smul_75278;
  wire [31:0] smul_75279;
  wire [31:0] smul_75280;
  wire [31:0] smul_75281;
  wire [31:0] smul_75282;
  wire [31:0] smul_75283;
  wire [31:0] smul_75284;
  wire [31:0] smul_75285;
  wire [31:0] smul_75286;
  wire [31:0] smul_75287;
  wire [31:0] smul_75288;
  wire [31:0] smul_75289;
  wire [31:0] smul_75290;
  wire [31:0] smul_75291;
  wire [31:0] smul_75292;
  wire [31:0] smul_75293;
  wire [31:0] smul_75294;
  wire [31:0] smul_75295;
  wire [31:0] smul_75296;
  wire [31:0] smul_75297;
  wire [31:0] smul_75298;
  wire [31:0] smul_75299;
  wire [31:0] smul_75300;
  wire [31:0] smul_75301;
  wire [31:0] smul_75302;
  wire [31:0] smul_75303;
  wire [31:0] smul_75304;
  wire [31:0] smul_75305;
  wire [31:0] smul_75306;
  wire [31:0] smul_75307;
  wire [31:0] smul_75308;
  wire [31:0] smul_75309;
  wire [31:0] smul_75310;
  wire [31:0] smul_75311;
  wire [31:0] smul_75312;
  wire [31:0] smul_75313;
  wire [31:0] smul_75314;
  wire [31:0] smul_75315;
  wire [31:0] smul_75316;
  wire [31:0] smul_75317;
  wire [31:0] smul_75318;
  wire [31:0] smul_75319;
  wire [31:0] smul_75320;
  wire [31:0] smul_75321;
  wire [31:0] smul_75322;
  wire [31:0] smul_75323;
  wire [31:0] smul_75324;
  wire [31:0] smul_75325;
  wire [31:0] smul_75326;
  wire [31:0] smul_75327;
  wire [31:0] smul_75328;
  wire [31:0] smul_75329;
  wire [31:0] smul_75330;
  wire [31:0] smul_75331;
  wire [31:0] smul_75332;
  wire [31:0] smul_75333;
  wire [31:0] smul_75334;
  wire [31:0] smul_75335;
  wire [31:0] smul_75336;
  wire [31:0] smul_75337;
  wire [31:0] smul_75338;
  wire [31:0] smul_75339;
  wire [31:0] smul_75340;
  wire [31:0] smul_75341;
  wire [31:0] smul_75342;
  wire [31:0] smul_75343;
  wire [31:0] smul_75344;
  wire [31:0] smul_75345;
  wire [31:0] smul_75346;
  wire [31:0] smul_75347;
  wire [31:0] smul_75348;
  wire [31:0] smul_75349;
  wire [31:0] smul_75350;
  wire [31:0] smul_75351;
  wire [31:0] smul_75352;
  wire [31:0] smul_75353;
  wire [31:0] smul_75354;
  wire [31:0] smul_75355;
  wire [31:0] smul_75356;
  wire [31:0] smul_75357;
  wire [31:0] smul_75358;
  wire [31:0] smul_75359;
  wire [31:0] smul_75360;
  wire [31:0] smul_75361;
  wire [31:0] smul_75362;
  wire [31:0] smul_75363;
  wire [31:0] smul_75364;
  wire [31:0] smul_75365;
  wire [31:0] smul_75366;
  wire [31:0] smul_75367;
  wire [31:0] smul_75368;
  wire [31:0] smul_75369;
  wire [31:0] smul_75370;
  wire [31:0] smul_75371;
  wire [31:0] smul_75372;
  wire [31:0] smul_75373;
  wire [31:0] smul_75374;
  wire [31:0] smul_75375;
  wire [31:0] smul_75376;
  wire [31:0] smul_75377;
  wire [31:0] smul_75378;
  wire [31:0] smul_75379;
  wire [31:0] smul_75380;
  wire [31:0] smul_75381;
  wire [31:0] smul_75382;
  wire [31:0] smul_75383;
  wire [31:0] smul_75384;
  wire [31:0] smul_75385;
  wire [31:0] smul_75386;
  wire [31:0] smul_75387;
  wire [31:0] smul_75388;
  wire [31:0] smul_75389;
  wire [31:0] smul_75390;
  wire [31:0] smul_75391;
  wire [31:0] smul_75392;
  wire [31:0] smul_75393;
  wire [31:0] smul_75394;
  wire [31:0] smul_75395;
  wire [31:0] smul_75396;
  wire [31:0] smul_75397;
  wire [31:0] smul_75398;
  wire [31:0] smul_75399;
  wire [31:0] smul_75400;
  wire [31:0] smul_75401;
  wire [31:0] smul_75402;
  wire [31:0] smul_75403;
  wire [31:0] smul_75404;
  wire [31:0] smul_75405;
  wire [31:0] smul_75406;
  wire [31:0] smul_75407;
  wire [31:0] smul_75408;
  wire [31:0] smul_75409;
  wire [31:0] smul_75410;
  wire [31:0] smul_75411;
  wire [31:0] smul_75412;
  wire [31:0] smul_75413;
  wire [31:0] smul_75414;
  wire [31:0] smul_75415;
  wire [31:0] smul_75416;
  wire [31:0] smul_75417;
  wire [31:0] smul_75418;
  wire [31:0] smul_75419;
  wire [31:0] smul_75420;
  wire [31:0] smul_75421;
  wire [31:0] smul_75422;
  wire [31:0] smul_75423;
  wire [31:0] smul_75424;
  wire [31:0] smul_75425;
  wire [31:0] smul_75426;
  wire [31:0] smul_75427;
  wire [31:0] smul_75428;
  wire [31:0] smul_75429;
  wire [31:0] smul_75430;
  wire [31:0] smul_75431;
  wire [31:0] smul_75432;
  wire [31:0] smul_75433;
  wire [31:0] smul_75434;
  wire [31:0] smul_75435;
  wire [31:0] smul_75436;
  wire [31:0] smul_75437;
  wire [31:0] smul_75438;
  wire [31:0] smul_75439;
  wire [31:0] smul_75440;
  wire [31:0] smul_75441;
  wire [31:0] smul_75442;
  wire [31:0] smul_75443;
  wire [31:0] smul_75444;
  wire [31:0] smul_75445;
  wire [31:0] smul_75446;
  wire [31:0] smul_75447;
  wire [31:0] smul_75448;
  wire [31:0] smul_75449;
  wire [31:0] smul_75450;
  wire [31:0] smul_75451;
  wire [31:0] smul_75452;
  wire [31:0] smul_75453;
  wire [31:0] smul_75454;
  wire [31:0] smul_75455;
  wire [31:0] smul_75456;
  wire [31:0] smul_75457;
  wire [31:0] smul_75458;
  wire [31:0] smul_75459;
  wire [31:0] smul_75460;
  wire [31:0] smul_75461;
  wire [31:0] smul_75462;
  wire [31:0] smul_75463;
  wire [31:0] smul_75464;
  wire [31:0] smul_75465;
  wire [31:0] smul_75466;
  wire [31:0] smul_75467;
  wire [31:0] smul_75468;
  wire [31:0] smul_75469;
  wire [31:0] smul_75470;
  wire [31:0] smul_75471;
  wire [31:0] smul_75472;
  wire [31:0] smul_75473;
  wire [31:0] smul_75474;
  wire [31:0] smul_75475;
  wire [31:0] smul_75476;
  wire [31:0] smul_75477;
  wire [31:0] smul_75478;
  wire [31:0] smul_75479;
  wire [31:0] smul_75480;
  wire [31:0] smul_75481;
  wire [31:0] smul_75482;
  wire [31:0] smul_75483;
  wire [31:0] smul_75484;
  wire [31:0] smul_75485;
  wire [31:0] smul_75486;
  wire [31:0] smul_75487;
  wire [31:0] smul_75488;
  wire [31:0] smul_75489;
  wire [31:0] smul_75490;
  wire [31:0] smul_75491;
  wire [31:0] smul_75492;
  wire [31:0] smul_75493;
  wire [31:0] smul_75494;
  wire [31:0] smul_75495;
  wire [31:0] smul_75496;
  wire [31:0] smul_75497;
  wire [31:0] smul_75498;
  wire [31:0] smul_75499;
  wire [31:0] smul_75500;
  wire [31:0] smul_75501;
  wire [31:0] smul_75502;
  wire [31:0] smul_75503;
  wire [31:0] smul_75504;
  wire [31:0] smul_75505;
  wire [31:0] smul_75506;
  wire [31:0] smul_75507;
  wire [31:0] smul_75508;
  wire [31:0] smul_75509;
  wire [31:0] smul_75510;
  wire [31:0] smul_75511;
  wire [31:0] smul_75512;
  wire [31:0] smul_75513;
  wire [31:0] smul_75514;
  wire [31:0] smul_75515;
  wire [31:0] smul_75516;
  wire [31:0] smul_75517;
  wire [31:0] smul_75518;
  wire [31:0] smul_75519;
  wire [31:0] smul_75520;
  wire [31:0] smul_75521;
  wire [31:0] smul_75522;
  wire [31:0] smul_75523;
  wire [31:0] smul_75524;
  wire [31:0] smul_75525;
  wire [31:0] smul_75526;
  wire [31:0] smul_75527;
  wire [31:0] smul_75528;
  wire [31:0] smul_75529;
  wire [31:0] smul_75530;
  wire [31:0] smul_75531;
  wire [31:0] smul_75532;
  wire [31:0] smul_75533;
  wire [31:0] smul_75534;
  wire [31:0] smul_75535;
  wire [31:0] smul_75536;
  wire [31:0] smul_75537;
  wire [31:0] smul_75538;
  wire [31:0] smul_75539;
  wire [31:0] smul_75540;
  wire [31:0] smul_75541;
  wire [31:0] smul_75542;
  wire [31:0] smul_75543;
  wire [31:0] smul_75544;
  wire [31:0] smul_75545;
  wire [31:0] smul_75546;
  wire [31:0] smul_75547;
  wire [31:0] smul_75548;
  wire [31:0] smul_75549;
  wire [31:0] smul_75550;
  wire [31:0] smul_75551;
  wire [31:0] smul_75552;
  wire [31:0] smul_75553;
  wire [31:0] smul_75554;
  wire [31:0] smul_75555;
  wire [31:0] smul_75556;
  wire [31:0] smul_75557;
  wire [31:0] smul_75558;
  wire [31:0] smul_75559;
  wire [31:0] smul_75560;
  wire [31:0] smul_75561;
  wire [31:0] smul_75562;
  wire [31:0] smul_75563;
  wire [31:0] smul_75564;
  wire [31:0] smul_75565;
  wire [31:0] smul_75566;
  wire [31:0] smul_75567;
  wire [31:0] smul_75568;
  wire [31:0] smul_75569;
  wire [31:0] smul_75570;
  wire [31:0] smul_75571;
  wire [31:0] smul_75572;
  wire [31:0] smul_75573;
  wire [31:0] smul_75574;
  wire [31:0] smul_75575;
  wire [31:0] smul_75576;
  wire [31:0] smul_75577;
  wire [31:0] smul_75578;
  wire [31:0] smul_75579;
  wire [31:0] smul_75580;
  wire [31:0] smul_75581;
  wire [31:0] smul_75582;
  wire [31:0] smul_75583;
  wire [31:0] smul_75584;
  wire [31:0] smul_75585;
  wire [31:0] smul_75586;
  wire [31:0] smul_75587;
  wire [31:0] smul_75588;
  wire [31:0] smul_75589;
  wire [31:0] smul_75590;
  wire [31:0] smul_75591;
  wire [31:0] smul_75592;
  wire [31:0] smul_75593;
  wire [31:0] smul_75594;
  wire [31:0] smul_75595;
  wire [31:0] smul_75596;
  wire [31:0] smul_75597;
  wire [31:0] smul_75598;
  wire [31:0] smul_75599;
  wire [31:0] smul_75600;
  wire [31:0] smul_75601;
  wire [31:0] smul_75602;
  wire [31:0] smul_75603;
  wire [31:0] smul_75604;
  wire [31:0] smul_75605;
  wire [31:0] smul_75606;
  wire [31:0] smul_75607;
  wire [31:0] smul_75608;
  wire [31:0] smul_75609;
  wire [31:0] smul_75610;
  wire [31:0] smul_75611;
  wire [31:0] smul_75612;
  wire [31:0] smul_75613;
  wire [31:0] smul_75614;
  wire [31:0] smul_75615;
  wire [31:0] smul_75616;
  wire [31:0] smul_75617;
  wire [31:0] smul_75618;
  wire [31:0] smul_75619;
  wire [31:0] smul_75620;
  wire [31:0] smul_75621;
  wire [31:0] smul_75622;
  wire [31:0] smul_75623;
  wire [31:0] smul_75624;
  wire [31:0] smul_75625;
  wire [31:0] smul_75626;
  wire [31:0] smul_75627;
  wire [31:0] smul_75628;
  wire [31:0] smul_75629;
  wire [31:0] smul_75630;
  wire [31:0] smul_75631;
  wire [31:0] smul_75632;
  wire [31:0] smul_75633;
  wire [31:0] smul_75634;
  wire [31:0] smul_75635;
  wire [31:0] smul_75636;
  wire [31:0] smul_75637;
  wire [31:0] smul_75638;
  wire [31:0] smul_75639;
  wire [31:0] smul_75640;
  wire [31:0] smul_75641;
  wire [31:0] smul_75642;
  wire [31:0] smul_75643;
  wire [31:0] smul_75644;
  wire [31:0] smul_75645;
  wire [31:0] smul_75646;
  wire [31:0] smul_75647;
  wire [31:0] smul_75648;
  wire [31:0] smul_75649;
  wire [31:0] smul_75650;
  wire [31:0] smul_75651;
  wire [31:0] smul_75652;
  wire [31:0] smul_75653;
  wire [31:0] smul_75654;
  wire [31:0] smul_75655;
  wire [31:0] smul_75656;
  wire [31:0] smul_75657;
  wire [31:0] smul_75658;
  wire [31:0] smul_75659;
  wire [31:0] smul_75660;
  wire [31:0] smul_75661;
  wire [31:0] smul_75662;
  wire [31:0] smul_75663;
  wire [31:0] smul_75664;
  wire [31:0] smul_75665;
  wire [31:0] smul_75666;
  wire [31:0] smul_75667;
  wire [31:0] smul_75668;
  wire [31:0] smul_75669;
  wire [31:0] smul_75670;
  wire [31:0] smul_75671;
  wire [31:0] smul_75672;
  wire [31:0] add_75673;
  wire [31:0] add_75674;
  wire [31:0] smul_75675;
  wire [31:0] smul_75676;
  wire [31:0] smul_75677;
  wire [31:0] smul_75678;
  wire [31:0] smul_75679;
  wire [31:0] smul_75680;
  wire [31:0] add_75681;
  wire [31:0] add_75682;
  wire [31:0] smul_75683;
  wire [31:0] smul_75684;
  wire [31:0] smul_75685;
  wire [31:0] smul_75686;
  wire [31:0] smul_75687;
  wire [31:0] smul_75688;
  wire [31:0] add_75689;
  wire [31:0] add_75690;
  wire [31:0] smul_75691;
  wire [31:0] smul_75692;
  wire [31:0] smul_75693;
  wire [31:0] smul_75694;
  wire [31:0] smul_75695;
  wire [31:0] smul_75696;
  wire [31:0] add_75697;
  wire [31:0] add_75698;
  wire [31:0] smul_75699;
  wire [31:0] smul_75700;
  wire [31:0] smul_75701;
  wire [31:0] smul_75702;
  wire [31:0] smul_75703;
  wire [31:0] smul_75704;
  wire [31:0] add_75705;
  wire [31:0] add_75706;
  wire [31:0] smul_75707;
  wire [31:0] smul_75708;
  wire [31:0] smul_75709;
  wire [31:0] smul_75710;
  wire [31:0] smul_75711;
  wire [31:0] smul_75712;
  wire [31:0] add_75713;
  wire [31:0] add_75714;
  wire [31:0] smul_75715;
  wire [31:0] smul_75716;
  wire [31:0] smul_75717;
  wire [31:0] smul_75718;
  wire [31:0] smul_75719;
  wire [31:0] smul_75720;
  wire [31:0] add_75721;
  wire [31:0] add_75722;
  wire [31:0] smul_75723;
  wire [31:0] smul_75724;
  wire [31:0] smul_75725;
  wire [31:0] smul_75726;
  wire [31:0] smul_75727;
  wire [31:0] smul_75728;
  wire [31:0] add_75729;
  wire [31:0] add_75730;
  wire [31:0] smul_75731;
  wire [31:0] smul_75732;
  wire [31:0] smul_75733;
  wire [31:0] smul_75734;
  wire [31:0] smul_75735;
  wire [31:0] smul_75736;
  wire [31:0] add_75737;
  wire [31:0] add_75738;
  wire [31:0] smul_75739;
  wire [31:0] smul_75740;
  wire [31:0] smul_75741;
  wire [31:0] smul_75742;
  wire [31:0] smul_75743;
  wire [31:0] smul_75744;
  wire [31:0] add_75745;
  wire [31:0] add_75746;
  wire [31:0] smul_75747;
  wire [31:0] smul_75748;
  wire [31:0] smul_75749;
  wire [31:0] smul_75750;
  wire [31:0] smul_75751;
  wire [31:0] smul_75752;
  wire [31:0] add_75753;
  wire [31:0] add_75754;
  wire [31:0] smul_75755;
  wire [31:0] smul_75756;
  wire [31:0] smul_75757;
  wire [31:0] smul_75758;
  wire [31:0] smul_75759;
  wire [31:0] smul_75760;
  wire [31:0] add_75761;
  wire [31:0] add_75762;
  wire [31:0] smul_75763;
  wire [31:0] smul_75764;
  wire [31:0] smul_75765;
  wire [31:0] smul_75766;
  wire [31:0] smul_75767;
  wire [31:0] smul_75768;
  wire [31:0] add_75769;
  wire [31:0] add_75770;
  wire [31:0] smul_75771;
  wire [31:0] smul_75772;
  wire [31:0] smul_75773;
  wire [31:0] smul_75774;
  wire [31:0] smul_75775;
  wire [31:0] smul_75776;
  wire [31:0] add_75777;
  wire [31:0] add_75778;
  wire [31:0] smul_75779;
  wire [31:0] smul_75780;
  wire [31:0] smul_75781;
  wire [31:0] smul_75782;
  wire [31:0] smul_75783;
  wire [31:0] smul_75784;
  wire [31:0] add_75785;
  wire [31:0] add_75786;
  wire [31:0] smul_75787;
  wire [31:0] smul_75788;
  wire [31:0] smul_75789;
  wire [31:0] smul_75790;
  wire [31:0] smul_75791;
  wire [31:0] smul_75792;
  wire [31:0] add_75793;
  wire [31:0] add_75794;
  wire [31:0] smul_75795;
  wire [31:0] smul_75796;
  wire [31:0] smul_75797;
  wire [31:0] smul_75798;
  wire [31:0] smul_75799;
  wire [31:0] smul_75800;
  wire [31:0] add_75801;
  wire [31:0] add_75802;
  wire [31:0] smul_75803;
  wire [31:0] smul_75804;
  wire [31:0] smul_75805;
  wire [31:0] smul_75806;
  wire [31:0] smul_75807;
  wire [31:0] smul_75808;
  wire [31:0] add_75809;
  wire [31:0] add_75810;
  wire [31:0] smul_75811;
  wire [31:0] smul_75812;
  wire [31:0] smul_75813;
  wire [31:0] smul_75814;
  wire [31:0] smul_75815;
  wire [31:0] smul_75816;
  wire [31:0] add_75817;
  wire [31:0] add_75818;
  wire [31:0] smul_75819;
  wire [31:0] smul_75820;
  wire [31:0] smul_75821;
  wire [31:0] smul_75822;
  wire [31:0] smul_75823;
  wire [31:0] smul_75824;
  wire [31:0] add_75825;
  wire [31:0] add_75826;
  wire [31:0] smul_75827;
  wire [31:0] smul_75828;
  wire [31:0] smul_75829;
  wire [31:0] smul_75830;
  wire [31:0] smul_75831;
  wire [31:0] smul_75832;
  wire [31:0] add_75833;
  wire [31:0] add_75834;
  wire [31:0] smul_75835;
  wire [31:0] smul_75836;
  wire [31:0] smul_75837;
  wire [31:0] smul_75838;
  wire [31:0] smul_75839;
  wire [31:0] smul_75840;
  wire [31:0] add_75841;
  wire [31:0] add_75842;
  wire [31:0] smul_75843;
  wire [31:0] smul_75844;
  wire [31:0] smul_75845;
  wire [31:0] smul_75846;
  wire [31:0] smul_75847;
  wire [31:0] smul_75848;
  wire [31:0] add_75849;
  wire [31:0] add_75850;
  wire [31:0] smul_75851;
  wire [31:0] smul_75852;
  wire [31:0] smul_75853;
  wire [31:0] smul_75854;
  wire [31:0] smul_75855;
  wire [31:0] smul_75856;
  wire [31:0] add_75857;
  wire [31:0] add_75858;
  wire [31:0] smul_75859;
  wire [31:0] smul_75860;
  wire [31:0] smul_75861;
  wire [31:0] smul_75862;
  wire [31:0] smul_75863;
  wire [31:0] smul_75864;
  wire [31:0] add_75865;
  wire [31:0] add_75866;
  wire [31:0] smul_75867;
  wire [31:0] smul_75868;
  wire [31:0] smul_75869;
  wire [31:0] smul_75870;
  wire [31:0] smul_75871;
  wire [31:0] smul_75872;
  wire [31:0] add_75873;
  wire [31:0] add_75874;
  wire [31:0] smul_75875;
  wire [31:0] smul_75876;
  wire [31:0] smul_75877;
  wire [31:0] smul_75878;
  wire [31:0] smul_75879;
  wire [31:0] smul_75880;
  wire [31:0] add_75881;
  wire [31:0] add_75882;
  wire [31:0] smul_75883;
  wire [31:0] smul_75884;
  wire [31:0] smul_75885;
  wire [31:0] smul_75886;
  wire [31:0] smul_75887;
  wire [31:0] smul_75888;
  wire [31:0] add_75889;
  wire [31:0] add_75890;
  wire [31:0] smul_75891;
  wire [31:0] smul_75892;
  wire [31:0] smul_75893;
  wire [31:0] smul_75894;
  wire [31:0] smul_75895;
  wire [31:0] smul_75896;
  wire [31:0] add_75897;
  wire [31:0] add_75898;
  wire [31:0] smul_75899;
  wire [31:0] smul_75900;
  wire [31:0] smul_75901;
  wire [31:0] smul_75902;
  wire [31:0] smul_75903;
  wire [31:0] smul_75904;
  wire [31:0] add_75905;
  wire [31:0] add_75906;
  wire [31:0] smul_75907;
  wire [31:0] smul_75908;
  wire [31:0] smul_75909;
  wire [31:0] smul_75910;
  wire [31:0] smul_75911;
  wire [31:0] smul_75912;
  wire [31:0] add_75913;
  wire [31:0] add_75914;
  wire [31:0] smul_75915;
  wire [31:0] smul_75916;
  wire [31:0] smul_75917;
  wire [31:0] smul_75918;
  wire [31:0] smul_75919;
  wire [31:0] smul_75920;
  wire [31:0] add_75921;
  wire [31:0] add_75922;
  wire [31:0] smul_75923;
  wire [31:0] smul_75924;
  wire [31:0] smul_75925;
  wire [31:0] smul_75926;
  wire [31:0] smul_75927;
  wire [31:0] smul_75928;
  wire [31:0] add_75929;
  wire [31:0] add_75930;
  wire [31:0] smul_75931;
  wire [31:0] smul_75932;
  wire [31:0] smul_75933;
  wire [31:0] smul_75934;
  wire [31:0] smul_75935;
  wire [31:0] smul_75936;
  wire [31:0] add_75937;
  wire [31:0] add_75938;
  wire [31:0] smul_75939;
  wire [31:0] smul_75940;
  wire [31:0] smul_75941;
  wire [31:0] smul_75942;
  wire [31:0] smul_75943;
  wire [31:0] smul_75944;
  wire [31:0] add_75945;
  wire [31:0] add_75946;
  wire [31:0] smul_75947;
  wire [31:0] smul_75948;
  wire [31:0] smul_75949;
  wire [31:0] smul_75950;
  wire [31:0] smul_75951;
  wire [31:0] smul_75952;
  wire [31:0] add_75953;
  wire [31:0] add_75954;
  wire [31:0] smul_75955;
  wire [31:0] smul_75956;
  wire [31:0] smul_75957;
  wire [31:0] smul_75958;
  wire [31:0] smul_75959;
  wire [31:0] smul_75960;
  wire [31:0] add_75961;
  wire [31:0] add_75962;
  wire [31:0] smul_75963;
  wire [31:0] smul_75964;
  wire [31:0] smul_75965;
  wire [31:0] smul_75966;
  wire [31:0] smul_75967;
  wire [31:0] smul_75968;
  wire [31:0] add_75969;
  wire [31:0] add_75970;
  wire [31:0] smul_75971;
  wire [31:0] smul_75972;
  wire [31:0] smul_75973;
  wire [31:0] smul_75974;
  wire [31:0] smul_75975;
  wire [31:0] smul_75976;
  wire [31:0] add_75977;
  wire [31:0] add_75978;
  wire [31:0] smul_75979;
  wire [31:0] smul_75980;
  wire [31:0] smul_75981;
  wire [31:0] smul_75982;
  wire [31:0] smul_75983;
  wire [31:0] smul_75984;
  wire [31:0] add_75985;
  wire [31:0] add_75986;
  wire [31:0] smul_75987;
  wire [31:0] smul_75988;
  wire [31:0] smul_75989;
  wire [31:0] smul_75990;
  wire [31:0] smul_75991;
  wire [31:0] smul_75992;
  wire [31:0] add_75993;
  wire [31:0] add_75994;
  wire [31:0] smul_75995;
  wire [31:0] smul_75996;
  wire [31:0] smul_75997;
  wire [31:0] smul_75998;
  wire [31:0] smul_75999;
  wire [31:0] smul_76000;
  wire [31:0] add_76001;
  wire [31:0] add_76002;
  wire [31:0] smul_76003;
  wire [31:0] smul_76004;
  wire [31:0] smul_76005;
  wire [31:0] smul_76006;
  wire [31:0] smul_76007;
  wire [31:0] smul_76008;
  wire [31:0] add_76009;
  wire [31:0] add_76010;
  wire [31:0] smul_76011;
  wire [31:0] smul_76012;
  wire [31:0] smul_76013;
  wire [31:0] smul_76014;
  wire [31:0] smul_76015;
  wire [31:0] smul_76016;
  wire [31:0] add_76017;
  wire [31:0] add_76018;
  wire [31:0] smul_76019;
  wire [31:0] smul_76020;
  wire [31:0] smul_76021;
  wire [31:0] smul_76022;
  wire [31:0] smul_76023;
  wire [31:0] smul_76024;
  wire [31:0] add_76025;
  wire [31:0] add_76026;
  wire [31:0] smul_76027;
  wire [31:0] smul_76028;
  wire [31:0] smul_76029;
  wire [31:0] smul_76030;
  wire [31:0] smul_76031;
  wire [31:0] smul_76032;
  wire [31:0] add_76033;
  wire [31:0] add_76034;
  wire [31:0] smul_76035;
  wire [31:0] smul_76036;
  wire [31:0] smul_76037;
  wire [31:0] smul_76038;
  wire [31:0] smul_76039;
  wire [31:0] smul_76040;
  wire [31:0] add_76041;
  wire [31:0] add_76042;
  wire [31:0] smul_76043;
  wire [31:0] smul_76044;
  wire [31:0] smul_76045;
  wire [31:0] smul_76046;
  wire [31:0] smul_76047;
  wire [31:0] smul_76048;
  wire [31:0] add_76049;
  wire [31:0] add_76050;
  wire [31:0] smul_76051;
  wire [31:0] smul_76052;
  wire [31:0] smul_76053;
  wire [31:0] smul_76054;
  wire [31:0] smul_76055;
  wire [31:0] smul_76056;
  wire [31:0] add_76057;
  wire [31:0] add_76058;
  wire [31:0] smul_76059;
  wire [31:0] smul_76060;
  wire [31:0] smul_76061;
  wire [31:0] smul_76062;
  wire [31:0] smul_76063;
  wire [31:0] smul_76064;
  wire [31:0] add_76065;
  wire [31:0] add_76066;
  wire [31:0] smul_76067;
  wire [31:0] smul_76068;
  wire [31:0] smul_76069;
  wire [31:0] smul_76070;
  wire [31:0] smul_76071;
  wire [31:0] smul_76072;
  wire [31:0] add_76073;
  wire [31:0] add_76074;
  wire [31:0] smul_76075;
  wire [31:0] smul_76076;
  wire [31:0] smul_76077;
  wire [31:0] smul_76078;
  wire [31:0] smul_76079;
  wire [31:0] smul_76080;
  wire [31:0] add_76081;
  wire [31:0] add_76082;
  wire [31:0] smul_76083;
  wire [31:0] smul_76084;
  wire [31:0] smul_76085;
  wire [31:0] smul_76086;
  wire [31:0] smul_76087;
  wire [31:0] smul_76088;
  wire [31:0] add_76089;
  wire [31:0] add_76090;
  wire [31:0] smul_76091;
  wire [31:0] smul_76092;
  wire [31:0] smul_76093;
  wire [31:0] smul_76094;
  wire [31:0] smul_76095;
  wire [31:0] smul_76096;
  wire [31:0] add_76097;
  wire [31:0] add_76098;
  wire [31:0] smul_76099;
  wire [31:0] smul_76100;
  wire [31:0] smul_76101;
  wire [31:0] smul_76102;
  wire [31:0] smul_76103;
  wire [31:0] smul_76104;
  wire [31:0] add_76105;
  wire [31:0] add_76106;
  wire [31:0] smul_76107;
  wire [31:0] smul_76108;
  wire [31:0] smul_76109;
  wire [31:0] smul_76110;
  wire [31:0] smul_76111;
  wire [31:0] smul_76112;
  wire [31:0] add_76113;
  wire [31:0] add_76114;
  wire [31:0] smul_76115;
  wire [31:0] smul_76116;
  wire [31:0] smul_76117;
  wire [31:0] smul_76118;
  wire [31:0] smul_76119;
  wire [31:0] smul_76120;
  wire [31:0] add_76121;
  wire [31:0] add_76122;
  wire [31:0] smul_76123;
  wire [31:0] smul_76124;
  wire [31:0] smul_76125;
  wire [31:0] smul_76126;
  wire [31:0] smul_76127;
  wire [31:0] smul_76128;
  wire [31:0] add_76129;
  wire [31:0] add_76130;
  wire [31:0] smul_76131;
  wire [31:0] smul_76132;
  wire [31:0] smul_76133;
  wire [31:0] smul_76134;
  wire [31:0] smul_76135;
  wire [31:0] smul_76136;
  wire [31:0] add_76137;
  wire [31:0] add_76138;
  wire [31:0] smul_76139;
  wire [31:0] smul_76140;
  wire [31:0] smul_76141;
  wire [31:0] smul_76142;
  wire [31:0] smul_76143;
  wire [31:0] smul_76144;
  wire [31:0] add_76145;
  wire [31:0] add_76146;
  wire [31:0] smul_76147;
  wire [31:0] smul_76148;
  wire [31:0] smul_76149;
  wire [31:0] smul_76150;
  wire [31:0] smul_76151;
  wire [31:0] smul_76152;
  wire [31:0] add_76153;
  wire [31:0] add_76154;
  wire [31:0] smul_76155;
  wire [31:0] smul_76156;
  wire [31:0] smul_76157;
  wire [31:0] smul_76158;
  wire [31:0] smul_76159;
  wire [31:0] smul_76160;
  wire [31:0] add_76161;
  wire [31:0] add_76162;
  wire [31:0] smul_76163;
  wire [31:0] smul_76164;
  wire [31:0] smul_76165;
  wire [31:0] smul_76166;
  wire [31:0] smul_76167;
  wire [31:0] smul_76168;
  wire [31:0] add_76169;
  wire [31:0] add_76170;
  wire [31:0] smul_76171;
  wire [31:0] smul_76172;
  wire [31:0] smul_76173;
  wire [31:0] smul_76174;
  wire [31:0] smul_76175;
  wire [31:0] smul_76176;
  wire [31:0] add_76177;
  wire [31:0] add_76178;
  wire [31:0] smul_76179;
  wire [31:0] smul_76180;
  wire [31:0] smul_76181;
  wire [31:0] smul_76182;
  wire [31:0] smul_76183;
  wire [31:0] smul_76184;
  wire [31:0] add_76185;
  wire [31:0] add_76186;
  wire [31:0] smul_76187;
  wire [31:0] smul_76188;
  wire [31:0] smul_76189;
  wire [31:0] smul_76190;
  wire [31:0] smul_76191;
  wire [31:0] smul_76192;
  wire [31:0] add_76193;
  wire [31:0] add_76194;
  wire [31:0] smul_76195;
  wire [31:0] smul_76196;
  wire [31:0] smul_76197;
  wire [31:0] smul_76198;
  wire [31:0] smul_76199;
  wire [31:0] smul_76200;
  wire [31:0] add_76201;
  wire [31:0] add_76202;
  wire [31:0] smul_76203;
  wire [31:0] smul_76204;
  wire [31:0] smul_76205;
  wire [31:0] smul_76206;
  wire [31:0] smul_76207;
  wire [31:0] smul_76208;
  wire [31:0] add_76209;
  wire [31:0] add_76210;
  wire [31:0] smul_76211;
  wire [31:0] smul_76212;
  wire [31:0] smul_76213;
  wire [31:0] smul_76214;
  wire [31:0] smul_76215;
  wire [31:0] smul_76216;
  wire [31:0] add_76217;
  wire [31:0] add_76218;
  wire [31:0] smul_76219;
  wire [31:0] smul_76220;
  wire [31:0] smul_76221;
  wire [31:0] smul_76222;
  wire [31:0] smul_76223;
  wire [31:0] smul_76224;
  wire [31:0] add_76225;
  wire [31:0] add_76226;
  wire [31:0] smul_76227;
  wire [31:0] smul_76228;
  wire [31:0] smul_76229;
  wire [31:0] smul_76230;
  wire [31:0] smul_76231;
  wire [31:0] smul_76232;
  wire [31:0] add_76233;
  wire [31:0] add_76234;
  wire [31:0] smul_76235;
  wire [31:0] smul_76236;
  wire [31:0] smul_76237;
  wire [31:0] smul_76238;
  wire [31:0] smul_76239;
  wire [31:0] smul_76240;
  wire [31:0] add_76241;
  wire [31:0] add_76242;
  wire [31:0] smul_76243;
  wire [31:0] smul_76244;
  wire [31:0] smul_76245;
  wire [31:0] smul_76246;
  wire [31:0] smul_76247;
  wire [31:0] smul_76248;
  wire [31:0] add_76249;
  wire [31:0] add_76250;
  wire [31:0] smul_76251;
  wire [31:0] smul_76252;
  wire [31:0] smul_76253;
  wire [31:0] smul_76254;
  wire [31:0] smul_76255;
  wire [31:0] smul_76256;
  wire [31:0] add_76257;
  wire [31:0] add_76258;
  wire [31:0] smul_76259;
  wire [31:0] smul_76260;
  wire [31:0] smul_76261;
  wire [31:0] smul_76262;
  wire [31:0] smul_76263;
  wire [31:0] smul_76264;
  wire [31:0] add_76265;
  wire [31:0] add_76266;
  wire [31:0] smul_76267;
  wire [31:0] smul_76268;
  wire [31:0] smul_76269;
  wire [31:0] smul_76270;
  wire [31:0] smul_76271;
  wire [31:0] smul_76272;
  wire [31:0] add_76273;
  wire [31:0] add_76274;
  wire [31:0] smul_76275;
  wire [31:0] smul_76276;
  wire [31:0] smul_76277;
  wire [31:0] smul_76278;
  wire [31:0] smul_76279;
  wire [31:0] smul_76280;
  wire [31:0] add_76281;
  wire [31:0] add_76282;
  wire [31:0] smul_76283;
  wire [31:0] smul_76284;
  wire [31:0] smul_76285;
  wire [31:0] smul_76286;
  wire [31:0] smul_76287;
  wire [31:0] smul_76288;
  wire [31:0] add_76289;
  wire [31:0] add_76290;
  wire [31:0] smul_76291;
  wire [31:0] smul_76292;
  wire [31:0] smul_76293;
  wire [31:0] smul_76294;
  wire [31:0] smul_76295;
  wire [31:0] smul_76296;
  wire [31:0] add_76297;
  wire [31:0] add_76298;
  wire [31:0] smul_76299;
  wire [31:0] smul_76300;
  wire [31:0] smul_76301;
  wire [31:0] smul_76302;
  wire [31:0] smul_76303;
  wire [31:0] smul_76304;
  wire [31:0] add_76305;
  wire [31:0] add_76306;
  wire [31:0] smul_76307;
  wire [31:0] smul_76308;
  wire [31:0] smul_76309;
  wire [31:0] smul_76310;
  wire [31:0] smul_76311;
  wire [31:0] smul_76312;
  wire [31:0] add_76313;
  wire [31:0] add_76314;
  wire [31:0] smul_76315;
  wire [31:0] smul_76316;
  wire [31:0] smul_76317;
  wire [31:0] smul_76318;
  wire [31:0] smul_76319;
  wire [31:0] smul_76320;
  wire [31:0] add_76321;
  wire [31:0] add_76322;
  wire [31:0] smul_76323;
  wire [31:0] smul_76324;
  wire [31:0] smul_76325;
  wire [31:0] smul_76326;
  wire [31:0] smul_76327;
  wire [31:0] smul_76328;
  wire [31:0] add_76329;
  wire [31:0] add_76330;
  wire [31:0] smul_76331;
  wire [31:0] smul_76332;
  wire [31:0] smul_76333;
  wire [31:0] smul_76334;
  wire [31:0] smul_76335;
  wire [31:0] smul_76336;
  wire [31:0] add_76337;
  wire [31:0] add_76338;
  wire [31:0] smul_76339;
  wire [31:0] smul_76340;
  wire [31:0] smul_76341;
  wire [31:0] smul_76342;
  wire [31:0] smul_76343;
  wire [31:0] smul_76344;
  wire [31:0] add_76345;
  wire [31:0] add_76346;
  wire [31:0] smul_76347;
  wire [31:0] smul_76348;
  wire [31:0] smul_76349;
  wire [31:0] smul_76350;
  wire [31:0] smul_76351;
  wire [31:0] smul_76352;
  wire [31:0] add_76353;
  wire [31:0] add_76354;
  wire [31:0] smul_76355;
  wire [31:0] smul_76356;
  wire [31:0] smul_76357;
  wire [31:0] smul_76358;
  wire [31:0] smul_76359;
  wire [31:0] smul_76360;
  wire [31:0] add_76361;
  wire [31:0] add_76362;
  wire [31:0] smul_76363;
  wire [31:0] smul_76364;
  wire [31:0] smul_76365;
  wire [31:0] smul_76366;
  wire [31:0] smul_76367;
  wire [31:0] smul_76368;
  wire [31:0] add_76369;
  wire [31:0] add_76370;
  wire [31:0] smul_76371;
  wire [31:0] smul_76372;
  wire [31:0] smul_76373;
  wire [31:0] smul_76374;
  wire [31:0] smul_76375;
  wire [31:0] smul_76376;
  wire [31:0] add_76377;
  wire [31:0] add_76378;
  wire [31:0] smul_76379;
  wire [31:0] smul_76380;
  wire [31:0] smul_76381;
  wire [31:0] smul_76382;
  wire [31:0] smul_76383;
  wire [31:0] smul_76384;
  wire [31:0] add_76385;
  wire [31:0] add_76386;
  wire [31:0] smul_76387;
  wire [31:0] smul_76388;
  wire [31:0] smul_76389;
  wire [31:0] smul_76390;
  wire [31:0] smul_76391;
  wire [31:0] smul_76392;
  wire [31:0] add_76393;
  wire [31:0] add_76394;
  wire [31:0] smul_76395;
  wire [31:0] smul_76396;
  wire [31:0] smul_76397;
  wire [31:0] smul_76398;
  wire [31:0] smul_76399;
  wire [31:0] smul_76400;
  wire [31:0] add_76401;
  wire [31:0] add_76402;
  wire [31:0] smul_76403;
  wire [31:0] smul_76404;
  wire [31:0] smul_76405;
  wire [31:0] smul_76406;
  wire [31:0] smul_76407;
  wire [31:0] smul_76408;
  wire [31:0] add_76409;
  wire [31:0] add_76410;
  wire [31:0] smul_76411;
  wire [31:0] smul_76412;
  wire [31:0] smul_76413;
  wire [31:0] smul_76414;
  wire [31:0] smul_76415;
  wire [31:0] smul_76416;
  wire [31:0] add_76417;
  wire [31:0] add_76418;
  wire [31:0] smul_76419;
  wire [31:0] smul_76420;
  wire [31:0] smul_76421;
  wire [31:0] smul_76422;
  wire [31:0] smul_76423;
  wire [31:0] smul_76424;
  wire [31:0] add_76425;
  wire [31:0] add_76426;
  wire [31:0] smul_76427;
  wire [31:0] smul_76428;
  wire [31:0] smul_76429;
  wire [31:0] smul_76430;
  wire [31:0] smul_76431;
  wire [31:0] smul_76432;
  wire [31:0] add_76433;
  wire [31:0] add_76434;
  wire [31:0] smul_76435;
  wire [31:0] smul_76436;
  wire [31:0] smul_76437;
  wire [31:0] smul_76438;
  wire [31:0] smul_76439;
  wire [31:0] smul_76440;
  wire [31:0] add_76441;
  wire [31:0] add_76442;
  wire [31:0] smul_76443;
  wire [31:0] smul_76444;
  wire [31:0] smul_76445;
  wire [31:0] smul_76446;
  wire [31:0] smul_76447;
  wire [31:0] smul_76448;
  wire [31:0] add_76449;
  wire [31:0] add_76450;
  wire [31:0] smul_76451;
  wire [31:0] smul_76452;
  wire [31:0] smul_76453;
  wire [31:0] smul_76454;
  wire [31:0] smul_76455;
  wire [31:0] smul_76456;
  wire [31:0] add_76457;
  wire [31:0] add_76458;
  wire [31:0] smul_76459;
  wire [31:0] smul_76460;
  wire [31:0] smul_76461;
  wire [31:0] smul_76462;
  wire [31:0] smul_76463;
  wire [31:0] smul_76464;
  wire [31:0] add_76465;
  wire [31:0] add_76466;
  wire [31:0] smul_76467;
  wire [31:0] smul_76468;
  wire [31:0] smul_76469;
  wire [31:0] smul_76470;
  wire [31:0] smul_76471;
  wire [31:0] smul_76472;
  wire [31:0] add_76473;
  wire [31:0] add_76474;
  wire [31:0] add_76475;
  wire [31:0] add_76476;
  wire [31:0] add_76477;
  wire [31:0] add_76478;
  wire [31:0] add_76479;
  wire [31:0] add_76480;
  wire [31:0] add_76481;
  wire [31:0] add_76482;
  wire [31:0] add_76483;
  wire [31:0] add_76484;
  wire [31:0] add_76485;
  wire [31:0] add_76486;
  wire [31:0] add_76487;
  wire [31:0] add_76488;
  wire [31:0] add_76489;
  wire [31:0] add_76490;
  wire [31:0] add_76491;
  wire [31:0] add_76492;
  wire [31:0] add_76493;
  wire [31:0] add_76494;
  wire [31:0] add_76495;
  wire [31:0] add_76496;
  wire [31:0] add_76497;
  wire [31:0] add_76498;
  wire [31:0] add_76499;
  wire [31:0] add_76500;
  wire [31:0] add_76501;
  wire [31:0] add_76502;
  wire [31:0] add_76503;
  wire [31:0] add_76504;
  wire [31:0] add_76505;
  wire [31:0] add_76506;
  wire [31:0] add_76507;
  wire [31:0] add_76508;
  wire [31:0] add_76509;
  wire [31:0] add_76510;
  wire [31:0] add_76511;
  wire [31:0] add_76512;
  wire [31:0] add_76513;
  wire [31:0] add_76514;
  wire [31:0] add_76515;
  wire [31:0] add_76516;
  wire [31:0] add_76517;
  wire [31:0] add_76518;
  wire [31:0] add_76519;
  wire [31:0] add_76520;
  wire [31:0] add_76521;
  wire [31:0] add_76522;
  wire [31:0] add_76523;
  wire [31:0] add_76524;
  wire [31:0] add_76525;
  wire [31:0] add_76526;
  wire [31:0] add_76527;
  wire [31:0] add_76528;
  wire [31:0] add_76529;
  wire [31:0] add_76530;
  wire [31:0] add_76531;
  wire [31:0] add_76532;
  wire [31:0] add_76533;
  wire [31:0] add_76534;
  wire [31:0] add_76535;
  wire [31:0] add_76536;
  wire [31:0] add_76537;
  wire [31:0] add_76538;
  wire [31:0] add_76539;
  wire [31:0] add_76540;
  wire [31:0] add_76541;
  wire [31:0] add_76542;
  wire [31:0] add_76543;
  wire [31:0] add_76544;
  wire [31:0] add_76545;
  wire [31:0] add_76546;
  wire [31:0] add_76547;
  wire [31:0] add_76548;
  wire [31:0] add_76549;
  wire [31:0] add_76550;
  wire [31:0] add_76551;
  wire [31:0] add_76552;
  wire [31:0] add_76553;
  wire [31:0] add_76554;
  wire [31:0] add_76555;
  wire [31:0] add_76556;
  wire [31:0] add_76557;
  wire [31:0] add_76558;
  wire [31:0] add_76559;
  wire [31:0] add_76560;
  wire [31:0] add_76561;
  wire [31:0] add_76562;
  wire [31:0] add_76563;
  wire [31:0] add_76564;
  wire [31:0] add_76565;
  wire [31:0] add_76566;
  wire [31:0] add_76567;
  wire [31:0] add_76568;
  wire [31:0] add_76569;
  wire [31:0] add_76570;
  wire [31:0] add_76571;
  wire [31:0] add_76572;
  wire [31:0] add_76573;
  wire [31:0] add_76574;
  wire [31:0] add_76575;
  wire [31:0] add_76576;
  wire [31:0] add_76577;
  wire [31:0] add_76578;
  wire [31:0] add_76579;
  wire [31:0] add_76580;
  wire [31:0] add_76581;
  wire [31:0] add_76582;
  wire [31:0] add_76583;
  wire [31:0] add_76584;
  wire [31:0] add_76585;
  wire [31:0] add_76586;
  wire [31:0] add_76587;
  wire [31:0] add_76588;
  wire [31:0] add_76589;
  wire [31:0] add_76590;
  wire [31:0] add_76591;
  wire [31:0] add_76592;
  wire [31:0] add_76593;
  wire [31:0] add_76594;
  wire [31:0] add_76595;
  wire [31:0] add_76596;
  wire [31:0] add_76597;
  wire [31:0] add_76598;
  wire [31:0] add_76599;
  wire [31:0] add_76600;
  wire [31:0] add_76601;
  wire [31:0] add_76602;
  wire [31:0] add_76603;
  wire [31:0] add_76604;
  wire [31:0] add_76605;
  wire [31:0] add_76606;
  wire [31:0] add_76607;
  wire [31:0] add_76608;
  wire [31:0] add_76609;
  wire [31:0] add_76610;
  wire [31:0] add_76611;
  wire [31:0] add_76612;
  wire [31:0] add_76613;
  wire [31:0] add_76614;
  wire [31:0] add_76615;
  wire [31:0] add_76616;
  wire [31:0] add_76617;
  wire [31:0] add_76618;
  wire [31:0] add_76619;
  wire [31:0] add_76620;
  wire [31:0] add_76621;
  wire [31:0] add_76622;
  wire [31:0] add_76623;
  wire [31:0] add_76624;
  wire [31:0] add_76625;
  wire [31:0] add_76626;
  wire [31:0] add_76627;
  wire [31:0] add_76628;
  wire [31:0] add_76629;
  wire [31:0] add_76630;
  wire [31:0] add_76631;
  wire [31:0] add_76632;
  wire [31:0] add_76633;
  wire [31:0] add_76634;
  wire [31:0] add_76635;
  wire [31:0] add_76636;
  wire [31:0] add_76637;
  wire [31:0] add_76638;
  wire [31:0] add_76639;
  wire [31:0] add_76640;
  wire [31:0] add_76641;
  wire [31:0] add_76642;
  wire [31:0] add_76643;
  wire [31:0] add_76644;
  wire [31:0] add_76645;
  wire [31:0] add_76646;
  wire [31:0] add_76647;
  wire [31:0] add_76648;
  wire [31:0] add_76649;
  wire [31:0] add_76650;
  wire [31:0] add_76651;
  wire [31:0] add_76652;
  wire [31:0] add_76653;
  wire [31:0] add_76654;
  wire [31:0] add_76655;
  wire [31:0] add_76656;
  wire [31:0] add_76657;
  wire [31:0] add_76658;
  wire [31:0] add_76659;
  wire [31:0] add_76660;
  wire [31:0] add_76661;
  wire [31:0] add_76662;
  wire [31:0] add_76663;
  wire [31:0] add_76664;
  wire [31:0] add_76665;
  wire [31:0] add_76666;
  wire [31:0] add_76667;
  wire [31:0] add_76668;
  wire [31:0] add_76669;
  wire [31:0] add_76670;
  wire [31:0] add_76671;
  wire [31:0] add_76672;
  wire [31:0] add_76673;
  wire [31:0] add_76674;
  wire [31:0] add_76675;
  wire [31:0] add_76676;
  wire [31:0] add_76677;
  wire [31:0] add_76678;
  wire [31:0] add_76679;
  wire [31:0] add_76680;
  wire [31:0] add_76681;
  wire [31:0] add_76682;
  wire [31:0] add_76683;
  wire [31:0] add_76684;
  wire [31:0] add_76685;
  wire [31:0] add_76686;
  wire [31:0] add_76687;
  wire [31:0] add_76688;
  wire [31:0] add_76689;
  wire [31:0] add_76690;
  wire [31:0] add_76691;
  wire [31:0] add_76692;
  wire [31:0] add_76693;
  wire [31:0] add_76694;
  wire [31:0] add_76695;
  wire [31:0] add_76696;
  wire [31:0] add_76697;
  wire [31:0] add_76698;
  wire [31:0] add_76699;
  wire [31:0] add_76700;
  wire [31:0] add_76701;
  wire [31:0] add_76702;
  wire [31:0] add_76703;
  wire [31:0] add_76704;
  wire [31:0] add_76705;
  wire [31:0] add_76706;
  wire [31:0] add_76707;
  wire [31:0] add_76708;
  wire [31:0] add_76709;
  wire [31:0] add_76710;
  wire [31:0] add_76711;
  wire [31:0] add_76712;
  wire [31:0] add_76713;
  wire [31:0] add_76714;
  wire [31:0] add_76715;
  wire [31:0] add_76716;
  wire [31:0] add_76717;
  wire [31:0] add_76718;
  wire [31:0] add_76719;
  wire [31:0] add_76720;
  wire [31:0] add_76721;
  wire [31:0] add_76722;
  wire [31:0] add_76723;
  wire [31:0] add_76724;
  wire [31:0] add_76725;
  wire [31:0] add_76726;
  wire [31:0] add_76727;
  wire [31:0] add_76728;
  wire [31:0] add_76729;
  wire [31:0] add_76730;
  wire [31:0] add_76731;
  wire [31:0] add_76732;
  wire [31:0] add_76733;
  wire [31:0] add_76734;
  wire [31:0] add_76735;
  wire [31:0] add_76736;
  wire [31:0] add_76737;
  wire [31:0] add_76738;
  wire [31:0] add_76739;
  wire [31:0] add_76740;
  wire [31:0] add_76741;
  wire [31:0] add_76742;
  wire [31:0] add_76743;
  wire [31:0] add_76744;
  wire [31:0] add_76745;
  wire [31:0] add_76746;
  wire [31:0] add_76747;
  wire [31:0] add_76748;
  wire [31:0] add_76749;
  wire [31:0] add_76750;
  wire [31:0] add_76751;
  wire [31:0] add_76752;
  wire [31:0] add_76753;
  wire [31:0] add_76754;
  wire [31:0] add_76755;
  wire [31:0] add_76756;
  wire [31:0] add_76757;
  wire [31:0] add_76758;
  wire [31:0] add_76759;
  wire [31:0] add_76760;
  wire [31:0] add_76761;
  wire [31:0] add_76762;
  wire [31:0] add_76763;
  wire [31:0] add_76764;
  wire [31:0] add_76765;
  wire [31:0] add_76766;
  wire [31:0] add_76767;
  wire [31:0] add_76768;
  wire [31:0] add_76769;
  wire [31:0] add_76770;
  wire [31:0] add_76771;
  wire [31:0] add_76772;
  wire [31:0] add_76773;
  wire [31:0] add_76774;
  wire [31:0] add_76775;
  wire [31:0] add_76776;
  wire [31:0] add_76777;
  wire [31:0] add_76778;
  wire [31:0] add_76779;
  wire [31:0] add_76780;
  wire [31:0] add_76781;
  wire [31:0] add_76782;
  wire [31:0] add_76783;
  wire [31:0] add_76784;
  wire [31:0] add_76785;
  wire [31:0] add_76786;
  wire [31:0] add_76787;
  wire [31:0] add_76788;
  wire [31:0] add_76789;
  wire [31:0] add_76790;
  wire [31:0] add_76791;
  wire [31:0] add_76792;
  wire [31:0] add_76793;
  wire [31:0] add_76794;
  wire [31:0] add_76795;
  wire [31:0] add_76796;
  wire [31:0] add_76797;
  wire [31:0] add_76798;
  wire [31:0] add_76799;
  wire [31:0] add_76800;
  wire [31:0] add_76801;
  wire [31:0] add_76802;
  wire [31:0] add_76803;
  wire [31:0] add_76804;
  wire [31:0] add_76805;
  wire [31:0] add_76806;
  wire [31:0] add_76807;
  wire [31:0] add_76808;
  wire [31:0] add_76809;
  wire [31:0] add_76810;
  wire [31:0] add_76811;
  wire [31:0] add_76812;
  wire [31:0] add_76813;
  wire [31:0] add_76814;
  wire [31:0] add_76815;
  wire [31:0] add_76816;
  wire [31:0] add_76817;
  wire [31:0] add_76818;
  wire [31:0] add_76819;
  wire [31:0] add_76820;
  wire [31:0] add_76821;
  wire [31:0] add_76822;
  wire [31:0] add_76823;
  wire [31:0] add_76824;
  wire [31:0] add_76825;
  wire [31:0] add_76826;
  wire [31:0] add_76827;
  wire [31:0] add_76828;
  wire [31:0] add_76829;
  wire [31:0] add_76830;
  wire [31:0] add_76831;
  wire [31:0] add_76832;
  wire [31:0] add_76833;
  wire [31:0] add_76834;
  wire [31:0] add_76835;
  wire [31:0] add_76836;
  wire [31:0] add_76837;
  wire [31:0] add_76838;
  wire [31:0] add_76839;
  wire [31:0] add_76840;
  wire [31:0] add_76841;
  wire [31:0] add_76842;
  wire [31:0] add_76843;
  wire [31:0] add_76844;
  wire [31:0] add_76845;
  wire [31:0] add_76846;
  wire [31:0] add_76847;
  wire [31:0] add_76848;
  wire [31:0] add_76849;
  wire [31:0] add_76850;
  wire [31:0] add_76851;
  wire [31:0] add_76852;
  wire [31:0] add_76853;
  wire [31:0] add_76854;
  wire [31:0] add_76855;
  wire [31:0] add_76856;
  wire [31:0] add_76857;
  wire [31:0] add_76858;
  wire [31:0] add_76859;
  wire [31:0] add_76860;
  wire [31:0] add_76861;
  wire [31:0] add_76862;
  wire [31:0] add_76863;
  wire [31:0] add_76864;
  wire [31:0] add_76865;
  wire [31:0] add_76866;
  wire [31:0] add_76867;
  wire [31:0] add_76868;
  wire [31:0] add_76869;
  wire [31:0] add_76870;
  wire [31:0] add_76871;
  wire [31:0] add_76872;
  wire [31:0] add_76873;
  wire [31:0] add_76874;
  wire [31:0] add_76875;
  wire [31:0] add_76876;
  wire [31:0] add_76877;
  wire [31:0] add_76878;
  wire [31:0] add_76879;
  wire [31:0] add_76880;
  wire [31:0] add_76881;
  wire [31:0] add_76882;
  wire [31:0] add_76883;
  wire [31:0] add_76884;
  wire [31:0] add_76885;
  wire [31:0] add_76886;
  wire [31:0] add_76887;
  wire [31:0] add_76888;
  wire [31:0] add_76889;
  wire [31:0] add_76890;
  wire [31:0] add_76891;
  wire [31:0] add_76892;
  wire [31:0] add_76893;
  wire [31:0] add_76894;
  wire [31:0] add_76895;
  wire [31:0] add_76896;
  wire [31:0] add_76897;
  wire [31:0] add_76898;
  wire [31:0] add_76899;
  wire [31:0] add_76900;
  wire [31:0] add_76901;
  wire [31:0] add_76902;
  wire [31:0] add_76903;
  wire [31:0] add_76904;
  wire [31:0] add_76905;
  wire [31:0] add_76906;
  wire [31:0] add_76907;
  wire [31:0] add_76908;
  wire [31:0] add_76909;
  wire [31:0] add_76910;
  wire [31:0] add_76911;
  wire [31:0] add_76912;
  wire [31:0] add_76913;
  wire [31:0] add_76914;
  wire [31:0] add_76915;
  wire [31:0] add_76916;
  wire [31:0] add_76917;
  wire [31:0] add_76918;
  wire [31:0] add_76919;
  wire [31:0] add_76920;
  wire [31:0] add_76921;
  wire [31:0] add_76922;
  wire [31:0] add_76923;
  wire [31:0] add_76924;
  wire [31:0] add_76925;
  wire [31:0] add_76926;
  wire [31:0] add_76927;
  wire [31:0] add_76928;
  wire [31:0] add_76929;
  wire [31:0] add_76930;
  wire [31:0] add_76931;
  wire [31:0] add_76932;
  wire [31:0] add_76933;
  wire [31:0] add_76934;
  wire [31:0] add_76935;
  wire [31:0] add_76936;
  wire [31:0] add_76937;
  wire [31:0] add_76938;
  wire [31:0] add_76939;
  wire [31:0] add_76940;
  wire [31:0] add_76941;
  wire [31:0] add_76942;
  wire [31:0] add_76943;
  wire [31:0] add_76944;
  wire [31:0] add_76945;
  wire [31:0] add_76946;
  wire [31:0] add_76947;
  wire [31:0] add_76948;
  wire [31:0] add_76949;
  wire [31:0] add_76950;
  wire [31:0] add_76951;
  wire [31:0] add_76952;
  wire [31:0] add_76953;
  wire [31:0] add_76954;
  wire [31:0] add_76955;
  wire [31:0] add_76956;
  wire [31:0] add_76957;
  wire [31:0] add_76958;
  wire [31:0] add_76959;
  wire [31:0] add_76960;
  wire [31:0] add_76961;
  wire [31:0] add_76962;
  wire [31:0] add_76963;
  wire [31:0] add_76964;
  wire [31:0] add_76965;
  wire [31:0] add_76966;
  wire [31:0] add_76967;
  wire [31:0] add_76968;
  wire [31:0] add_76969;
  wire [31:0] add_76970;
  wire [31:0] add_76971;
  wire [31:0] add_76972;
  wire [31:0] add_76973;
  wire [31:0] add_76974;
  wire [31:0] add_76975;
  wire [31:0] add_76976;
  wire [31:0] add_76977;
  wire [31:0] add_76978;
  wire [31:0] add_76979;
  wire [31:0] add_76980;
  wire [31:0] add_76981;
  wire [31:0] add_76982;
  wire [31:0] add_76983;
  wire [31:0] add_76984;
  wire [31:0] add_76985;
  wire [31:0] add_76986;
  wire [31:0] add_76987;
  wire [31:0] add_76988;
  wire [31:0] add_76989;
  wire [31:0] add_76990;
  wire [31:0] add_76991;
  wire [31:0] add_76992;
  wire [31:0] add_76993;
  wire [31:0] add_76994;
  wire [31:0] add_76995;
  wire [31:0] add_76996;
  wire [31:0] add_76997;
  wire [31:0] add_76998;
  wire [31:0] add_76999;
  wire [31:0] add_77000;
  wire [31:0] add_77001;
  wire [31:0] add_77002;
  wire [31:0] add_77003;
  wire [31:0] add_77004;
  wire [31:0] add_77005;
  wire [31:0] add_77006;
  wire [31:0] add_77007;
  wire [31:0] add_77008;
  wire [31:0] add_77009;
  wire [31:0] add_77010;
  wire [31:0] add_77011;
  wire [31:0] add_77012;
  wire [31:0] add_77013;
  wire [31:0] add_77014;
  wire [31:0] add_77015;
  wire [31:0] add_77016;
  wire [31:0] add_77017;
  wire [31:0] add_77018;
  wire [31:0] add_77019;
  wire [31:0] add_77020;
  wire [31:0] add_77021;
  wire [31:0] add_77022;
  wire [31:0] add_77023;
  wire [31:0] add_77024;
  wire [31:0] add_77025;
  wire [31:0] add_77026;
  wire [31:0] add_77027;
  wire [31:0] add_77028;
  wire [31:0] add_77029;
  wire [31:0] add_77030;
  wire [31:0] add_77031;
  wire [31:0] add_77032;
  wire [31:0] add_77033;
  wire [31:0] add_77034;
  wire [31:0] add_77035;
  wire [31:0] add_77036;
  wire [31:0] add_77037;
  wire [31:0] add_77038;
  wire [31:0] add_77039;
  wire [31:0] add_77040;
  wire [31:0] add_77041;
  wire [31:0] add_77042;
  wire [31:0] add_77043;
  wire [31:0] add_77044;
  wire [31:0] add_77045;
  wire [31:0] add_77046;
  wire [31:0] add_77047;
  wire [31:0] add_77048;
  wire [31:0] add_77049;
  wire [31:0] add_77050;
  wire [31:0] add_77051;
  wire [31:0] add_77052;
  wire [31:0] add_77053;
  wire [31:0] add_77054;
  wire [31:0] add_77055;
  wire [31:0] add_77056;
  wire [31:0] add_77057;
  wire [31:0] add_77058;
  wire [31:0] add_77059;
  wire [31:0] add_77060;
  wire [31:0] add_77061;
  wire [31:0] add_77062;
  wire [31:0] add_77063;
  wire [31:0] add_77064;
  wire [31:0] add_77065;
  wire [31:0] add_77066;
  wire [31:0] add_77067;
  wire [31:0] add_77068;
  wire [31:0] add_77069;
  wire [31:0] add_77070;
  wire [31:0] add_77071;
  wire [31:0] add_77072;
  wire [31:0] add_77073;
  wire literal_77074;
  wire [31:0] add_77075;
  wire [31:0] add_77076;
  wire [31:0] add_77077;
  wire [31:0] add_77078;
  wire [31:0] add_77079;
  wire [31:0] add_77080;
  wire [31:0] add_77081;
  wire [31:0] add_77082;
  wire [31:0] add_77083;
  wire [31:0] add_77084;
  wire [31:0] add_77085;
  wire [31:0] add_77086;
  wire [31:0] add_77087;
  wire [31:0] add_77088;
  wire [31:0] add_77089;
  wire [31:0] add_77090;
  wire [31:0] add_77091;
  wire [31:0] add_77092;
  wire [31:0] add_77093;
  wire [31:0] add_77094;
  wire [31:0] add_77095;
  wire [31:0] add_77096;
  wire [31:0] add_77097;
  wire [31:0] add_77098;
  wire [31:0] add_77099;
  wire [31:0] add_77100;
  wire [31:0] add_77101;
  wire [31:0] add_77102;
  wire [31:0] add_77103;
  wire [31:0] add_77104;
  wire [31:0] add_77105;
  wire [31:0] add_77106;
  wire [31:0] add_77107;
  wire [31:0] add_77108;
  wire [31:0] add_77109;
  wire [31:0] add_77110;
  wire [31:0] add_77111;
  wire [31:0] add_77112;
  wire [31:0] add_77113;
  wire [31:0] add_77114;
  wire [31:0] add_77115;
  wire [31:0] add_77116;
  wire [31:0] add_77117;
  wire [31:0] add_77118;
  wire [31:0] add_77119;
  wire [31:0] add_77120;
  wire [31:0] add_77121;
  wire [31:0] add_77122;
  wire [31:0] add_77123;
  wire [31:0] add_77124;
  wire [31:0] add_77125;
  wire [31:0] add_77126;
  wire [31:0] add_77127;
  wire [31:0] add_77128;
  wire [31:0] add_77129;
  wire [31:0] add_77130;
  wire [31:0] add_77131;
  wire [31:0] add_77132;
  wire [31:0] add_77133;
  wire [31:0] add_77134;
  wire [31:0] add_77135;
  wire [31:0] add_77136;
  wire [31:0] add_77137;
  wire [31:0] add_77138;
  wire [31:0] add_77139;
  wire [31:0] add_77140;
  wire [31:0] add_77141;
  wire [31:0] add_77142;
  wire [31:0] add_77143;
  wire [31:0] add_77144;
  wire [31:0] add_77145;
  wire [31:0] add_77146;
  wire [31:0] add_77147;
  wire [31:0] add_77148;
  wire [31:0] add_77149;
  wire [31:0] add_77150;
  wire [31:0] add_77151;
  wire [31:0] add_77152;
  wire [31:0] add_77153;
  wire [31:0] add_77154;
  wire [31:0] add_77155;
  wire [31:0] add_77156;
  wire [31:0] add_77157;
  wire [31:0] add_77158;
  wire [31:0] add_77159;
  wire [31:0] add_77160;
  wire [31:0] add_77161;
  wire [31:0] add_77162;
  wire [31:0] add_77163;
  wire [31:0] add_77164;
  wire [31:0] add_77165;
  wire [31:0] add_77166;
  wire [31:0] add_77167;
  wire [31:0] add_77168;
  wire [31:0] add_77169;
  wire [31:0] add_77170;
  wire [31:0] add_77171;
  wire [31:0] add_77172;
  wire [31:0] add_77173;
  assign smul_75273 = smul32b_32b_x_32b(TestBlock__A_op0, TestBlock__B_op0);
  assign smul_75274 = smul32b_32b_x_32b(TestBlock__A_op1, TestBlock__B_op10);
  assign smul_75275 = smul32b_32b_x_32b(TestBlock__A_op2, TestBlock__B_op20);
  assign smul_75276 = smul32b_32b_x_32b(TestBlock__A_op3, TestBlock__B_op30);
  assign smul_75277 = smul32b_32b_x_32b(TestBlock__A_op0, TestBlock__B_op1);
  assign smul_75278 = smul32b_32b_x_32b(TestBlock__A_op1, TestBlock__B_op11);
  assign smul_75279 = smul32b_32b_x_32b(TestBlock__A_op2, TestBlock__B_op21);
  assign smul_75280 = smul32b_32b_x_32b(TestBlock__A_op3, TestBlock__B_op31);
  assign smul_75281 = smul32b_32b_x_32b(TestBlock__A_op0, TestBlock__B_op2);
  assign smul_75282 = smul32b_32b_x_32b(TestBlock__A_op1, TestBlock__B_op12);
  assign smul_75283 = smul32b_32b_x_32b(TestBlock__A_op2, TestBlock__B_op22);
  assign smul_75284 = smul32b_32b_x_32b(TestBlock__A_op3, TestBlock__B_op32);
  assign smul_75285 = smul32b_32b_x_32b(TestBlock__A_op0, TestBlock__B_op3);
  assign smul_75286 = smul32b_32b_x_32b(TestBlock__A_op1, TestBlock__B_op13);
  assign smul_75287 = smul32b_32b_x_32b(TestBlock__A_op2, TestBlock__B_op23);
  assign smul_75288 = smul32b_32b_x_32b(TestBlock__A_op3, TestBlock__B_op33);
  assign smul_75289 = smul32b_32b_x_32b(TestBlock__A_op0, TestBlock__B_op4);
  assign smul_75290 = smul32b_32b_x_32b(TestBlock__A_op1, TestBlock__B_op14);
  assign smul_75291 = smul32b_32b_x_32b(TestBlock__A_op2, TestBlock__B_op24);
  assign smul_75292 = smul32b_32b_x_32b(TestBlock__A_op3, TestBlock__B_op34);
  assign smul_75293 = smul32b_32b_x_32b(TestBlock__A_op0, TestBlock__B_op5);
  assign smul_75294 = smul32b_32b_x_32b(TestBlock__A_op1, TestBlock__B_op15);
  assign smul_75295 = smul32b_32b_x_32b(TestBlock__A_op2, TestBlock__B_op25);
  assign smul_75296 = smul32b_32b_x_32b(TestBlock__A_op3, TestBlock__B_op35);
  assign smul_75297 = smul32b_32b_x_32b(TestBlock__A_op0, TestBlock__B_op6);
  assign smul_75298 = smul32b_32b_x_32b(TestBlock__A_op1, TestBlock__B_op16);
  assign smul_75299 = smul32b_32b_x_32b(TestBlock__A_op2, TestBlock__B_op26);
  assign smul_75300 = smul32b_32b_x_32b(TestBlock__A_op3, TestBlock__B_op36);
  assign smul_75301 = smul32b_32b_x_32b(TestBlock__A_op0, TestBlock__B_op7);
  assign smul_75302 = smul32b_32b_x_32b(TestBlock__A_op1, TestBlock__B_op17);
  assign smul_75303 = smul32b_32b_x_32b(TestBlock__A_op2, TestBlock__B_op27);
  assign smul_75304 = smul32b_32b_x_32b(TestBlock__A_op3, TestBlock__B_op37);
  assign smul_75305 = smul32b_32b_x_32b(TestBlock__A_op0, TestBlock__B_op8);
  assign smul_75306 = smul32b_32b_x_32b(TestBlock__A_op1, TestBlock__B_op18);
  assign smul_75307 = smul32b_32b_x_32b(TestBlock__A_op2, TestBlock__B_op28);
  assign smul_75308 = smul32b_32b_x_32b(TestBlock__A_op3, TestBlock__B_op38);
  assign smul_75309 = smul32b_32b_x_32b(TestBlock__A_op0, TestBlock__B_op9);
  assign smul_75310 = smul32b_32b_x_32b(TestBlock__A_op1, TestBlock__B_op19);
  assign smul_75311 = smul32b_32b_x_32b(TestBlock__A_op2, TestBlock__B_op29);
  assign smul_75312 = smul32b_32b_x_32b(TestBlock__A_op3, TestBlock__B_op39);
  assign smul_75313 = smul32b_32b_x_32b(TestBlock__A_op10, TestBlock__B_op0);
  assign smul_75314 = smul32b_32b_x_32b(TestBlock__A_op11, TestBlock__B_op10);
  assign smul_75315 = smul32b_32b_x_32b(TestBlock__A_op12, TestBlock__B_op20);
  assign smul_75316 = smul32b_32b_x_32b(TestBlock__A_op13, TestBlock__B_op30);
  assign smul_75317 = smul32b_32b_x_32b(TestBlock__A_op10, TestBlock__B_op1);
  assign smul_75318 = smul32b_32b_x_32b(TestBlock__A_op11, TestBlock__B_op11);
  assign smul_75319 = smul32b_32b_x_32b(TestBlock__A_op12, TestBlock__B_op21);
  assign smul_75320 = smul32b_32b_x_32b(TestBlock__A_op13, TestBlock__B_op31);
  assign smul_75321 = smul32b_32b_x_32b(TestBlock__A_op10, TestBlock__B_op2);
  assign smul_75322 = smul32b_32b_x_32b(TestBlock__A_op11, TestBlock__B_op12);
  assign smul_75323 = smul32b_32b_x_32b(TestBlock__A_op12, TestBlock__B_op22);
  assign smul_75324 = smul32b_32b_x_32b(TestBlock__A_op13, TestBlock__B_op32);
  assign smul_75325 = smul32b_32b_x_32b(TestBlock__A_op10, TestBlock__B_op3);
  assign smul_75326 = smul32b_32b_x_32b(TestBlock__A_op11, TestBlock__B_op13);
  assign smul_75327 = smul32b_32b_x_32b(TestBlock__A_op12, TestBlock__B_op23);
  assign smul_75328 = smul32b_32b_x_32b(TestBlock__A_op13, TestBlock__B_op33);
  assign smul_75329 = smul32b_32b_x_32b(TestBlock__A_op10, TestBlock__B_op4);
  assign smul_75330 = smul32b_32b_x_32b(TestBlock__A_op11, TestBlock__B_op14);
  assign smul_75331 = smul32b_32b_x_32b(TestBlock__A_op12, TestBlock__B_op24);
  assign smul_75332 = smul32b_32b_x_32b(TestBlock__A_op13, TestBlock__B_op34);
  assign smul_75333 = smul32b_32b_x_32b(TestBlock__A_op10, TestBlock__B_op5);
  assign smul_75334 = smul32b_32b_x_32b(TestBlock__A_op11, TestBlock__B_op15);
  assign smul_75335 = smul32b_32b_x_32b(TestBlock__A_op12, TestBlock__B_op25);
  assign smul_75336 = smul32b_32b_x_32b(TestBlock__A_op13, TestBlock__B_op35);
  assign smul_75337 = smul32b_32b_x_32b(TestBlock__A_op10, TestBlock__B_op6);
  assign smul_75338 = smul32b_32b_x_32b(TestBlock__A_op11, TestBlock__B_op16);
  assign smul_75339 = smul32b_32b_x_32b(TestBlock__A_op12, TestBlock__B_op26);
  assign smul_75340 = smul32b_32b_x_32b(TestBlock__A_op13, TestBlock__B_op36);
  assign smul_75341 = smul32b_32b_x_32b(TestBlock__A_op10, TestBlock__B_op7);
  assign smul_75342 = smul32b_32b_x_32b(TestBlock__A_op11, TestBlock__B_op17);
  assign smul_75343 = smul32b_32b_x_32b(TestBlock__A_op12, TestBlock__B_op27);
  assign smul_75344 = smul32b_32b_x_32b(TestBlock__A_op13, TestBlock__B_op37);
  assign smul_75345 = smul32b_32b_x_32b(TestBlock__A_op10, TestBlock__B_op8);
  assign smul_75346 = smul32b_32b_x_32b(TestBlock__A_op11, TestBlock__B_op18);
  assign smul_75347 = smul32b_32b_x_32b(TestBlock__A_op12, TestBlock__B_op28);
  assign smul_75348 = smul32b_32b_x_32b(TestBlock__A_op13, TestBlock__B_op38);
  assign smul_75349 = smul32b_32b_x_32b(TestBlock__A_op10, TestBlock__B_op9);
  assign smul_75350 = smul32b_32b_x_32b(TestBlock__A_op11, TestBlock__B_op19);
  assign smul_75351 = smul32b_32b_x_32b(TestBlock__A_op12, TestBlock__B_op29);
  assign smul_75352 = smul32b_32b_x_32b(TestBlock__A_op13, TestBlock__B_op39);
  assign smul_75353 = smul32b_32b_x_32b(TestBlock__A_op20, TestBlock__B_op0);
  assign smul_75354 = smul32b_32b_x_32b(TestBlock__A_op21, TestBlock__B_op10);
  assign smul_75355 = smul32b_32b_x_32b(TestBlock__A_op22, TestBlock__B_op20);
  assign smul_75356 = smul32b_32b_x_32b(TestBlock__A_op23, TestBlock__B_op30);
  assign smul_75357 = smul32b_32b_x_32b(TestBlock__A_op20, TestBlock__B_op1);
  assign smul_75358 = smul32b_32b_x_32b(TestBlock__A_op21, TestBlock__B_op11);
  assign smul_75359 = smul32b_32b_x_32b(TestBlock__A_op22, TestBlock__B_op21);
  assign smul_75360 = smul32b_32b_x_32b(TestBlock__A_op23, TestBlock__B_op31);
  assign smul_75361 = smul32b_32b_x_32b(TestBlock__A_op20, TestBlock__B_op2);
  assign smul_75362 = smul32b_32b_x_32b(TestBlock__A_op21, TestBlock__B_op12);
  assign smul_75363 = smul32b_32b_x_32b(TestBlock__A_op22, TestBlock__B_op22);
  assign smul_75364 = smul32b_32b_x_32b(TestBlock__A_op23, TestBlock__B_op32);
  assign smul_75365 = smul32b_32b_x_32b(TestBlock__A_op20, TestBlock__B_op3);
  assign smul_75366 = smul32b_32b_x_32b(TestBlock__A_op21, TestBlock__B_op13);
  assign smul_75367 = smul32b_32b_x_32b(TestBlock__A_op22, TestBlock__B_op23);
  assign smul_75368 = smul32b_32b_x_32b(TestBlock__A_op23, TestBlock__B_op33);
  assign smul_75369 = smul32b_32b_x_32b(TestBlock__A_op20, TestBlock__B_op4);
  assign smul_75370 = smul32b_32b_x_32b(TestBlock__A_op21, TestBlock__B_op14);
  assign smul_75371 = smul32b_32b_x_32b(TestBlock__A_op22, TestBlock__B_op24);
  assign smul_75372 = smul32b_32b_x_32b(TestBlock__A_op23, TestBlock__B_op34);
  assign smul_75373 = smul32b_32b_x_32b(TestBlock__A_op20, TestBlock__B_op5);
  assign smul_75374 = smul32b_32b_x_32b(TestBlock__A_op21, TestBlock__B_op15);
  assign smul_75375 = smul32b_32b_x_32b(TestBlock__A_op22, TestBlock__B_op25);
  assign smul_75376 = smul32b_32b_x_32b(TestBlock__A_op23, TestBlock__B_op35);
  assign smul_75377 = smul32b_32b_x_32b(TestBlock__A_op20, TestBlock__B_op6);
  assign smul_75378 = smul32b_32b_x_32b(TestBlock__A_op21, TestBlock__B_op16);
  assign smul_75379 = smul32b_32b_x_32b(TestBlock__A_op22, TestBlock__B_op26);
  assign smul_75380 = smul32b_32b_x_32b(TestBlock__A_op23, TestBlock__B_op36);
  assign smul_75381 = smul32b_32b_x_32b(TestBlock__A_op20, TestBlock__B_op7);
  assign smul_75382 = smul32b_32b_x_32b(TestBlock__A_op21, TestBlock__B_op17);
  assign smul_75383 = smul32b_32b_x_32b(TestBlock__A_op22, TestBlock__B_op27);
  assign smul_75384 = smul32b_32b_x_32b(TestBlock__A_op23, TestBlock__B_op37);
  assign smul_75385 = smul32b_32b_x_32b(TestBlock__A_op20, TestBlock__B_op8);
  assign smul_75386 = smul32b_32b_x_32b(TestBlock__A_op21, TestBlock__B_op18);
  assign smul_75387 = smul32b_32b_x_32b(TestBlock__A_op22, TestBlock__B_op28);
  assign smul_75388 = smul32b_32b_x_32b(TestBlock__A_op23, TestBlock__B_op38);
  assign smul_75389 = smul32b_32b_x_32b(TestBlock__A_op20, TestBlock__B_op9);
  assign smul_75390 = smul32b_32b_x_32b(TestBlock__A_op21, TestBlock__B_op19);
  assign smul_75391 = smul32b_32b_x_32b(TestBlock__A_op22, TestBlock__B_op29);
  assign smul_75392 = smul32b_32b_x_32b(TestBlock__A_op23, TestBlock__B_op39);
  assign smul_75393 = smul32b_32b_x_32b(TestBlock__A_op30, TestBlock__B_op0);
  assign smul_75394 = smul32b_32b_x_32b(TestBlock__A_op31, TestBlock__B_op10);
  assign smul_75395 = smul32b_32b_x_32b(TestBlock__A_op32, TestBlock__B_op20);
  assign smul_75396 = smul32b_32b_x_32b(TestBlock__A_op33, TestBlock__B_op30);
  assign smul_75397 = smul32b_32b_x_32b(TestBlock__A_op30, TestBlock__B_op1);
  assign smul_75398 = smul32b_32b_x_32b(TestBlock__A_op31, TestBlock__B_op11);
  assign smul_75399 = smul32b_32b_x_32b(TestBlock__A_op32, TestBlock__B_op21);
  assign smul_75400 = smul32b_32b_x_32b(TestBlock__A_op33, TestBlock__B_op31);
  assign smul_75401 = smul32b_32b_x_32b(TestBlock__A_op30, TestBlock__B_op2);
  assign smul_75402 = smul32b_32b_x_32b(TestBlock__A_op31, TestBlock__B_op12);
  assign smul_75403 = smul32b_32b_x_32b(TestBlock__A_op32, TestBlock__B_op22);
  assign smul_75404 = smul32b_32b_x_32b(TestBlock__A_op33, TestBlock__B_op32);
  assign smul_75405 = smul32b_32b_x_32b(TestBlock__A_op30, TestBlock__B_op3);
  assign smul_75406 = smul32b_32b_x_32b(TestBlock__A_op31, TestBlock__B_op13);
  assign smul_75407 = smul32b_32b_x_32b(TestBlock__A_op32, TestBlock__B_op23);
  assign smul_75408 = smul32b_32b_x_32b(TestBlock__A_op33, TestBlock__B_op33);
  assign smul_75409 = smul32b_32b_x_32b(TestBlock__A_op30, TestBlock__B_op4);
  assign smul_75410 = smul32b_32b_x_32b(TestBlock__A_op31, TestBlock__B_op14);
  assign smul_75411 = smul32b_32b_x_32b(TestBlock__A_op32, TestBlock__B_op24);
  assign smul_75412 = smul32b_32b_x_32b(TestBlock__A_op33, TestBlock__B_op34);
  assign smul_75413 = smul32b_32b_x_32b(TestBlock__A_op30, TestBlock__B_op5);
  assign smul_75414 = smul32b_32b_x_32b(TestBlock__A_op31, TestBlock__B_op15);
  assign smul_75415 = smul32b_32b_x_32b(TestBlock__A_op32, TestBlock__B_op25);
  assign smul_75416 = smul32b_32b_x_32b(TestBlock__A_op33, TestBlock__B_op35);
  assign smul_75417 = smul32b_32b_x_32b(TestBlock__A_op30, TestBlock__B_op6);
  assign smul_75418 = smul32b_32b_x_32b(TestBlock__A_op31, TestBlock__B_op16);
  assign smul_75419 = smul32b_32b_x_32b(TestBlock__A_op32, TestBlock__B_op26);
  assign smul_75420 = smul32b_32b_x_32b(TestBlock__A_op33, TestBlock__B_op36);
  assign smul_75421 = smul32b_32b_x_32b(TestBlock__A_op30, TestBlock__B_op7);
  assign smul_75422 = smul32b_32b_x_32b(TestBlock__A_op31, TestBlock__B_op17);
  assign smul_75423 = smul32b_32b_x_32b(TestBlock__A_op32, TestBlock__B_op27);
  assign smul_75424 = smul32b_32b_x_32b(TestBlock__A_op33, TestBlock__B_op37);
  assign smul_75425 = smul32b_32b_x_32b(TestBlock__A_op30, TestBlock__B_op8);
  assign smul_75426 = smul32b_32b_x_32b(TestBlock__A_op31, TestBlock__B_op18);
  assign smul_75427 = smul32b_32b_x_32b(TestBlock__A_op32, TestBlock__B_op28);
  assign smul_75428 = smul32b_32b_x_32b(TestBlock__A_op33, TestBlock__B_op38);
  assign smul_75429 = smul32b_32b_x_32b(TestBlock__A_op30, TestBlock__B_op9);
  assign smul_75430 = smul32b_32b_x_32b(TestBlock__A_op31, TestBlock__B_op19);
  assign smul_75431 = smul32b_32b_x_32b(TestBlock__A_op32, TestBlock__B_op29);
  assign smul_75432 = smul32b_32b_x_32b(TestBlock__A_op33, TestBlock__B_op39);
  assign smul_75433 = smul32b_32b_x_32b(TestBlock__A_op40, TestBlock__B_op0);
  assign smul_75434 = smul32b_32b_x_32b(TestBlock__A_op41, TestBlock__B_op10);
  assign smul_75435 = smul32b_32b_x_32b(TestBlock__A_op42, TestBlock__B_op20);
  assign smul_75436 = smul32b_32b_x_32b(TestBlock__A_op43, TestBlock__B_op30);
  assign smul_75437 = smul32b_32b_x_32b(TestBlock__A_op40, TestBlock__B_op1);
  assign smul_75438 = smul32b_32b_x_32b(TestBlock__A_op41, TestBlock__B_op11);
  assign smul_75439 = smul32b_32b_x_32b(TestBlock__A_op42, TestBlock__B_op21);
  assign smul_75440 = smul32b_32b_x_32b(TestBlock__A_op43, TestBlock__B_op31);
  assign smul_75441 = smul32b_32b_x_32b(TestBlock__A_op40, TestBlock__B_op2);
  assign smul_75442 = smul32b_32b_x_32b(TestBlock__A_op41, TestBlock__B_op12);
  assign smul_75443 = smul32b_32b_x_32b(TestBlock__A_op42, TestBlock__B_op22);
  assign smul_75444 = smul32b_32b_x_32b(TestBlock__A_op43, TestBlock__B_op32);
  assign smul_75445 = smul32b_32b_x_32b(TestBlock__A_op40, TestBlock__B_op3);
  assign smul_75446 = smul32b_32b_x_32b(TestBlock__A_op41, TestBlock__B_op13);
  assign smul_75447 = smul32b_32b_x_32b(TestBlock__A_op42, TestBlock__B_op23);
  assign smul_75448 = smul32b_32b_x_32b(TestBlock__A_op43, TestBlock__B_op33);
  assign smul_75449 = smul32b_32b_x_32b(TestBlock__A_op40, TestBlock__B_op4);
  assign smul_75450 = smul32b_32b_x_32b(TestBlock__A_op41, TestBlock__B_op14);
  assign smul_75451 = smul32b_32b_x_32b(TestBlock__A_op42, TestBlock__B_op24);
  assign smul_75452 = smul32b_32b_x_32b(TestBlock__A_op43, TestBlock__B_op34);
  assign smul_75453 = smul32b_32b_x_32b(TestBlock__A_op40, TestBlock__B_op5);
  assign smul_75454 = smul32b_32b_x_32b(TestBlock__A_op41, TestBlock__B_op15);
  assign smul_75455 = smul32b_32b_x_32b(TestBlock__A_op42, TestBlock__B_op25);
  assign smul_75456 = smul32b_32b_x_32b(TestBlock__A_op43, TestBlock__B_op35);
  assign smul_75457 = smul32b_32b_x_32b(TestBlock__A_op40, TestBlock__B_op6);
  assign smul_75458 = smul32b_32b_x_32b(TestBlock__A_op41, TestBlock__B_op16);
  assign smul_75459 = smul32b_32b_x_32b(TestBlock__A_op42, TestBlock__B_op26);
  assign smul_75460 = smul32b_32b_x_32b(TestBlock__A_op43, TestBlock__B_op36);
  assign smul_75461 = smul32b_32b_x_32b(TestBlock__A_op40, TestBlock__B_op7);
  assign smul_75462 = smul32b_32b_x_32b(TestBlock__A_op41, TestBlock__B_op17);
  assign smul_75463 = smul32b_32b_x_32b(TestBlock__A_op42, TestBlock__B_op27);
  assign smul_75464 = smul32b_32b_x_32b(TestBlock__A_op43, TestBlock__B_op37);
  assign smul_75465 = smul32b_32b_x_32b(TestBlock__A_op40, TestBlock__B_op8);
  assign smul_75466 = smul32b_32b_x_32b(TestBlock__A_op41, TestBlock__B_op18);
  assign smul_75467 = smul32b_32b_x_32b(TestBlock__A_op42, TestBlock__B_op28);
  assign smul_75468 = smul32b_32b_x_32b(TestBlock__A_op43, TestBlock__B_op38);
  assign smul_75469 = smul32b_32b_x_32b(TestBlock__A_op40, TestBlock__B_op9);
  assign smul_75470 = smul32b_32b_x_32b(TestBlock__A_op41, TestBlock__B_op19);
  assign smul_75471 = smul32b_32b_x_32b(TestBlock__A_op42, TestBlock__B_op29);
  assign smul_75472 = smul32b_32b_x_32b(TestBlock__A_op43, TestBlock__B_op39);
  assign smul_75473 = smul32b_32b_x_32b(TestBlock__A_op50, TestBlock__B_op0);
  assign smul_75474 = smul32b_32b_x_32b(TestBlock__A_op51, TestBlock__B_op10);
  assign smul_75475 = smul32b_32b_x_32b(TestBlock__A_op52, TestBlock__B_op20);
  assign smul_75476 = smul32b_32b_x_32b(TestBlock__A_op53, TestBlock__B_op30);
  assign smul_75477 = smul32b_32b_x_32b(TestBlock__A_op50, TestBlock__B_op1);
  assign smul_75478 = smul32b_32b_x_32b(TestBlock__A_op51, TestBlock__B_op11);
  assign smul_75479 = smul32b_32b_x_32b(TestBlock__A_op52, TestBlock__B_op21);
  assign smul_75480 = smul32b_32b_x_32b(TestBlock__A_op53, TestBlock__B_op31);
  assign smul_75481 = smul32b_32b_x_32b(TestBlock__A_op50, TestBlock__B_op2);
  assign smul_75482 = smul32b_32b_x_32b(TestBlock__A_op51, TestBlock__B_op12);
  assign smul_75483 = smul32b_32b_x_32b(TestBlock__A_op52, TestBlock__B_op22);
  assign smul_75484 = smul32b_32b_x_32b(TestBlock__A_op53, TestBlock__B_op32);
  assign smul_75485 = smul32b_32b_x_32b(TestBlock__A_op50, TestBlock__B_op3);
  assign smul_75486 = smul32b_32b_x_32b(TestBlock__A_op51, TestBlock__B_op13);
  assign smul_75487 = smul32b_32b_x_32b(TestBlock__A_op52, TestBlock__B_op23);
  assign smul_75488 = smul32b_32b_x_32b(TestBlock__A_op53, TestBlock__B_op33);
  assign smul_75489 = smul32b_32b_x_32b(TestBlock__A_op50, TestBlock__B_op4);
  assign smul_75490 = smul32b_32b_x_32b(TestBlock__A_op51, TestBlock__B_op14);
  assign smul_75491 = smul32b_32b_x_32b(TestBlock__A_op52, TestBlock__B_op24);
  assign smul_75492 = smul32b_32b_x_32b(TestBlock__A_op53, TestBlock__B_op34);
  assign smul_75493 = smul32b_32b_x_32b(TestBlock__A_op50, TestBlock__B_op5);
  assign smul_75494 = smul32b_32b_x_32b(TestBlock__A_op51, TestBlock__B_op15);
  assign smul_75495 = smul32b_32b_x_32b(TestBlock__A_op52, TestBlock__B_op25);
  assign smul_75496 = smul32b_32b_x_32b(TestBlock__A_op53, TestBlock__B_op35);
  assign smul_75497 = smul32b_32b_x_32b(TestBlock__A_op50, TestBlock__B_op6);
  assign smul_75498 = smul32b_32b_x_32b(TestBlock__A_op51, TestBlock__B_op16);
  assign smul_75499 = smul32b_32b_x_32b(TestBlock__A_op52, TestBlock__B_op26);
  assign smul_75500 = smul32b_32b_x_32b(TestBlock__A_op53, TestBlock__B_op36);
  assign smul_75501 = smul32b_32b_x_32b(TestBlock__A_op50, TestBlock__B_op7);
  assign smul_75502 = smul32b_32b_x_32b(TestBlock__A_op51, TestBlock__B_op17);
  assign smul_75503 = smul32b_32b_x_32b(TestBlock__A_op52, TestBlock__B_op27);
  assign smul_75504 = smul32b_32b_x_32b(TestBlock__A_op53, TestBlock__B_op37);
  assign smul_75505 = smul32b_32b_x_32b(TestBlock__A_op50, TestBlock__B_op8);
  assign smul_75506 = smul32b_32b_x_32b(TestBlock__A_op51, TestBlock__B_op18);
  assign smul_75507 = smul32b_32b_x_32b(TestBlock__A_op52, TestBlock__B_op28);
  assign smul_75508 = smul32b_32b_x_32b(TestBlock__A_op53, TestBlock__B_op38);
  assign smul_75509 = smul32b_32b_x_32b(TestBlock__A_op50, TestBlock__B_op9);
  assign smul_75510 = smul32b_32b_x_32b(TestBlock__A_op51, TestBlock__B_op19);
  assign smul_75511 = smul32b_32b_x_32b(TestBlock__A_op52, TestBlock__B_op29);
  assign smul_75512 = smul32b_32b_x_32b(TestBlock__A_op53, TestBlock__B_op39);
  assign smul_75513 = smul32b_32b_x_32b(TestBlock__A_op60, TestBlock__B_op0);
  assign smul_75514 = smul32b_32b_x_32b(TestBlock__A_op61, TestBlock__B_op10);
  assign smul_75515 = smul32b_32b_x_32b(TestBlock__A_op62, TestBlock__B_op20);
  assign smul_75516 = smul32b_32b_x_32b(TestBlock__A_op63, TestBlock__B_op30);
  assign smul_75517 = smul32b_32b_x_32b(TestBlock__A_op60, TestBlock__B_op1);
  assign smul_75518 = smul32b_32b_x_32b(TestBlock__A_op61, TestBlock__B_op11);
  assign smul_75519 = smul32b_32b_x_32b(TestBlock__A_op62, TestBlock__B_op21);
  assign smul_75520 = smul32b_32b_x_32b(TestBlock__A_op63, TestBlock__B_op31);
  assign smul_75521 = smul32b_32b_x_32b(TestBlock__A_op60, TestBlock__B_op2);
  assign smul_75522 = smul32b_32b_x_32b(TestBlock__A_op61, TestBlock__B_op12);
  assign smul_75523 = smul32b_32b_x_32b(TestBlock__A_op62, TestBlock__B_op22);
  assign smul_75524 = smul32b_32b_x_32b(TestBlock__A_op63, TestBlock__B_op32);
  assign smul_75525 = smul32b_32b_x_32b(TestBlock__A_op60, TestBlock__B_op3);
  assign smul_75526 = smul32b_32b_x_32b(TestBlock__A_op61, TestBlock__B_op13);
  assign smul_75527 = smul32b_32b_x_32b(TestBlock__A_op62, TestBlock__B_op23);
  assign smul_75528 = smul32b_32b_x_32b(TestBlock__A_op63, TestBlock__B_op33);
  assign smul_75529 = smul32b_32b_x_32b(TestBlock__A_op60, TestBlock__B_op4);
  assign smul_75530 = smul32b_32b_x_32b(TestBlock__A_op61, TestBlock__B_op14);
  assign smul_75531 = smul32b_32b_x_32b(TestBlock__A_op62, TestBlock__B_op24);
  assign smul_75532 = smul32b_32b_x_32b(TestBlock__A_op63, TestBlock__B_op34);
  assign smul_75533 = smul32b_32b_x_32b(TestBlock__A_op60, TestBlock__B_op5);
  assign smul_75534 = smul32b_32b_x_32b(TestBlock__A_op61, TestBlock__B_op15);
  assign smul_75535 = smul32b_32b_x_32b(TestBlock__A_op62, TestBlock__B_op25);
  assign smul_75536 = smul32b_32b_x_32b(TestBlock__A_op63, TestBlock__B_op35);
  assign smul_75537 = smul32b_32b_x_32b(TestBlock__A_op60, TestBlock__B_op6);
  assign smul_75538 = smul32b_32b_x_32b(TestBlock__A_op61, TestBlock__B_op16);
  assign smul_75539 = smul32b_32b_x_32b(TestBlock__A_op62, TestBlock__B_op26);
  assign smul_75540 = smul32b_32b_x_32b(TestBlock__A_op63, TestBlock__B_op36);
  assign smul_75541 = smul32b_32b_x_32b(TestBlock__A_op60, TestBlock__B_op7);
  assign smul_75542 = smul32b_32b_x_32b(TestBlock__A_op61, TestBlock__B_op17);
  assign smul_75543 = smul32b_32b_x_32b(TestBlock__A_op62, TestBlock__B_op27);
  assign smul_75544 = smul32b_32b_x_32b(TestBlock__A_op63, TestBlock__B_op37);
  assign smul_75545 = smul32b_32b_x_32b(TestBlock__A_op60, TestBlock__B_op8);
  assign smul_75546 = smul32b_32b_x_32b(TestBlock__A_op61, TestBlock__B_op18);
  assign smul_75547 = smul32b_32b_x_32b(TestBlock__A_op62, TestBlock__B_op28);
  assign smul_75548 = smul32b_32b_x_32b(TestBlock__A_op63, TestBlock__B_op38);
  assign smul_75549 = smul32b_32b_x_32b(TestBlock__A_op60, TestBlock__B_op9);
  assign smul_75550 = smul32b_32b_x_32b(TestBlock__A_op61, TestBlock__B_op19);
  assign smul_75551 = smul32b_32b_x_32b(TestBlock__A_op62, TestBlock__B_op29);
  assign smul_75552 = smul32b_32b_x_32b(TestBlock__A_op63, TestBlock__B_op39);
  assign smul_75553 = smul32b_32b_x_32b(TestBlock__A_op70, TestBlock__B_op0);
  assign smul_75554 = smul32b_32b_x_32b(TestBlock__A_op71, TestBlock__B_op10);
  assign smul_75555 = smul32b_32b_x_32b(TestBlock__A_op72, TestBlock__B_op20);
  assign smul_75556 = smul32b_32b_x_32b(TestBlock__A_op73, TestBlock__B_op30);
  assign smul_75557 = smul32b_32b_x_32b(TestBlock__A_op70, TestBlock__B_op1);
  assign smul_75558 = smul32b_32b_x_32b(TestBlock__A_op71, TestBlock__B_op11);
  assign smul_75559 = smul32b_32b_x_32b(TestBlock__A_op72, TestBlock__B_op21);
  assign smul_75560 = smul32b_32b_x_32b(TestBlock__A_op73, TestBlock__B_op31);
  assign smul_75561 = smul32b_32b_x_32b(TestBlock__A_op70, TestBlock__B_op2);
  assign smul_75562 = smul32b_32b_x_32b(TestBlock__A_op71, TestBlock__B_op12);
  assign smul_75563 = smul32b_32b_x_32b(TestBlock__A_op72, TestBlock__B_op22);
  assign smul_75564 = smul32b_32b_x_32b(TestBlock__A_op73, TestBlock__B_op32);
  assign smul_75565 = smul32b_32b_x_32b(TestBlock__A_op70, TestBlock__B_op3);
  assign smul_75566 = smul32b_32b_x_32b(TestBlock__A_op71, TestBlock__B_op13);
  assign smul_75567 = smul32b_32b_x_32b(TestBlock__A_op72, TestBlock__B_op23);
  assign smul_75568 = smul32b_32b_x_32b(TestBlock__A_op73, TestBlock__B_op33);
  assign smul_75569 = smul32b_32b_x_32b(TestBlock__A_op70, TestBlock__B_op4);
  assign smul_75570 = smul32b_32b_x_32b(TestBlock__A_op71, TestBlock__B_op14);
  assign smul_75571 = smul32b_32b_x_32b(TestBlock__A_op72, TestBlock__B_op24);
  assign smul_75572 = smul32b_32b_x_32b(TestBlock__A_op73, TestBlock__B_op34);
  assign smul_75573 = smul32b_32b_x_32b(TestBlock__A_op70, TestBlock__B_op5);
  assign smul_75574 = smul32b_32b_x_32b(TestBlock__A_op71, TestBlock__B_op15);
  assign smul_75575 = smul32b_32b_x_32b(TestBlock__A_op72, TestBlock__B_op25);
  assign smul_75576 = smul32b_32b_x_32b(TestBlock__A_op73, TestBlock__B_op35);
  assign smul_75577 = smul32b_32b_x_32b(TestBlock__A_op70, TestBlock__B_op6);
  assign smul_75578 = smul32b_32b_x_32b(TestBlock__A_op71, TestBlock__B_op16);
  assign smul_75579 = smul32b_32b_x_32b(TestBlock__A_op72, TestBlock__B_op26);
  assign smul_75580 = smul32b_32b_x_32b(TestBlock__A_op73, TestBlock__B_op36);
  assign smul_75581 = smul32b_32b_x_32b(TestBlock__A_op70, TestBlock__B_op7);
  assign smul_75582 = smul32b_32b_x_32b(TestBlock__A_op71, TestBlock__B_op17);
  assign smul_75583 = smul32b_32b_x_32b(TestBlock__A_op72, TestBlock__B_op27);
  assign smul_75584 = smul32b_32b_x_32b(TestBlock__A_op73, TestBlock__B_op37);
  assign smul_75585 = smul32b_32b_x_32b(TestBlock__A_op70, TestBlock__B_op8);
  assign smul_75586 = smul32b_32b_x_32b(TestBlock__A_op71, TestBlock__B_op18);
  assign smul_75587 = smul32b_32b_x_32b(TestBlock__A_op72, TestBlock__B_op28);
  assign smul_75588 = smul32b_32b_x_32b(TestBlock__A_op73, TestBlock__B_op38);
  assign smul_75589 = smul32b_32b_x_32b(TestBlock__A_op70, TestBlock__B_op9);
  assign smul_75590 = smul32b_32b_x_32b(TestBlock__A_op71, TestBlock__B_op19);
  assign smul_75591 = smul32b_32b_x_32b(TestBlock__A_op72, TestBlock__B_op29);
  assign smul_75592 = smul32b_32b_x_32b(TestBlock__A_op73, TestBlock__B_op39);
  assign smul_75593 = smul32b_32b_x_32b(TestBlock__A_op80, TestBlock__B_op0);
  assign smul_75594 = smul32b_32b_x_32b(TestBlock__A_op81, TestBlock__B_op10);
  assign smul_75595 = smul32b_32b_x_32b(TestBlock__A_op82, TestBlock__B_op20);
  assign smul_75596 = smul32b_32b_x_32b(TestBlock__A_op83, TestBlock__B_op30);
  assign smul_75597 = smul32b_32b_x_32b(TestBlock__A_op80, TestBlock__B_op1);
  assign smul_75598 = smul32b_32b_x_32b(TestBlock__A_op81, TestBlock__B_op11);
  assign smul_75599 = smul32b_32b_x_32b(TestBlock__A_op82, TestBlock__B_op21);
  assign smul_75600 = smul32b_32b_x_32b(TestBlock__A_op83, TestBlock__B_op31);
  assign smul_75601 = smul32b_32b_x_32b(TestBlock__A_op80, TestBlock__B_op2);
  assign smul_75602 = smul32b_32b_x_32b(TestBlock__A_op81, TestBlock__B_op12);
  assign smul_75603 = smul32b_32b_x_32b(TestBlock__A_op82, TestBlock__B_op22);
  assign smul_75604 = smul32b_32b_x_32b(TestBlock__A_op83, TestBlock__B_op32);
  assign smul_75605 = smul32b_32b_x_32b(TestBlock__A_op80, TestBlock__B_op3);
  assign smul_75606 = smul32b_32b_x_32b(TestBlock__A_op81, TestBlock__B_op13);
  assign smul_75607 = smul32b_32b_x_32b(TestBlock__A_op82, TestBlock__B_op23);
  assign smul_75608 = smul32b_32b_x_32b(TestBlock__A_op83, TestBlock__B_op33);
  assign smul_75609 = smul32b_32b_x_32b(TestBlock__A_op80, TestBlock__B_op4);
  assign smul_75610 = smul32b_32b_x_32b(TestBlock__A_op81, TestBlock__B_op14);
  assign smul_75611 = smul32b_32b_x_32b(TestBlock__A_op82, TestBlock__B_op24);
  assign smul_75612 = smul32b_32b_x_32b(TestBlock__A_op83, TestBlock__B_op34);
  assign smul_75613 = smul32b_32b_x_32b(TestBlock__A_op80, TestBlock__B_op5);
  assign smul_75614 = smul32b_32b_x_32b(TestBlock__A_op81, TestBlock__B_op15);
  assign smul_75615 = smul32b_32b_x_32b(TestBlock__A_op82, TestBlock__B_op25);
  assign smul_75616 = smul32b_32b_x_32b(TestBlock__A_op83, TestBlock__B_op35);
  assign smul_75617 = smul32b_32b_x_32b(TestBlock__A_op80, TestBlock__B_op6);
  assign smul_75618 = smul32b_32b_x_32b(TestBlock__A_op81, TestBlock__B_op16);
  assign smul_75619 = smul32b_32b_x_32b(TestBlock__A_op82, TestBlock__B_op26);
  assign smul_75620 = smul32b_32b_x_32b(TestBlock__A_op83, TestBlock__B_op36);
  assign smul_75621 = smul32b_32b_x_32b(TestBlock__A_op80, TestBlock__B_op7);
  assign smul_75622 = smul32b_32b_x_32b(TestBlock__A_op81, TestBlock__B_op17);
  assign smul_75623 = smul32b_32b_x_32b(TestBlock__A_op82, TestBlock__B_op27);
  assign smul_75624 = smul32b_32b_x_32b(TestBlock__A_op83, TestBlock__B_op37);
  assign smul_75625 = smul32b_32b_x_32b(TestBlock__A_op80, TestBlock__B_op8);
  assign smul_75626 = smul32b_32b_x_32b(TestBlock__A_op81, TestBlock__B_op18);
  assign smul_75627 = smul32b_32b_x_32b(TestBlock__A_op82, TestBlock__B_op28);
  assign smul_75628 = smul32b_32b_x_32b(TestBlock__A_op83, TestBlock__B_op38);
  assign smul_75629 = smul32b_32b_x_32b(TestBlock__A_op80, TestBlock__B_op9);
  assign smul_75630 = smul32b_32b_x_32b(TestBlock__A_op81, TestBlock__B_op19);
  assign smul_75631 = smul32b_32b_x_32b(TestBlock__A_op82, TestBlock__B_op29);
  assign smul_75632 = smul32b_32b_x_32b(TestBlock__A_op83, TestBlock__B_op39);
  assign smul_75633 = smul32b_32b_x_32b(TestBlock__A_op90, TestBlock__B_op0);
  assign smul_75634 = smul32b_32b_x_32b(TestBlock__A_op91, TestBlock__B_op10);
  assign smul_75635 = smul32b_32b_x_32b(TestBlock__A_op92, TestBlock__B_op20);
  assign smul_75636 = smul32b_32b_x_32b(TestBlock__A_op93, TestBlock__B_op30);
  assign smul_75637 = smul32b_32b_x_32b(TestBlock__A_op90, TestBlock__B_op1);
  assign smul_75638 = smul32b_32b_x_32b(TestBlock__A_op91, TestBlock__B_op11);
  assign smul_75639 = smul32b_32b_x_32b(TestBlock__A_op92, TestBlock__B_op21);
  assign smul_75640 = smul32b_32b_x_32b(TestBlock__A_op93, TestBlock__B_op31);
  assign smul_75641 = smul32b_32b_x_32b(TestBlock__A_op90, TestBlock__B_op2);
  assign smul_75642 = smul32b_32b_x_32b(TestBlock__A_op91, TestBlock__B_op12);
  assign smul_75643 = smul32b_32b_x_32b(TestBlock__A_op92, TestBlock__B_op22);
  assign smul_75644 = smul32b_32b_x_32b(TestBlock__A_op93, TestBlock__B_op32);
  assign smul_75645 = smul32b_32b_x_32b(TestBlock__A_op90, TestBlock__B_op3);
  assign smul_75646 = smul32b_32b_x_32b(TestBlock__A_op91, TestBlock__B_op13);
  assign smul_75647 = smul32b_32b_x_32b(TestBlock__A_op92, TestBlock__B_op23);
  assign smul_75648 = smul32b_32b_x_32b(TestBlock__A_op93, TestBlock__B_op33);
  assign smul_75649 = smul32b_32b_x_32b(TestBlock__A_op90, TestBlock__B_op4);
  assign smul_75650 = smul32b_32b_x_32b(TestBlock__A_op91, TestBlock__B_op14);
  assign smul_75651 = smul32b_32b_x_32b(TestBlock__A_op92, TestBlock__B_op24);
  assign smul_75652 = smul32b_32b_x_32b(TestBlock__A_op93, TestBlock__B_op34);
  assign smul_75653 = smul32b_32b_x_32b(TestBlock__A_op90, TestBlock__B_op5);
  assign smul_75654 = smul32b_32b_x_32b(TestBlock__A_op91, TestBlock__B_op15);
  assign smul_75655 = smul32b_32b_x_32b(TestBlock__A_op92, TestBlock__B_op25);
  assign smul_75656 = smul32b_32b_x_32b(TestBlock__A_op93, TestBlock__B_op35);
  assign smul_75657 = smul32b_32b_x_32b(TestBlock__A_op90, TestBlock__B_op6);
  assign smul_75658 = smul32b_32b_x_32b(TestBlock__A_op91, TestBlock__B_op16);
  assign smul_75659 = smul32b_32b_x_32b(TestBlock__A_op92, TestBlock__B_op26);
  assign smul_75660 = smul32b_32b_x_32b(TestBlock__A_op93, TestBlock__B_op36);
  assign smul_75661 = smul32b_32b_x_32b(TestBlock__A_op90, TestBlock__B_op7);
  assign smul_75662 = smul32b_32b_x_32b(TestBlock__A_op91, TestBlock__B_op17);
  assign smul_75663 = smul32b_32b_x_32b(TestBlock__A_op92, TestBlock__B_op27);
  assign smul_75664 = smul32b_32b_x_32b(TestBlock__A_op93, TestBlock__B_op37);
  assign smul_75665 = smul32b_32b_x_32b(TestBlock__A_op90, TestBlock__B_op8);
  assign smul_75666 = smul32b_32b_x_32b(TestBlock__A_op91, TestBlock__B_op18);
  assign smul_75667 = smul32b_32b_x_32b(TestBlock__A_op92, TestBlock__B_op28);
  assign smul_75668 = smul32b_32b_x_32b(TestBlock__A_op93, TestBlock__B_op38);
  assign smul_75669 = smul32b_32b_x_32b(TestBlock__A_op90, TestBlock__B_op9);
  assign smul_75670 = smul32b_32b_x_32b(TestBlock__A_op91, TestBlock__B_op19);
  assign smul_75671 = smul32b_32b_x_32b(TestBlock__A_op92, TestBlock__B_op29);
  assign smul_75672 = smul32b_32b_x_32b(TestBlock__A_op93, TestBlock__B_op39);
  assign add_75673 = smul_75273 + smul_75274;
  assign add_75674 = smul_75275 + smul_75276;
  assign smul_75675 = smul32b_32b_x_32b(TestBlock__A_op4, TestBlock__B_op40);
  assign smul_75676 = smul32b_32b_x_32b(TestBlock__A_op5, TestBlock__B_op50);
  assign smul_75677 = smul32b_32b_x_32b(TestBlock__A_op6, TestBlock__B_op60);
  assign smul_75678 = smul32b_32b_x_32b(TestBlock__A_op7, TestBlock__B_op70);
  assign smul_75679 = smul32b_32b_x_32b(TestBlock__A_op8, TestBlock__B_op80);
  assign smul_75680 = smul32b_32b_x_32b(TestBlock__A_op9, TestBlock__B_op90);
  assign add_75681 = smul_75277 + smul_75278;
  assign add_75682 = smul_75279 + smul_75280;
  assign smul_75683 = smul32b_32b_x_32b(TestBlock__A_op4, TestBlock__B_op41);
  assign smul_75684 = smul32b_32b_x_32b(TestBlock__A_op5, TestBlock__B_op51);
  assign smul_75685 = smul32b_32b_x_32b(TestBlock__A_op6, TestBlock__B_op61);
  assign smul_75686 = smul32b_32b_x_32b(TestBlock__A_op7, TestBlock__B_op71);
  assign smul_75687 = smul32b_32b_x_32b(TestBlock__A_op8, TestBlock__B_op81);
  assign smul_75688 = smul32b_32b_x_32b(TestBlock__A_op9, TestBlock__B_op91);
  assign add_75689 = smul_75281 + smul_75282;
  assign add_75690 = smul_75283 + smul_75284;
  assign smul_75691 = smul32b_32b_x_32b(TestBlock__A_op4, TestBlock__B_op42);
  assign smul_75692 = smul32b_32b_x_32b(TestBlock__A_op5, TestBlock__B_op52);
  assign smul_75693 = smul32b_32b_x_32b(TestBlock__A_op6, TestBlock__B_op62);
  assign smul_75694 = smul32b_32b_x_32b(TestBlock__A_op7, TestBlock__B_op72);
  assign smul_75695 = smul32b_32b_x_32b(TestBlock__A_op8, TestBlock__B_op82);
  assign smul_75696 = smul32b_32b_x_32b(TestBlock__A_op9, TestBlock__B_op92);
  assign add_75697 = smul_75285 + smul_75286;
  assign add_75698 = smul_75287 + smul_75288;
  assign smul_75699 = smul32b_32b_x_32b(TestBlock__A_op4, TestBlock__B_op43);
  assign smul_75700 = smul32b_32b_x_32b(TestBlock__A_op5, TestBlock__B_op53);
  assign smul_75701 = smul32b_32b_x_32b(TestBlock__A_op6, TestBlock__B_op63);
  assign smul_75702 = smul32b_32b_x_32b(TestBlock__A_op7, TestBlock__B_op73);
  assign smul_75703 = smul32b_32b_x_32b(TestBlock__A_op8, TestBlock__B_op83);
  assign smul_75704 = smul32b_32b_x_32b(TestBlock__A_op9, TestBlock__B_op93);
  assign add_75705 = smul_75289 + smul_75290;
  assign add_75706 = smul_75291 + smul_75292;
  assign smul_75707 = smul32b_32b_x_32b(TestBlock__A_op4, TestBlock__B_op44);
  assign smul_75708 = smul32b_32b_x_32b(TestBlock__A_op5, TestBlock__B_op54);
  assign smul_75709 = smul32b_32b_x_32b(TestBlock__A_op6, TestBlock__B_op64);
  assign smul_75710 = smul32b_32b_x_32b(TestBlock__A_op7, TestBlock__B_op74);
  assign smul_75711 = smul32b_32b_x_32b(TestBlock__A_op8, TestBlock__B_op84);
  assign smul_75712 = smul32b_32b_x_32b(TestBlock__A_op9, TestBlock__B_op94);
  assign add_75713 = smul_75293 + smul_75294;
  assign add_75714 = smul_75295 + smul_75296;
  assign smul_75715 = smul32b_32b_x_32b(TestBlock__A_op4, TestBlock__B_op45);
  assign smul_75716 = smul32b_32b_x_32b(TestBlock__A_op5, TestBlock__B_op55);
  assign smul_75717 = smul32b_32b_x_32b(TestBlock__A_op6, TestBlock__B_op65);
  assign smul_75718 = smul32b_32b_x_32b(TestBlock__A_op7, TestBlock__B_op75);
  assign smul_75719 = smul32b_32b_x_32b(TestBlock__A_op8, TestBlock__B_op85);
  assign smul_75720 = smul32b_32b_x_32b(TestBlock__A_op9, TestBlock__B_op95);
  assign add_75721 = smul_75297 + smul_75298;
  assign add_75722 = smul_75299 + smul_75300;
  assign smul_75723 = smul32b_32b_x_32b(TestBlock__A_op4, TestBlock__B_op46);
  assign smul_75724 = smul32b_32b_x_32b(TestBlock__A_op5, TestBlock__B_op56);
  assign smul_75725 = smul32b_32b_x_32b(TestBlock__A_op6, TestBlock__B_op66);
  assign smul_75726 = smul32b_32b_x_32b(TestBlock__A_op7, TestBlock__B_op76);
  assign smul_75727 = smul32b_32b_x_32b(TestBlock__A_op8, TestBlock__B_op86);
  assign smul_75728 = smul32b_32b_x_32b(TestBlock__A_op9, TestBlock__B_op96);
  assign add_75729 = smul_75301 + smul_75302;
  assign add_75730 = smul_75303 + smul_75304;
  assign smul_75731 = smul32b_32b_x_32b(TestBlock__A_op4, TestBlock__B_op47);
  assign smul_75732 = smul32b_32b_x_32b(TestBlock__A_op5, TestBlock__B_op57);
  assign smul_75733 = smul32b_32b_x_32b(TestBlock__A_op6, TestBlock__B_op67);
  assign smul_75734 = smul32b_32b_x_32b(TestBlock__A_op7, TestBlock__B_op77);
  assign smul_75735 = smul32b_32b_x_32b(TestBlock__A_op8, TestBlock__B_op87);
  assign smul_75736 = smul32b_32b_x_32b(TestBlock__A_op9, TestBlock__B_op97);
  assign add_75737 = smul_75305 + smul_75306;
  assign add_75738 = smul_75307 + smul_75308;
  assign smul_75739 = smul32b_32b_x_32b(TestBlock__A_op4, TestBlock__B_op48);
  assign smul_75740 = smul32b_32b_x_32b(TestBlock__A_op5, TestBlock__B_op58);
  assign smul_75741 = smul32b_32b_x_32b(TestBlock__A_op6, TestBlock__B_op68);
  assign smul_75742 = smul32b_32b_x_32b(TestBlock__A_op7, TestBlock__B_op78);
  assign smul_75743 = smul32b_32b_x_32b(TestBlock__A_op8, TestBlock__B_op88);
  assign smul_75744 = smul32b_32b_x_32b(TestBlock__A_op9, TestBlock__B_op98);
  assign add_75745 = smul_75309 + smul_75310;
  assign add_75746 = smul_75311 + smul_75312;
  assign smul_75747 = smul32b_32b_x_32b(TestBlock__A_op4, TestBlock__B_op49);
  assign smul_75748 = smul32b_32b_x_32b(TestBlock__A_op5, TestBlock__B_op59);
  assign smul_75749 = smul32b_32b_x_32b(TestBlock__A_op6, TestBlock__B_op69);
  assign smul_75750 = smul32b_32b_x_32b(TestBlock__A_op7, TestBlock__B_op79);
  assign smul_75751 = smul32b_32b_x_32b(TestBlock__A_op8, TestBlock__B_op89);
  assign smul_75752 = smul32b_32b_x_32b(TestBlock__A_op9, TestBlock__B_op99);
  assign add_75753 = smul_75313 + smul_75314;
  assign add_75754 = smul_75315 + smul_75316;
  assign smul_75755 = smul32b_32b_x_32b(TestBlock__A_op14, TestBlock__B_op40);
  assign smul_75756 = smul32b_32b_x_32b(TestBlock__A_op15, TestBlock__B_op50);
  assign smul_75757 = smul32b_32b_x_32b(TestBlock__A_op16, TestBlock__B_op60);
  assign smul_75758 = smul32b_32b_x_32b(TestBlock__A_op17, TestBlock__B_op70);
  assign smul_75759 = smul32b_32b_x_32b(TestBlock__A_op18, TestBlock__B_op80);
  assign smul_75760 = smul32b_32b_x_32b(TestBlock__A_op19, TestBlock__B_op90);
  assign add_75761 = smul_75317 + smul_75318;
  assign add_75762 = smul_75319 + smul_75320;
  assign smul_75763 = smul32b_32b_x_32b(TestBlock__A_op14, TestBlock__B_op41);
  assign smul_75764 = smul32b_32b_x_32b(TestBlock__A_op15, TestBlock__B_op51);
  assign smul_75765 = smul32b_32b_x_32b(TestBlock__A_op16, TestBlock__B_op61);
  assign smul_75766 = smul32b_32b_x_32b(TestBlock__A_op17, TestBlock__B_op71);
  assign smul_75767 = smul32b_32b_x_32b(TestBlock__A_op18, TestBlock__B_op81);
  assign smul_75768 = smul32b_32b_x_32b(TestBlock__A_op19, TestBlock__B_op91);
  assign add_75769 = smul_75321 + smul_75322;
  assign add_75770 = smul_75323 + smul_75324;
  assign smul_75771 = smul32b_32b_x_32b(TestBlock__A_op14, TestBlock__B_op42);
  assign smul_75772 = smul32b_32b_x_32b(TestBlock__A_op15, TestBlock__B_op52);
  assign smul_75773 = smul32b_32b_x_32b(TestBlock__A_op16, TestBlock__B_op62);
  assign smul_75774 = smul32b_32b_x_32b(TestBlock__A_op17, TestBlock__B_op72);
  assign smul_75775 = smul32b_32b_x_32b(TestBlock__A_op18, TestBlock__B_op82);
  assign smul_75776 = smul32b_32b_x_32b(TestBlock__A_op19, TestBlock__B_op92);
  assign add_75777 = smul_75325 + smul_75326;
  assign add_75778 = smul_75327 + smul_75328;
  assign smul_75779 = smul32b_32b_x_32b(TestBlock__A_op14, TestBlock__B_op43);
  assign smul_75780 = smul32b_32b_x_32b(TestBlock__A_op15, TestBlock__B_op53);
  assign smul_75781 = smul32b_32b_x_32b(TestBlock__A_op16, TestBlock__B_op63);
  assign smul_75782 = smul32b_32b_x_32b(TestBlock__A_op17, TestBlock__B_op73);
  assign smul_75783 = smul32b_32b_x_32b(TestBlock__A_op18, TestBlock__B_op83);
  assign smul_75784 = smul32b_32b_x_32b(TestBlock__A_op19, TestBlock__B_op93);
  assign add_75785 = smul_75329 + smul_75330;
  assign add_75786 = smul_75331 + smul_75332;
  assign smul_75787 = smul32b_32b_x_32b(TestBlock__A_op14, TestBlock__B_op44);
  assign smul_75788 = smul32b_32b_x_32b(TestBlock__A_op15, TestBlock__B_op54);
  assign smul_75789 = smul32b_32b_x_32b(TestBlock__A_op16, TestBlock__B_op64);
  assign smul_75790 = smul32b_32b_x_32b(TestBlock__A_op17, TestBlock__B_op74);
  assign smul_75791 = smul32b_32b_x_32b(TestBlock__A_op18, TestBlock__B_op84);
  assign smul_75792 = smul32b_32b_x_32b(TestBlock__A_op19, TestBlock__B_op94);
  assign add_75793 = smul_75333 + smul_75334;
  assign add_75794 = smul_75335 + smul_75336;
  assign smul_75795 = smul32b_32b_x_32b(TestBlock__A_op14, TestBlock__B_op45);
  assign smul_75796 = smul32b_32b_x_32b(TestBlock__A_op15, TestBlock__B_op55);
  assign smul_75797 = smul32b_32b_x_32b(TestBlock__A_op16, TestBlock__B_op65);
  assign smul_75798 = smul32b_32b_x_32b(TestBlock__A_op17, TestBlock__B_op75);
  assign smul_75799 = smul32b_32b_x_32b(TestBlock__A_op18, TestBlock__B_op85);
  assign smul_75800 = smul32b_32b_x_32b(TestBlock__A_op19, TestBlock__B_op95);
  assign add_75801 = smul_75337 + smul_75338;
  assign add_75802 = smul_75339 + smul_75340;
  assign smul_75803 = smul32b_32b_x_32b(TestBlock__A_op14, TestBlock__B_op46);
  assign smul_75804 = smul32b_32b_x_32b(TestBlock__A_op15, TestBlock__B_op56);
  assign smul_75805 = smul32b_32b_x_32b(TestBlock__A_op16, TestBlock__B_op66);
  assign smul_75806 = smul32b_32b_x_32b(TestBlock__A_op17, TestBlock__B_op76);
  assign smul_75807 = smul32b_32b_x_32b(TestBlock__A_op18, TestBlock__B_op86);
  assign smul_75808 = smul32b_32b_x_32b(TestBlock__A_op19, TestBlock__B_op96);
  assign add_75809 = smul_75341 + smul_75342;
  assign add_75810 = smul_75343 + smul_75344;
  assign smul_75811 = smul32b_32b_x_32b(TestBlock__A_op14, TestBlock__B_op47);
  assign smul_75812 = smul32b_32b_x_32b(TestBlock__A_op15, TestBlock__B_op57);
  assign smul_75813 = smul32b_32b_x_32b(TestBlock__A_op16, TestBlock__B_op67);
  assign smul_75814 = smul32b_32b_x_32b(TestBlock__A_op17, TestBlock__B_op77);
  assign smul_75815 = smul32b_32b_x_32b(TestBlock__A_op18, TestBlock__B_op87);
  assign smul_75816 = smul32b_32b_x_32b(TestBlock__A_op19, TestBlock__B_op97);
  assign add_75817 = smul_75345 + smul_75346;
  assign add_75818 = smul_75347 + smul_75348;
  assign smul_75819 = smul32b_32b_x_32b(TestBlock__A_op14, TestBlock__B_op48);
  assign smul_75820 = smul32b_32b_x_32b(TestBlock__A_op15, TestBlock__B_op58);
  assign smul_75821 = smul32b_32b_x_32b(TestBlock__A_op16, TestBlock__B_op68);
  assign smul_75822 = smul32b_32b_x_32b(TestBlock__A_op17, TestBlock__B_op78);
  assign smul_75823 = smul32b_32b_x_32b(TestBlock__A_op18, TestBlock__B_op88);
  assign smul_75824 = smul32b_32b_x_32b(TestBlock__A_op19, TestBlock__B_op98);
  assign add_75825 = smul_75349 + smul_75350;
  assign add_75826 = smul_75351 + smul_75352;
  assign smul_75827 = smul32b_32b_x_32b(TestBlock__A_op14, TestBlock__B_op49);
  assign smul_75828 = smul32b_32b_x_32b(TestBlock__A_op15, TestBlock__B_op59);
  assign smul_75829 = smul32b_32b_x_32b(TestBlock__A_op16, TestBlock__B_op69);
  assign smul_75830 = smul32b_32b_x_32b(TestBlock__A_op17, TestBlock__B_op79);
  assign smul_75831 = smul32b_32b_x_32b(TestBlock__A_op18, TestBlock__B_op89);
  assign smul_75832 = smul32b_32b_x_32b(TestBlock__A_op19, TestBlock__B_op99);
  assign add_75833 = smul_75353 + smul_75354;
  assign add_75834 = smul_75355 + smul_75356;
  assign smul_75835 = smul32b_32b_x_32b(TestBlock__A_op24, TestBlock__B_op40);
  assign smul_75836 = smul32b_32b_x_32b(TestBlock__A_op25, TestBlock__B_op50);
  assign smul_75837 = smul32b_32b_x_32b(TestBlock__A_op26, TestBlock__B_op60);
  assign smul_75838 = smul32b_32b_x_32b(TestBlock__A_op27, TestBlock__B_op70);
  assign smul_75839 = smul32b_32b_x_32b(TestBlock__A_op28, TestBlock__B_op80);
  assign smul_75840 = smul32b_32b_x_32b(TestBlock__A_op29, TestBlock__B_op90);
  assign add_75841 = smul_75357 + smul_75358;
  assign add_75842 = smul_75359 + smul_75360;
  assign smul_75843 = smul32b_32b_x_32b(TestBlock__A_op24, TestBlock__B_op41);
  assign smul_75844 = smul32b_32b_x_32b(TestBlock__A_op25, TestBlock__B_op51);
  assign smul_75845 = smul32b_32b_x_32b(TestBlock__A_op26, TestBlock__B_op61);
  assign smul_75846 = smul32b_32b_x_32b(TestBlock__A_op27, TestBlock__B_op71);
  assign smul_75847 = smul32b_32b_x_32b(TestBlock__A_op28, TestBlock__B_op81);
  assign smul_75848 = smul32b_32b_x_32b(TestBlock__A_op29, TestBlock__B_op91);
  assign add_75849 = smul_75361 + smul_75362;
  assign add_75850 = smul_75363 + smul_75364;
  assign smul_75851 = smul32b_32b_x_32b(TestBlock__A_op24, TestBlock__B_op42);
  assign smul_75852 = smul32b_32b_x_32b(TestBlock__A_op25, TestBlock__B_op52);
  assign smul_75853 = smul32b_32b_x_32b(TestBlock__A_op26, TestBlock__B_op62);
  assign smul_75854 = smul32b_32b_x_32b(TestBlock__A_op27, TestBlock__B_op72);
  assign smul_75855 = smul32b_32b_x_32b(TestBlock__A_op28, TestBlock__B_op82);
  assign smul_75856 = smul32b_32b_x_32b(TestBlock__A_op29, TestBlock__B_op92);
  assign add_75857 = smul_75365 + smul_75366;
  assign add_75858 = smul_75367 + smul_75368;
  assign smul_75859 = smul32b_32b_x_32b(TestBlock__A_op24, TestBlock__B_op43);
  assign smul_75860 = smul32b_32b_x_32b(TestBlock__A_op25, TestBlock__B_op53);
  assign smul_75861 = smul32b_32b_x_32b(TestBlock__A_op26, TestBlock__B_op63);
  assign smul_75862 = smul32b_32b_x_32b(TestBlock__A_op27, TestBlock__B_op73);
  assign smul_75863 = smul32b_32b_x_32b(TestBlock__A_op28, TestBlock__B_op83);
  assign smul_75864 = smul32b_32b_x_32b(TestBlock__A_op29, TestBlock__B_op93);
  assign add_75865 = smul_75369 + smul_75370;
  assign add_75866 = smul_75371 + smul_75372;
  assign smul_75867 = smul32b_32b_x_32b(TestBlock__A_op24, TestBlock__B_op44);
  assign smul_75868 = smul32b_32b_x_32b(TestBlock__A_op25, TestBlock__B_op54);
  assign smul_75869 = smul32b_32b_x_32b(TestBlock__A_op26, TestBlock__B_op64);
  assign smul_75870 = smul32b_32b_x_32b(TestBlock__A_op27, TestBlock__B_op74);
  assign smul_75871 = smul32b_32b_x_32b(TestBlock__A_op28, TestBlock__B_op84);
  assign smul_75872 = smul32b_32b_x_32b(TestBlock__A_op29, TestBlock__B_op94);
  assign add_75873 = smul_75373 + smul_75374;
  assign add_75874 = smul_75375 + smul_75376;
  assign smul_75875 = smul32b_32b_x_32b(TestBlock__A_op24, TestBlock__B_op45);
  assign smul_75876 = smul32b_32b_x_32b(TestBlock__A_op25, TestBlock__B_op55);
  assign smul_75877 = smul32b_32b_x_32b(TestBlock__A_op26, TestBlock__B_op65);
  assign smul_75878 = smul32b_32b_x_32b(TestBlock__A_op27, TestBlock__B_op75);
  assign smul_75879 = smul32b_32b_x_32b(TestBlock__A_op28, TestBlock__B_op85);
  assign smul_75880 = smul32b_32b_x_32b(TestBlock__A_op29, TestBlock__B_op95);
  assign add_75881 = smul_75377 + smul_75378;
  assign add_75882 = smul_75379 + smul_75380;
  assign smul_75883 = smul32b_32b_x_32b(TestBlock__A_op24, TestBlock__B_op46);
  assign smul_75884 = smul32b_32b_x_32b(TestBlock__A_op25, TestBlock__B_op56);
  assign smul_75885 = smul32b_32b_x_32b(TestBlock__A_op26, TestBlock__B_op66);
  assign smul_75886 = smul32b_32b_x_32b(TestBlock__A_op27, TestBlock__B_op76);
  assign smul_75887 = smul32b_32b_x_32b(TestBlock__A_op28, TestBlock__B_op86);
  assign smul_75888 = smul32b_32b_x_32b(TestBlock__A_op29, TestBlock__B_op96);
  assign add_75889 = smul_75381 + smul_75382;
  assign add_75890 = smul_75383 + smul_75384;
  assign smul_75891 = smul32b_32b_x_32b(TestBlock__A_op24, TestBlock__B_op47);
  assign smul_75892 = smul32b_32b_x_32b(TestBlock__A_op25, TestBlock__B_op57);
  assign smul_75893 = smul32b_32b_x_32b(TestBlock__A_op26, TestBlock__B_op67);
  assign smul_75894 = smul32b_32b_x_32b(TestBlock__A_op27, TestBlock__B_op77);
  assign smul_75895 = smul32b_32b_x_32b(TestBlock__A_op28, TestBlock__B_op87);
  assign smul_75896 = smul32b_32b_x_32b(TestBlock__A_op29, TestBlock__B_op97);
  assign add_75897 = smul_75385 + smul_75386;
  assign add_75898 = smul_75387 + smul_75388;
  assign smul_75899 = smul32b_32b_x_32b(TestBlock__A_op24, TestBlock__B_op48);
  assign smul_75900 = smul32b_32b_x_32b(TestBlock__A_op25, TestBlock__B_op58);
  assign smul_75901 = smul32b_32b_x_32b(TestBlock__A_op26, TestBlock__B_op68);
  assign smul_75902 = smul32b_32b_x_32b(TestBlock__A_op27, TestBlock__B_op78);
  assign smul_75903 = smul32b_32b_x_32b(TestBlock__A_op28, TestBlock__B_op88);
  assign smul_75904 = smul32b_32b_x_32b(TestBlock__A_op29, TestBlock__B_op98);
  assign add_75905 = smul_75389 + smul_75390;
  assign add_75906 = smul_75391 + smul_75392;
  assign smul_75907 = smul32b_32b_x_32b(TestBlock__A_op24, TestBlock__B_op49);
  assign smul_75908 = smul32b_32b_x_32b(TestBlock__A_op25, TestBlock__B_op59);
  assign smul_75909 = smul32b_32b_x_32b(TestBlock__A_op26, TestBlock__B_op69);
  assign smul_75910 = smul32b_32b_x_32b(TestBlock__A_op27, TestBlock__B_op79);
  assign smul_75911 = smul32b_32b_x_32b(TestBlock__A_op28, TestBlock__B_op89);
  assign smul_75912 = smul32b_32b_x_32b(TestBlock__A_op29, TestBlock__B_op99);
  assign add_75913 = smul_75393 + smul_75394;
  assign add_75914 = smul_75395 + smul_75396;
  assign smul_75915 = smul32b_32b_x_32b(TestBlock__A_op34, TestBlock__B_op40);
  assign smul_75916 = smul32b_32b_x_32b(TestBlock__A_op35, TestBlock__B_op50);
  assign smul_75917 = smul32b_32b_x_32b(TestBlock__A_op36, TestBlock__B_op60);
  assign smul_75918 = smul32b_32b_x_32b(TestBlock__A_op37, TestBlock__B_op70);
  assign smul_75919 = smul32b_32b_x_32b(TestBlock__A_op38, TestBlock__B_op80);
  assign smul_75920 = smul32b_32b_x_32b(TestBlock__A_op39, TestBlock__B_op90);
  assign add_75921 = smul_75397 + smul_75398;
  assign add_75922 = smul_75399 + smul_75400;
  assign smul_75923 = smul32b_32b_x_32b(TestBlock__A_op34, TestBlock__B_op41);
  assign smul_75924 = smul32b_32b_x_32b(TestBlock__A_op35, TestBlock__B_op51);
  assign smul_75925 = smul32b_32b_x_32b(TestBlock__A_op36, TestBlock__B_op61);
  assign smul_75926 = smul32b_32b_x_32b(TestBlock__A_op37, TestBlock__B_op71);
  assign smul_75927 = smul32b_32b_x_32b(TestBlock__A_op38, TestBlock__B_op81);
  assign smul_75928 = smul32b_32b_x_32b(TestBlock__A_op39, TestBlock__B_op91);
  assign add_75929 = smul_75401 + smul_75402;
  assign add_75930 = smul_75403 + smul_75404;
  assign smul_75931 = smul32b_32b_x_32b(TestBlock__A_op34, TestBlock__B_op42);
  assign smul_75932 = smul32b_32b_x_32b(TestBlock__A_op35, TestBlock__B_op52);
  assign smul_75933 = smul32b_32b_x_32b(TestBlock__A_op36, TestBlock__B_op62);
  assign smul_75934 = smul32b_32b_x_32b(TestBlock__A_op37, TestBlock__B_op72);
  assign smul_75935 = smul32b_32b_x_32b(TestBlock__A_op38, TestBlock__B_op82);
  assign smul_75936 = smul32b_32b_x_32b(TestBlock__A_op39, TestBlock__B_op92);
  assign add_75937 = smul_75405 + smul_75406;
  assign add_75938 = smul_75407 + smul_75408;
  assign smul_75939 = smul32b_32b_x_32b(TestBlock__A_op34, TestBlock__B_op43);
  assign smul_75940 = smul32b_32b_x_32b(TestBlock__A_op35, TestBlock__B_op53);
  assign smul_75941 = smul32b_32b_x_32b(TestBlock__A_op36, TestBlock__B_op63);
  assign smul_75942 = smul32b_32b_x_32b(TestBlock__A_op37, TestBlock__B_op73);
  assign smul_75943 = smul32b_32b_x_32b(TestBlock__A_op38, TestBlock__B_op83);
  assign smul_75944 = smul32b_32b_x_32b(TestBlock__A_op39, TestBlock__B_op93);
  assign add_75945 = smul_75409 + smul_75410;
  assign add_75946 = smul_75411 + smul_75412;
  assign smul_75947 = smul32b_32b_x_32b(TestBlock__A_op34, TestBlock__B_op44);
  assign smul_75948 = smul32b_32b_x_32b(TestBlock__A_op35, TestBlock__B_op54);
  assign smul_75949 = smul32b_32b_x_32b(TestBlock__A_op36, TestBlock__B_op64);
  assign smul_75950 = smul32b_32b_x_32b(TestBlock__A_op37, TestBlock__B_op74);
  assign smul_75951 = smul32b_32b_x_32b(TestBlock__A_op38, TestBlock__B_op84);
  assign smul_75952 = smul32b_32b_x_32b(TestBlock__A_op39, TestBlock__B_op94);
  assign add_75953 = smul_75413 + smul_75414;
  assign add_75954 = smul_75415 + smul_75416;
  assign smul_75955 = smul32b_32b_x_32b(TestBlock__A_op34, TestBlock__B_op45);
  assign smul_75956 = smul32b_32b_x_32b(TestBlock__A_op35, TestBlock__B_op55);
  assign smul_75957 = smul32b_32b_x_32b(TestBlock__A_op36, TestBlock__B_op65);
  assign smul_75958 = smul32b_32b_x_32b(TestBlock__A_op37, TestBlock__B_op75);
  assign smul_75959 = smul32b_32b_x_32b(TestBlock__A_op38, TestBlock__B_op85);
  assign smul_75960 = smul32b_32b_x_32b(TestBlock__A_op39, TestBlock__B_op95);
  assign add_75961 = smul_75417 + smul_75418;
  assign add_75962 = smul_75419 + smul_75420;
  assign smul_75963 = smul32b_32b_x_32b(TestBlock__A_op34, TestBlock__B_op46);
  assign smul_75964 = smul32b_32b_x_32b(TestBlock__A_op35, TestBlock__B_op56);
  assign smul_75965 = smul32b_32b_x_32b(TestBlock__A_op36, TestBlock__B_op66);
  assign smul_75966 = smul32b_32b_x_32b(TestBlock__A_op37, TestBlock__B_op76);
  assign smul_75967 = smul32b_32b_x_32b(TestBlock__A_op38, TestBlock__B_op86);
  assign smul_75968 = smul32b_32b_x_32b(TestBlock__A_op39, TestBlock__B_op96);
  assign add_75969 = smul_75421 + smul_75422;
  assign add_75970 = smul_75423 + smul_75424;
  assign smul_75971 = smul32b_32b_x_32b(TestBlock__A_op34, TestBlock__B_op47);
  assign smul_75972 = smul32b_32b_x_32b(TestBlock__A_op35, TestBlock__B_op57);
  assign smul_75973 = smul32b_32b_x_32b(TestBlock__A_op36, TestBlock__B_op67);
  assign smul_75974 = smul32b_32b_x_32b(TestBlock__A_op37, TestBlock__B_op77);
  assign smul_75975 = smul32b_32b_x_32b(TestBlock__A_op38, TestBlock__B_op87);
  assign smul_75976 = smul32b_32b_x_32b(TestBlock__A_op39, TestBlock__B_op97);
  assign add_75977 = smul_75425 + smul_75426;
  assign add_75978 = smul_75427 + smul_75428;
  assign smul_75979 = smul32b_32b_x_32b(TestBlock__A_op34, TestBlock__B_op48);
  assign smul_75980 = smul32b_32b_x_32b(TestBlock__A_op35, TestBlock__B_op58);
  assign smul_75981 = smul32b_32b_x_32b(TestBlock__A_op36, TestBlock__B_op68);
  assign smul_75982 = smul32b_32b_x_32b(TestBlock__A_op37, TestBlock__B_op78);
  assign smul_75983 = smul32b_32b_x_32b(TestBlock__A_op38, TestBlock__B_op88);
  assign smul_75984 = smul32b_32b_x_32b(TestBlock__A_op39, TestBlock__B_op98);
  assign add_75985 = smul_75429 + smul_75430;
  assign add_75986 = smul_75431 + smul_75432;
  assign smul_75987 = smul32b_32b_x_32b(TestBlock__A_op34, TestBlock__B_op49);
  assign smul_75988 = smul32b_32b_x_32b(TestBlock__A_op35, TestBlock__B_op59);
  assign smul_75989 = smul32b_32b_x_32b(TestBlock__A_op36, TestBlock__B_op69);
  assign smul_75990 = smul32b_32b_x_32b(TestBlock__A_op37, TestBlock__B_op79);
  assign smul_75991 = smul32b_32b_x_32b(TestBlock__A_op38, TestBlock__B_op89);
  assign smul_75992 = smul32b_32b_x_32b(TestBlock__A_op39, TestBlock__B_op99);
  assign add_75993 = smul_75433 + smul_75434;
  assign add_75994 = smul_75435 + smul_75436;
  assign smul_75995 = smul32b_32b_x_32b(TestBlock__A_op44, TestBlock__B_op40);
  assign smul_75996 = smul32b_32b_x_32b(TestBlock__A_op45, TestBlock__B_op50);
  assign smul_75997 = smul32b_32b_x_32b(TestBlock__A_op46, TestBlock__B_op60);
  assign smul_75998 = smul32b_32b_x_32b(TestBlock__A_op47, TestBlock__B_op70);
  assign smul_75999 = smul32b_32b_x_32b(TestBlock__A_op48, TestBlock__B_op80);
  assign smul_76000 = smul32b_32b_x_32b(TestBlock__A_op49, TestBlock__B_op90);
  assign add_76001 = smul_75437 + smul_75438;
  assign add_76002 = smul_75439 + smul_75440;
  assign smul_76003 = smul32b_32b_x_32b(TestBlock__A_op44, TestBlock__B_op41);
  assign smul_76004 = smul32b_32b_x_32b(TestBlock__A_op45, TestBlock__B_op51);
  assign smul_76005 = smul32b_32b_x_32b(TestBlock__A_op46, TestBlock__B_op61);
  assign smul_76006 = smul32b_32b_x_32b(TestBlock__A_op47, TestBlock__B_op71);
  assign smul_76007 = smul32b_32b_x_32b(TestBlock__A_op48, TestBlock__B_op81);
  assign smul_76008 = smul32b_32b_x_32b(TestBlock__A_op49, TestBlock__B_op91);
  assign add_76009 = smul_75441 + smul_75442;
  assign add_76010 = smul_75443 + smul_75444;
  assign smul_76011 = smul32b_32b_x_32b(TestBlock__A_op44, TestBlock__B_op42);
  assign smul_76012 = smul32b_32b_x_32b(TestBlock__A_op45, TestBlock__B_op52);
  assign smul_76013 = smul32b_32b_x_32b(TestBlock__A_op46, TestBlock__B_op62);
  assign smul_76014 = smul32b_32b_x_32b(TestBlock__A_op47, TestBlock__B_op72);
  assign smul_76015 = smul32b_32b_x_32b(TestBlock__A_op48, TestBlock__B_op82);
  assign smul_76016 = smul32b_32b_x_32b(TestBlock__A_op49, TestBlock__B_op92);
  assign add_76017 = smul_75445 + smul_75446;
  assign add_76018 = smul_75447 + smul_75448;
  assign smul_76019 = smul32b_32b_x_32b(TestBlock__A_op44, TestBlock__B_op43);
  assign smul_76020 = smul32b_32b_x_32b(TestBlock__A_op45, TestBlock__B_op53);
  assign smul_76021 = smul32b_32b_x_32b(TestBlock__A_op46, TestBlock__B_op63);
  assign smul_76022 = smul32b_32b_x_32b(TestBlock__A_op47, TestBlock__B_op73);
  assign smul_76023 = smul32b_32b_x_32b(TestBlock__A_op48, TestBlock__B_op83);
  assign smul_76024 = smul32b_32b_x_32b(TestBlock__A_op49, TestBlock__B_op93);
  assign add_76025 = smul_75449 + smul_75450;
  assign add_76026 = smul_75451 + smul_75452;
  assign smul_76027 = smul32b_32b_x_32b(TestBlock__A_op44, TestBlock__B_op44);
  assign smul_76028 = smul32b_32b_x_32b(TestBlock__A_op45, TestBlock__B_op54);
  assign smul_76029 = smul32b_32b_x_32b(TestBlock__A_op46, TestBlock__B_op64);
  assign smul_76030 = smul32b_32b_x_32b(TestBlock__A_op47, TestBlock__B_op74);
  assign smul_76031 = smul32b_32b_x_32b(TestBlock__A_op48, TestBlock__B_op84);
  assign smul_76032 = smul32b_32b_x_32b(TestBlock__A_op49, TestBlock__B_op94);
  assign add_76033 = smul_75453 + smul_75454;
  assign add_76034 = smul_75455 + smul_75456;
  assign smul_76035 = smul32b_32b_x_32b(TestBlock__A_op44, TestBlock__B_op45);
  assign smul_76036 = smul32b_32b_x_32b(TestBlock__A_op45, TestBlock__B_op55);
  assign smul_76037 = smul32b_32b_x_32b(TestBlock__A_op46, TestBlock__B_op65);
  assign smul_76038 = smul32b_32b_x_32b(TestBlock__A_op47, TestBlock__B_op75);
  assign smul_76039 = smul32b_32b_x_32b(TestBlock__A_op48, TestBlock__B_op85);
  assign smul_76040 = smul32b_32b_x_32b(TestBlock__A_op49, TestBlock__B_op95);
  assign add_76041 = smul_75457 + smul_75458;
  assign add_76042 = smul_75459 + smul_75460;
  assign smul_76043 = smul32b_32b_x_32b(TestBlock__A_op44, TestBlock__B_op46);
  assign smul_76044 = smul32b_32b_x_32b(TestBlock__A_op45, TestBlock__B_op56);
  assign smul_76045 = smul32b_32b_x_32b(TestBlock__A_op46, TestBlock__B_op66);
  assign smul_76046 = smul32b_32b_x_32b(TestBlock__A_op47, TestBlock__B_op76);
  assign smul_76047 = smul32b_32b_x_32b(TestBlock__A_op48, TestBlock__B_op86);
  assign smul_76048 = smul32b_32b_x_32b(TestBlock__A_op49, TestBlock__B_op96);
  assign add_76049 = smul_75461 + smul_75462;
  assign add_76050 = smul_75463 + smul_75464;
  assign smul_76051 = smul32b_32b_x_32b(TestBlock__A_op44, TestBlock__B_op47);
  assign smul_76052 = smul32b_32b_x_32b(TestBlock__A_op45, TestBlock__B_op57);
  assign smul_76053 = smul32b_32b_x_32b(TestBlock__A_op46, TestBlock__B_op67);
  assign smul_76054 = smul32b_32b_x_32b(TestBlock__A_op47, TestBlock__B_op77);
  assign smul_76055 = smul32b_32b_x_32b(TestBlock__A_op48, TestBlock__B_op87);
  assign smul_76056 = smul32b_32b_x_32b(TestBlock__A_op49, TestBlock__B_op97);
  assign add_76057 = smul_75465 + smul_75466;
  assign add_76058 = smul_75467 + smul_75468;
  assign smul_76059 = smul32b_32b_x_32b(TestBlock__A_op44, TestBlock__B_op48);
  assign smul_76060 = smul32b_32b_x_32b(TestBlock__A_op45, TestBlock__B_op58);
  assign smul_76061 = smul32b_32b_x_32b(TestBlock__A_op46, TestBlock__B_op68);
  assign smul_76062 = smul32b_32b_x_32b(TestBlock__A_op47, TestBlock__B_op78);
  assign smul_76063 = smul32b_32b_x_32b(TestBlock__A_op48, TestBlock__B_op88);
  assign smul_76064 = smul32b_32b_x_32b(TestBlock__A_op49, TestBlock__B_op98);
  assign add_76065 = smul_75469 + smul_75470;
  assign add_76066 = smul_75471 + smul_75472;
  assign smul_76067 = smul32b_32b_x_32b(TestBlock__A_op44, TestBlock__B_op49);
  assign smul_76068 = smul32b_32b_x_32b(TestBlock__A_op45, TestBlock__B_op59);
  assign smul_76069 = smul32b_32b_x_32b(TestBlock__A_op46, TestBlock__B_op69);
  assign smul_76070 = smul32b_32b_x_32b(TestBlock__A_op47, TestBlock__B_op79);
  assign smul_76071 = smul32b_32b_x_32b(TestBlock__A_op48, TestBlock__B_op89);
  assign smul_76072 = smul32b_32b_x_32b(TestBlock__A_op49, TestBlock__B_op99);
  assign add_76073 = smul_75473 + smul_75474;
  assign add_76074 = smul_75475 + smul_75476;
  assign smul_76075 = smul32b_32b_x_32b(TestBlock__A_op54, TestBlock__B_op40);
  assign smul_76076 = smul32b_32b_x_32b(TestBlock__A_op55, TestBlock__B_op50);
  assign smul_76077 = smul32b_32b_x_32b(TestBlock__A_op56, TestBlock__B_op60);
  assign smul_76078 = smul32b_32b_x_32b(TestBlock__A_op57, TestBlock__B_op70);
  assign smul_76079 = smul32b_32b_x_32b(TestBlock__A_op58, TestBlock__B_op80);
  assign smul_76080 = smul32b_32b_x_32b(TestBlock__A_op59, TestBlock__B_op90);
  assign add_76081 = smul_75477 + smul_75478;
  assign add_76082 = smul_75479 + smul_75480;
  assign smul_76083 = smul32b_32b_x_32b(TestBlock__A_op54, TestBlock__B_op41);
  assign smul_76084 = smul32b_32b_x_32b(TestBlock__A_op55, TestBlock__B_op51);
  assign smul_76085 = smul32b_32b_x_32b(TestBlock__A_op56, TestBlock__B_op61);
  assign smul_76086 = smul32b_32b_x_32b(TestBlock__A_op57, TestBlock__B_op71);
  assign smul_76087 = smul32b_32b_x_32b(TestBlock__A_op58, TestBlock__B_op81);
  assign smul_76088 = smul32b_32b_x_32b(TestBlock__A_op59, TestBlock__B_op91);
  assign add_76089 = smul_75481 + smul_75482;
  assign add_76090 = smul_75483 + smul_75484;
  assign smul_76091 = smul32b_32b_x_32b(TestBlock__A_op54, TestBlock__B_op42);
  assign smul_76092 = smul32b_32b_x_32b(TestBlock__A_op55, TestBlock__B_op52);
  assign smul_76093 = smul32b_32b_x_32b(TestBlock__A_op56, TestBlock__B_op62);
  assign smul_76094 = smul32b_32b_x_32b(TestBlock__A_op57, TestBlock__B_op72);
  assign smul_76095 = smul32b_32b_x_32b(TestBlock__A_op58, TestBlock__B_op82);
  assign smul_76096 = smul32b_32b_x_32b(TestBlock__A_op59, TestBlock__B_op92);
  assign add_76097 = smul_75485 + smul_75486;
  assign add_76098 = smul_75487 + smul_75488;
  assign smul_76099 = smul32b_32b_x_32b(TestBlock__A_op54, TestBlock__B_op43);
  assign smul_76100 = smul32b_32b_x_32b(TestBlock__A_op55, TestBlock__B_op53);
  assign smul_76101 = smul32b_32b_x_32b(TestBlock__A_op56, TestBlock__B_op63);
  assign smul_76102 = smul32b_32b_x_32b(TestBlock__A_op57, TestBlock__B_op73);
  assign smul_76103 = smul32b_32b_x_32b(TestBlock__A_op58, TestBlock__B_op83);
  assign smul_76104 = smul32b_32b_x_32b(TestBlock__A_op59, TestBlock__B_op93);
  assign add_76105 = smul_75489 + smul_75490;
  assign add_76106 = smul_75491 + smul_75492;
  assign smul_76107 = smul32b_32b_x_32b(TestBlock__A_op54, TestBlock__B_op44);
  assign smul_76108 = smul32b_32b_x_32b(TestBlock__A_op55, TestBlock__B_op54);
  assign smul_76109 = smul32b_32b_x_32b(TestBlock__A_op56, TestBlock__B_op64);
  assign smul_76110 = smul32b_32b_x_32b(TestBlock__A_op57, TestBlock__B_op74);
  assign smul_76111 = smul32b_32b_x_32b(TestBlock__A_op58, TestBlock__B_op84);
  assign smul_76112 = smul32b_32b_x_32b(TestBlock__A_op59, TestBlock__B_op94);
  assign add_76113 = smul_75493 + smul_75494;
  assign add_76114 = smul_75495 + smul_75496;
  assign smul_76115 = smul32b_32b_x_32b(TestBlock__A_op54, TestBlock__B_op45);
  assign smul_76116 = smul32b_32b_x_32b(TestBlock__A_op55, TestBlock__B_op55);
  assign smul_76117 = smul32b_32b_x_32b(TestBlock__A_op56, TestBlock__B_op65);
  assign smul_76118 = smul32b_32b_x_32b(TestBlock__A_op57, TestBlock__B_op75);
  assign smul_76119 = smul32b_32b_x_32b(TestBlock__A_op58, TestBlock__B_op85);
  assign smul_76120 = smul32b_32b_x_32b(TestBlock__A_op59, TestBlock__B_op95);
  assign add_76121 = smul_75497 + smul_75498;
  assign add_76122 = smul_75499 + smul_75500;
  assign smul_76123 = smul32b_32b_x_32b(TestBlock__A_op54, TestBlock__B_op46);
  assign smul_76124 = smul32b_32b_x_32b(TestBlock__A_op55, TestBlock__B_op56);
  assign smul_76125 = smul32b_32b_x_32b(TestBlock__A_op56, TestBlock__B_op66);
  assign smul_76126 = smul32b_32b_x_32b(TestBlock__A_op57, TestBlock__B_op76);
  assign smul_76127 = smul32b_32b_x_32b(TestBlock__A_op58, TestBlock__B_op86);
  assign smul_76128 = smul32b_32b_x_32b(TestBlock__A_op59, TestBlock__B_op96);
  assign add_76129 = smul_75501 + smul_75502;
  assign add_76130 = smul_75503 + smul_75504;
  assign smul_76131 = smul32b_32b_x_32b(TestBlock__A_op54, TestBlock__B_op47);
  assign smul_76132 = smul32b_32b_x_32b(TestBlock__A_op55, TestBlock__B_op57);
  assign smul_76133 = smul32b_32b_x_32b(TestBlock__A_op56, TestBlock__B_op67);
  assign smul_76134 = smul32b_32b_x_32b(TestBlock__A_op57, TestBlock__B_op77);
  assign smul_76135 = smul32b_32b_x_32b(TestBlock__A_op58, TestBlock__B_op87);
  assign smul_76136 = smul32b_32b_x_32b(TestBlock__A_op59, TestBlock__B_op97);
  assign add_76137 = smul_75505 + smul_75506;
  assign add_76138 = smul_75507 + smul_75508;
  assign smul_76139 = smul32b_32b_x_32b(TestBlock__A_op54, TestBlock__B_op48);
  assign smul_76140 = smul32b_32b_x_32b(TestBlock__A_op55, TestBlock__B_op58);
  assign smul_76141 = smul32b_32b_x_32b(TestBlock__A_op56, TestBlock__B_op68);
  assign smul_76142 = smul32b_32b_x_32b(TestBlock__A_op57, TestBlock__B_op78);
  assign smul_76143 = smul32b_32b_x_32b(TestBlock__A_op58, TestBlock__B_op88);
  assign smul_76144 = smul32b_32b_x_32b(TestBlock__A_op59, TestBlock__B_op98);
  assign add_76145 = smul_75509 + smul_75510;
  assign add_76146 = smul_75511 + smul_75512;
  assign smul_76147 = smul32b_32b_x_32b(TestBlock__A_op54, TestBlock__B_op49);
  assign smul_76148 = smul32b_32b_x_32b(TestBlock__A_op55, TestBlock__B_op59);
  assign smul_76149 = smul32b_32b_x_32b(TestBlock__A_op56, TestBlock__B_op69);
  assign smul_76150 = smul32b_32b_x_32b(TestBlock__A_op57, TestBlock__B_op79);
  assign smul_76151 = smul32b_32b_x_32b(TestBlock__A_op58, TestBlock__B_op89);
  assign smul_76152 = smul32b_32b_x_32b(TestBlock__A_op59, TestBlock__B_op99);
  assign add_76153 = smul_75513 + smul_75514;
  assign add_76154 = smul_75515 + smul_75516;
  assign smul_76155 = smul32b_32b_x_32b(TestBlock__A_op64, TestBlock__B_op40);
  assign smul_76156 = smul32b_32b_x_32b(TestBlock__A_op65, TestBlock__B_op50);
  assign smul_76157 = smul32b_32b_x_32b(TestBlock__A_op66, TestBlock__B_op60);
  assign smul_76158 = smul32b_32b_x_32b(TestBlock__A_op67, TestBlock__B_op70);
  assign smul_76159 = smul32b_32b_x_32b(TestBlock__A_op68, TestBlock__B_op80);
  assign smul_76160 = smul32b_32b_x_32b(TestBlock__A_op69, TestBlock__B_op90);
  assign add_76161 = smul_75517 + smul_75518;
  assign add_76162 = smul_75519 + smul_75520;
  assign smul_76163 = smul32b_32b_x_32b(TestBlock__A_op64, TestBlock__B_op41);
  assign smul_76164 = smul32b_32b_x_32b(TestBlock__A_op65, TestBlock__B_op51);
  assign smul_76165 = smul32b_32b_x_32b(TestBlock__A_op66, TestBlock__B_op61);
  assign smul_76166 = smul32b_32b_x_32b(TestBlock__A_op67, TestBlock__B_op71);
  assign smul_76167 = smul32b_32b_x_32b(TestBlock__A_op68, TestBlock__B_op81);
  assign smul_76168 = smul32b_32b_x_32b(TestBlock__A_op69, TestBlock__B_op91);
  assign add_76169 = smul_75521 + smul_75522;
  assign add_76170 = smul_75523 + smul_75524;
  assign smul_76171 = smul32b_32b_x_32b(TestBlock__A_op64, TestBlock__B_op42);
  assign smul_76172 = smul32b_32b_x_32b(TestBlock__A_op65, TestBlock__B_op52);
  assign smul_76173 = smul32b_32b_x_32b(TestBlock__A_op66, TestBlock__B_op62);
  assign smul_76174 = smul32b_32b_x_32b(TestBlock__A_op67, TestBlock__B_op72);
  assign smul_76175 = smul32b_32b_x_32b(TestBlock__A_op68, TestBlock__B_op82);
  assign smul_76176 = smul32b_32b_x_32b(TestBlock__A_op69, TestBlock__B_op92);
  assign add_76177 = smul_75525 + smul_75526;
  assign add_76178 = smul_75527 + smul_75528;
  assign smul_76179 = smul32b_32b_x_32b(TestBlock__A_op64, TestBlock__B_op43);
  assign smul_76180 = smul32b_32b_x_32b(TestBlock__A_op65, TestBlock__B_op53);
  assign smul_76181 = smul32b_32b_x_32b(TestBlock__A_op66, TestBlock__B_op63);
  assign smul_76182 = smul32b_32b_x_32b(TestBlock__A_op67, TestBlock__B_op73);
  assign smul_76183 = smul32b_32b_x_32b(TestBlock__A_op68, TestBlock__B_op83);
  assign smul_76184 = smul32b_32b_x_32b(TestBlock__A_op69, TestBlock__B_op93);
  assign add_76185 = smul_75529 + smul_75530;
  assign add_76186 = smul_75531 + smul_75532;
  assign smul_76187 = smul32b_32b_x_32b(TestBlock__A_op64, TestBlock__B_op44);
  assign smul_76188 = smul32b_32b_x_32b(TestBlock__A_op65, TestBlock__B_op54);
  assign smul_76189 = smul32b_32b_x_32b(TestBlock__A_op66, TestBlock__B_op64);
  assign smul_76190 = smul32b_32b_x_32b(TestBlock__A_op67, TestBlock__B_op74);
  assign smul_76191 = smul32b_32b_x_32b(TestBlock__A_op68, TestBlock__B_op84);
  assign smul_76192 = smul32b_32b_x_32b(TestBlock__A_op69, TestBlock__B_op94);
  assign add_76193 = smul_75533 + smul_75534;
  assign add_76194 = smul_75535 + smul_75536;
  assign smul_76195 = smul32b_32b_x_32b(TestBlock__A_op64, TestBlock__B_op45);
  assign smul_76196 = smul32b_32b_x_32b(TestBlock__A_op65, TestBlock__B_op55);
  assign smul_76197 = smul32b_32b_x_32b(TestBlock__A_op66, TestBlock__B_op65);
  assign smul_76198 = smul32b_32b_x_32b(TestBlock__A_op67, TestBlock__B_op75);
  assign smul_76199 = smul32b_32b_x_32b(TestBlock__A_op68, TestBlock__B_op85);
  assign smul_76200 = smul32b_32b_x_32b(TestBlock__A_op69, TestBlock__B_op95);
  assign add_76201 = smul_75537 + smul_75538;
  assign add_76202 = smul_75539 + smul_75540;
  assign smul_76203 = smul32b_32b_x_32b(TestBlock__A_op64, TestBlock__B_op46);
  assign smul_76204 = smul32b_32b_x_32b(TestBlock__A_op65, TestBlock__B_op56);
  assign smul_76205 = smul32b_32b_x_32b(TestBlock__A_op66, TestBlock__B_op66);
  assign smul_76206 = smul32b_32b_x_32b(TestBlock__A_op67, TestBlock__B_op76);
  assign smul_76207 = smul32b_32b_x_32b(TestBlock__A_op68, TestBlock__B_op86);
  assign smul_76208 = smul32b_32b_x_32b(TestBlock__A_op69, TestBlock__B_op96);
  assign add_76209 = smul_75541 + smul_75542;
  assign add_76210 = smul_75543 + smul_75544;
  assign smul_76211 = smul32b_32b_x_32b(TestBlock__A_op64, TestBlock__B_op47);
  assign smul_76212 = smul32b_32b_x_32b(TestBlock__A_op65, TestBlock__B_op57);
  assign smul_76213 = smul32b_32b_x_32b(TestBlock__A_op66, TestBlock__B_op67);
  assign smul_76214 = smul32b_32b_x_32b(TestBlock__A_op67, TestBlock__B_op77);
  assign smul_76215 = smul32b_32b_x_32b(TestBlock__A_op68, TestBlock__B_op87);
  assign smul_76216 = smul32b_32b_x_32b(TestBlock__A_op69, TestBlock__B_op97);
  assign add_76217 = smul_75545 + smul_75546;
  assign add_76218 = smul_75547 + smul_75548;
  assign smul_76219 = smul32b_32b_x_32b(TestBlock__A_op64, TestBlock__B_op48);
  assign smul_76220 = smul32b_32b_x_32b(TestBlock__A_op65, TestBlock__B_op58);
  assign smul_76221 = smul32b_32b_x_32b(TestBlock__A_op66, TestBlock__B_op68);
  assign smul_76222 = smul32b_32b_x_32b(TestBlock__A_op67, TestBlock__B_op78);
  assign smul_76223 = smul32b_32b_x_32b(TestBlock__A_op68, TestBlock__B_op88);
  assign smul_76224 = smul32b_32b_x_32b(TestBlock__A_op69, TestBlock__B_op98);
  assign add_76225 = smul_75549 + smul_75550;
  assign add_76226 = smul_75551 + smul_75552;
  assign smul_76227 = smul32b_32b_x_32b(TestBlock__A_op64, TestBlock__B_op49);
  assign smul_76228 = smul32b_32b_x_32b(TestBlock__A_op65, TestBlock__B_op59);
  assign smul_76229 = smul32b_32b_x_32b(TestBlock__A_op66, TestBlock__B_op69);
  assign smul_76230 = smul32b_32b_x_32b(TestBlock__A_op67, TestBlock__B_op79);
  assign smul_76231 = smul32b_32b_x_32b(TestBlock__A_op68, TestBlock__B_op89);
  assign smul_76232 = smul32b_32b_x_32b(TestBlock__A_op69, TestBlock__B_op99);
  assign add_76233 = smul_75553 + smul_75554;
  assign add_76234 = smul_75555 + smul_75556;
  assign smul_76235 = smul32b_32b_x_32b(TestBlock__A_op74, TestBlock__B_op40);
  assign smul_76236 = smul32b_32b_x_32b(TestBlock__A_op75, TestBlock__B_op50);
  assign smul_76237 = smul32b_32b_x_32b(TestBlock__A_op76, TestBlock__B_op60);
  assign smul_76238 = smul32b_32b_x_32b(TestBlock__A_op77, TestBlock__B_op70);
  assign smul_76239 = smul32b_32b_x_32b(TestBlock__A_op78, TestBlock__B_op80);
  assign smul_76240 = smul32b_32b_x_32b(TestBlock__A_op79, TestBlock__B_op90);
  assign add_76241 = smul_75557 + smul_75558;
  assign add_76242 = smul_75559 + smul_75560;
  assign smul_76243 = smul32b_32b_x_32b(TestBlock__A_op74, TestBlock__B_op41);
  assign smul_76244 = smul32b_32b_x_32b(TestBlock__A_op75, TestBlock__B_op51);
  assign smul_76245 = smul32b_32b_x_32b(TestBlock__A_op76, TestBlock__B_op61);
  assign smul_76246 = smul32b_32b_x_32b(TestBlock__A_op77, TestBlock__B_op71);
  assign smul_76247 = smul32b_32b_x_32b(TestBlock__A_op78, TestBlock__B_op81);
  assign smul_76248 = smul32b_32b_x_32b(TestBlock__A_op79, TestBlock__B_op91);
  assign add_76249 = smul_75561 + smul_75562;
  assign add_76250 = smul_75563 + smul_75564;
  assign smul_76251 = smul32b_32b_x_32b(TestBlock__A_op74, TestBlock__B_op42);
  assign smul_76252 = smul32b_32b_x_32b(TestBlock__A_op75, TestBlock__B_op52);
  assign smul_76253 = smul32b_32b_x_32b(TestBlock__A_op76, TestBlock__B_op62);
  assign smul_76254 = smul32b_32b_x_32b(TestBlock__A_op77, TestBlock__B_op72);
  assign smul_76255 = smul32b_32b_x_32b(TestBlock__A_op78, TestBlock__B_op82);
  assign smul_76256 = smul32b_32b_x_32b(TestBlock__A_op79, TestBlock__B_op92);
  assign add_76257 = smul_75565 + smul_75566;
  assign add_76258 = smul_75567 + smul_75568;
  assign smul_76259 = smul32b_32b_x_32b(TestBlock__A_op74, TestBlock__B_op43);
  assign smul_76260 = smul32b_32b_x_32b(TestBlock__A_op75, TestBlock__B_op53);
  assign smul_76261 = smul32b_32b_x_32b(TestBlock__A_op76, TestBlock__B_op63);
  assign smul_76262 = smul32b_32b_x_32b(TestBlock__A_op77, TestBlock__B_op73);
  assign smul_76263 = smul32b_32b_x_32b(TestBlock__A_op78, TestBlock__B_op83);
  assign smul_76264 = smul32b_32b_x_32b(TestBlock__A_op79, TestBlock__B_op93);
  assign add_76265 = smul_75569 + smul_75570;
  assign add_76266 = smul_75571 + smul_75572;
  assign smul_76267 = smul32b_32b_x_32b(TestBlock__A_op74, TestBlock__B_op44);
  assign smul_76268 = smul32b_32b_x_32b(TestBlock__A_op75, TestBlock__B_op54);
  assign smul_76269 = smul32b_32b_x_32b(TestBlock__A_op76, TestBlock__B_op64);
  assign smul_76270 = smul32b_32b_x_32b(TestBlock__A_op77, TestBlock__B_op74);
  assign smul_76271 = smul32b_32b_x_32b(TestBlock__A_op78, TestBlock__B_op84);
  assign smul_76272 = smul32b_32b_x_32b(TestBlock__A_op79, TestBlock__B_op94);
  assign add_76273 = smul_75573 + smul_75574;
  assign add_76274 = smul_75575 + smul_75576;
  assign smul_76275 = smul32b_32b_x_32b(TestBlock__A_op74, TestBlock__B_op45);
  assign smul_76276 = smul32b_32b_x_32b(TestBlock__A_op75, TestBlock__B_op55);
  assign smul_76277 = smul32b_32b_x_32b(TestBlock__A_op76, TestBlock__B_op65);
  assign smul_76278 = smul32b_32b_x_32b(TestBlock__A_op77, TestBlock__B_op75);
  assign smul_76279 = smul32b_32b_x_32b(TestBlock__A_op78, TestBlock__B_op85);
  assign smul_76280 = smul32b_32b_x_32b(TestBlock__A_op79, TestBlock__B_op95);
  assign add_76281 = smul_75577 + smul_75578;
  assign add_76282 = smul_75579 + smul_75580;
  assign smul_76283 = smul32b_32b_x_32b(TestBlock__A_op74, TestBlock__B_op46);
  assign smul_76284 = smul32b_32b_x_32b(TestBlock__A_op75, TestBlock__B_op56);
  assign smul_76285 = smul32b_32b_x_32b(TestBlock__A_op76, TestBlock__B_op66);
  assign smul_76286 = smul32b_32b_x_32b(TestBlock__A_op77, TestBlock__B_op76);
  assign smul_76287 = smul32b_32b_x_32b(TestBlock__A_op78, TestBlock__B_op86);
  assign smul_76288 = smul32b_32b_x_32b(TestBlock__A_op79, TestBlock__B_op96);
  assign add_76289 = smul_75581 + smul_75582;
  assign add_76290 = smul_75583 + smul_75584;
  assign smul_76291 = smul32b_32b_x_32b(TestBlock__A_op74, TestBlock__B_op47);
  assign smul_76292 = smul32b_32b_x_32b(TestBlock__A_op75, TestBlock__B_op57);
  assign smul_76293 = smul32b_32b_x_32b(TestBlock__A_op76, TestBlock__B_op67);
  assign smul_76294 = smul32b_32b_x_32b(TestBlock__A_op77, TestBlock__B_op77);
  assign smul_76295 = smul32b_32b_x_32b(TestBlock__A_op78, TestBlock__B_op87);
  assign smul_76296 = smul32b_32b_x_32b(TestBlock__A_op79, TestBlock__B_op97);
  assign add_76297 = smul_75585 + smul_75586;
  assign add_76298 = smul_75587 + smul_75588;
  assign smul_76299 = smul32b_32b_x_32b(TestBlock__A_op74, TestBlock__B_op48);
  assign smul_76300 = smul32b_32b_x_32b(TestBlock__A_op75, TestBlock__B_op58);
  assign smul_76301 = smul32b_32b_x_32b(TestBlock__A_op76, TestBlock__B_op68);
  assign smul_76302 = smul32b_32b_x_32b(TestBlock__A_op77, TestBlock__B_op78);
  assign smul_76303 = smul32b_32b_x_32b(TestBlock__A_op78, TestBlock__B_op88);
  assign smul_76304 = smul32b_32b_x_32b(TestBlock__A_op79, TestBlock__B_op98);
  assign add_76305 = smul_75589 + smul_75590;
  assign add_76306 = smul_75591 + smul_75592;
  assign smul_76307 = smul32b_32b_x_32b(TestBlock__A_op74, TestBlock__B_op49);
  assign smul_76308 = smul32b_32b_x_32b(TestBlock__A_op75, TestBlock__B_op59);
  assign smul_76309 = smul32b_32b_x_32b(TestBlock__A_op76, TestBlock__B_op69);
  assign smul_76310 = smul32b_32b_x_32b(TestBlock__A_op77, TestBlock__B_op79);
  assign smul_76311 = smul32b_32b_x_32b(TestBlock__A_op78, TestBlock__B_op89);
  assign smul_76312 = smul32b_32b_x_32b(TestBlock__A_op79, TestBlock__B_op99);
  assign add_76313 = smul_75593 + smul_75594;
  assign add_76314 = smul_75595 + smul_75596;
  assign smul_76315 = smul32b_32b_x_32b(TestBlock__A_op84, TestBlock__B_op40);
  assign smul_76316 = smul32b_32b_x_32b(TestBlock__A_op85, TestBlock__B_op50);
  assign smul_76317 = smul32b_32b_x_32b(TestBlock__A_op86, TestBlock__B_op60);
  assign smul_76318 = smul32b_32b_x_32b(TestBlock__A_op87, TestBlock__B_op70);
  assign smul_76319 = smul32b_32b_x_32b(TestBlock__A_op88, TestBlock__B_op80);
  assign smul_76320 = smul32b_32b_x_32b(TestBlock__A_op89, TestBlock__B_op90);
  assign add_76321 = smul_75597 + smul_75598;
  assign add_76322 = smul_75599 + smul_75600;
  assign smul_76323 = smul32b_32b_x_32b(TestBlock__A_op84, TestBlock__B_op41);
  assign smul_76324 = smul32b_32b_x_32b(TestBlock__A_op85, TestBlock__B_op51);
  assign smul_76325 = smul32b_32b_x_32b(TestBlock__A_op86, TestBlock__B_op61);
  assign smul_76326 = smul32b_32b_x_32b(TestBlock__A_op87, TestBlock__B_op71);
  assign smul_76327 = smul32b_32b_x_32b(TestBlock__A_op88, TestBlock__B_op81);
  assign smul_76328 = smul32b_32b_x_32b(TestBlock__A_op89, TestBlock__B_op91);
  assign add_76329 = smul_75601 + smul_75602;
  assign add_76330 = smul_75603 + smul_75604;
  assign smul_76331 = smul32b_32b_x_32b(TestBlock__A_op84, TestBlock__B_op42);
  assign smul_76332 = smul32b_32b_x_32b(TestBlock__A_op85, TestBlock__B_op52);
  assign smul_76333 = smul32b_32b_x_32b(TestBlock__A_op86, TestBlock__B_op62);
  assign smul_76334 = smul32b_32b_x_32b(TestBlock__A_op87, TestBlock__B_op72);
  assign smul_76335 = smul32b_32b_x_32b(TestBlock__A_op88, TestBlock__B_op82);
  assign smul_76336 = smul32b_32b_x_32b(TestBlock__A_op89, TestBlock__B_op92);
  assign add_76337 = smul_75605 + smul_75606;
  assign add_76338 = smul_75607 + smul_75608;
  assign smul_76339 = smul32b_32b_x_32b(TestBlock__A_op84, TestBlock__B_op43);
  assign smul_76340 = smul32b_32b_x_32b(TestBlock__A_op85, TestBlock__B_op53);
  assign smul_76341 = smul32b_32b_x_32b(TestBlock__A_op86, TestBlock__B_op63);
  assign smul_76342 = smul32b_32b_x_32b(TestBlock__A_op87, TestBlock__B_op73);
  assign smul_76343 = smul32b_32b_x_32b(TestBlock__A_op88, TestBlock__B_op83);
  assign smul_76344 = smul32b_32b_x_32b(TestBlock__A_op89, TestBlock__B_op93);
  assign add_76345 = smul_75609 + smul_75610;
  assign add_76346 = smul_75611 + smul_75612;
  assign smul_76347 = smul32b_32b_x_32b(TestBlock__A_op84, TestBlock__B_op44);
  assign smul_76348 = smul32b_32b_x_32b(TestBlock__A_op85, TestBlock__B_op54);
  assign smul_76349 = smul32b_32b_x_32b(TestBlock__A_op86, TestBlock__B_op64);
  assign smul_76350 = smul32b_32b_x_32b(TestBlock__A_op87, TestBlock__B_op74);
  assign smul_76351 = smul32b_32b_x_32b(TestBlock__A_op88, TestBlock__B_op84);
  assign smul_76352 = smul32b_32b_x_32b(TestBlock__A_op89, TestBlock__B_op94);
  assign add_76353 = smul_75613 + smul_75614;
  assign add_76354 = smul_75615 + smul_75616;
  assign smul_76355 = smul32b_32b_x_32b(TestBlock__A_op84, TestBlock__B_op45);
  assign smul_76356 = smul32b_32b_x_32b(TestBlock__A_op85, TestBlock__B_op55);
  assign smul_76357 = smul32b_32b_x_32b(TestBlock__A_op86, TestBlock__B_op65);
  assign smul_76358 = smul32b_32b_x_32b(TestBlock__A_op87, TestBlock__B_op75);
  assign smul_76359 = smul32b_32b_x_32b(TestBlock__A_op88, TestBlock__B_op85);
  assign smul_76360 = smul32b_32b_x_32b(TestBlock__A_op89, TestBlock__B_op95);
  assign add_76361 = smul_75617 + smul_75618;
  assign add_76362 = smul_75619 + smul_75620;
  assign smul_76363 = smul32b_32b_x_32b(TestBlock__A_op84, TestBlock__B_op46);
  assign smul_76364 = smul32b_32b_x_32b(TestBlock__A_op85, TestBlock__B_op56);
  assign smul_76365 = smul32b_32b_x_32b(TestBlock__A_op86, TestBlock__B_op66);
  assign smul_76366 = smul32b_32b_x_32b(TestBlock__A_op87, TestBlock__B_op76);
  assign smul_76367 = smul32b_32b_x_32b(TestBlock__A_op88, TestBlock__B_op86);
  assign smul_76368 = smul32b_32b_x_32b(TestBlock__A_op89, TestBlock__B_op96);
  assign add_76369 = smul_75621 + smul_75622;
  assign add_76370 = smul_75623 + smul_75624;
  assign smul_76371 = smul32b_32b_x_32b(TestBlock__A_op84, TestBlock__B_op47);
  assign smul_76372 = smul32b_32b_x_32b(TestBlock__A_op85, TestBlock__B_op57);
  assign smul_76373 = smul32b_32b_x_32b(TestBlock__A_op86, TestBlock__B_op67);
  assign smul_76374 = smul32b_32b_x_32b(TestBlock__A_op87, TestBlock__B_op77);
  assign smul_76375 = smul32b_32b_x_32b(TestBlock__A_op88, TestBlock__B_op87);
  assign smul_76376 = smul32b_32b_x_32b(TestBlock__A_op89, TestBlock__B_op97);
  assign add_76377 = smul_75625 + smul_75626;
  assign add_76378 = smul_75627 + smul_75628;
  assign smul_76379 = smul32b_32b_x_32b(TestBlock__A_op84, TestBlock__B_op48);
  assign smul_76380 = smul32b_32b_x_32b(TestBlock__A_op85, TestBlock__B_op58);
  assign smul_76381 = smul32b_32b_x_32b(TestBlock__A_op86, TestBlock__B_op68);
  assign smul_76382 = smul32b_32b_x_32b(TestBlock__A_op87, TestBlock__B_op78);
  assign smul_76383 = smul32b_32b_x_32b(TestBlock__A_op88, TestBlock__B_op88);
  assign smul_76384 = smul32b_32b_x_32b(TestBlock__A_op89, TestBlock__B_op98);
  assign add_76385 = smul_75629 + smul_75630;
  assign add_76386 = smul_75631 + smul_75632;
  assign smul_76387 = smul32b_32b_x_32b(TestBlock__A_op84, TestBlock__B_op49);
  assign smul_76388 = smul32b_32b_x_32b(TestBlock__A_op85, TestBlock__B_op59);
  assign smul_76389 = smul32b_32b_x_32b(TestBlock__A_op86, TestBlock__B_op69);
  assign smul_76390 = smul32b_32b_x_32b(TestBlock__A_op87, TestBlock__B_op79);
  assign smul_76391 = smul32b_32b_x_32b(TestBlock__A_op88, TestBlock__B_op89);
  assign smul_76392 = smul32b_32b_x_32b(TestBlock__A_op89, TestBlock__B_op99);
  assign add_76393 = smul_75633 + smul_75634;
  assign add_76394 = smul_75635 + smul_75636;
  assign smul_76395 = smul32b_32b_x_32b(TestBlock__A_op94, TestBlock__B_op40);
  assign smul_76396 = smul32b_32b_x_32b(TestBlock__A_op95, TestBlock__B_op50);
  assign smul_76397 = smul32b_32b_x_32b(TestBlock__A_op96, TestBlock__B_op60);
  assign smul_76398 = smul32b_32b_x_32b(TestBlock__A_op97, TestBlock__B_op70);
  assign smul_76399 = smul32b_32b_x_32b(TestBlock__A_op98, TestBlock__B_op80);
  assign smul_76400 = smul32b_32b_x_32b(TestBlock__A_op99, TestBlock__B_op90);
  assign add_76401 = smul_75637 + smul_75638;
  assign add_76402 = smul_75639 + smul_75640;
  assign smul_76403 = smul32b_32b_x_32b(TestBlock__A_op94, TestBlock__B_op41);
  assign smul_76404 = smul32b_32b_x_32b(TestBlock__A_op95, TestBlock__B_op51);
  assign smul_76405 = smul32b_32b_x_32b(TestBlock__A_op96, TestBlock__B_op61);
  assign smul_76406 = smul32b_32b_x_32b(TestBlock__A_op97, TestBlock__B_op71);
  assign smul_76407 = smul32b_32b_x_32b(TestBlock__A_op98, TestBlock__B_op81);
  assign smul_76408 = smul32b_32b_x_32b(TestBlock__A_op99, TestBlock__B_op91);
  assign add_76409 = smul_75641 + smul_75642;
  assign add_76410 = smul_75643 + smul_75644;
  assign smul_76411 = smul32b_32b_x_32b(TestBlock__A_op94, TestBlock__B_op42);
  assign smul_76412 = smul32b_32b_x_32b(TestBlock__A_op95, TestBlock__B_op52);
  assign smul_76413 = smul32b_32b_x_32b(TestBlock__A_op96, TestBlock__B_op62);
  assign smul_76414 = smul32b_32b_x_32b(TestBlock__A_op97, TestBlock__B_op72);
  assign smul_76415 = smul32b_32b_x_32b(TestBlock__A_op98, TestBlock__B_op82);
  assign smul_76416 = smul32b_32b_x_32b(TestBlock__A_op99, TestBlock__B_op92);
  assign add_76417 = smul_75645 + smul_75646;
  assign add_76418 = smul_75647 + smul_75648;
  assign smul_76419 = smul32b_32b_x_32b(TestBlock__A_op94, TestBlock__B_op43);
  assign smul_76420 = smul32b_32b_x_32b(TestBlock__A_op95, TestBlock__B_op53);
  assign smul_76421 = smul32b_32b_x_32b(TestBlock__A_op96, TestBlock__B_op63);
  assign smul_76422 = smul32b_32b_x_32b(TestBlock__A_op97, TestBlock__B_op73);
  assign smul_76423 = smul32b_32b_x_32b(TestBlock__A_op98, TestBlock__B_op83);
  assign smul_76424 = smul32b_32b_x_32b(TestBlock__A_op99, TestBlock__B_op93);
  assign add_76425 = smul_75649 + smul_75650;
  assign add_76426 = smul_75651 + smul_75652;
  assign smul_76427 = smul32b_32b_x_32b(TestBlock__A_op94, TestBlock__B_op44);
  assign smul_76428 = smul32b_32b_x_32b(TestBlock__A_op95, TestBlock__B_op54);
  assign smul_76429 = smul32b_32b_x_32b(TestBlock__A_op96, TestBlock__B_op64);
  assign smul_76430 = smul32b_32b_x_32b(TestBlock__A_op97, TestBlock__B_op74);
  assign smul_76431 = smul32b_32b_x_32b(TestBlock__A_op98, TestBlock__B_op84);
  assign smul_76432 = smul32b_32b_x_32b(TestBlock__A_op99, TestBlock__B_op94);
  assign add_76433 = smul_75653 + smul_75654;
  assign add_76434 = smul_75655 + smul_75656;
  assign smul_76435 = smul32b_32b_x_32b(TestBlock__A_op94, TestBlock__B_op45);
  assign smul_76436 = smul32b_32b_x_32b(TestBlock__A_op95, TestBlock__B_op55);
  assign smul_76437 = smul32b_32b_x_32b(TestBlock__A_op96, TestBlock__B_op65);
  assign smul_76438 = smul32b_32b_x_32b(TestBlock__A_op97, TestBlock__B_op75);
  assign smul_76439 = smul32b_32b_x_32b(TestBlock__A_op98, TestBlock__B_op85);
  assign smul_76440 = smul32b_32b_x_32b(TestBlock__A_op99, TestBlock__B_op95);
  assign add_76441 = smul_75657 + smul_75658;
  assign add_76442 = smul_75659 + smul_75660;
  assign smul_76443 = smul32b_32b_x_32b(TestBlock__A_op94, TestBlock__B_op46);
  assign smul_76444 = smul32b_32b_x_32b(TestBlock__A_op95, TestBlock__B_op56);
  assign smul_76445 = smul32b_32b_x_32b(TestBlock__A_op96, TestBlock__B_op66);
  assign smul_76446 = smul32b_32b_x_32b(TestBlock__A_op97, TestBlock__B_op76);
  assign smul_76447 = smul32b_32b_x_32b(TestBlock__A_op98, TestBlock__B_op86);
  assign smul_76448 = smul32b_32b_x_32b(TestBlock__A_op99, TestBlock__B_op96);
  assign add_76449 = smul_75661 + smul_75662;
  assign add_76450 = smul_75663 + smul_75664;
  assign smul_76451 = smul32b_32b_x_32b(TestBlock__A_op94, TestBlock__B_op47);
  assign smul_76452 = smul32b_32b_x_32b(TestBlock__A_op95, TestBlock__B_op57);
  assign smul_76453 = smul32b_32b_x_32b(TestBlock__A_op96, TestBlock__B_op67);
  assign smul_76454 = smul32b_32b_x_32b(TestBlock__A_op97, TestBlock__B_op77);
  assign smul_76455 = smul32b_32b_x_32b(TestBlock__A_op98, TestBlock__B_op87);
  assign smul_76456 = smul32b_32b_x_32b(TestBlock__A_op99, TestBlock__B_op97);
  assign add_76457 = smul_75665 + smul_75666;
  assign add_76458 = smul_75667 + smul_75668;
  assign smul_76459 = smul32b_32b_x_32b(TestBlock__A_op94, TestBlock__B_op48);
  assign smul_76460 = smul32b_32b_x_32b(TestBlock__A_op95, TestBlock__B_op58);
  assign smul_76461 = smul32b_32b_x_32b(TestBlock__A_op96, TestBlock__B_op68);
  assign smul_76462 = smul32b_32b_x_32b(TestBlock__A_op97, TestBlock__B_op78);
  assign smul_76463 = smul32b_32b_x_32b(TestBlock__A_op98, TestBlock__B_op88);
  assign smul_76464 = smul32b_32b_x_32b(TestBlock__A_op99, TestBlock__B_op98);
  assign add_76465 = smul_75669 + smul_75670;
  assign add_76466 = smul_75671 + smul_75672;
  assign smul_76467 = smul32b_32b_x_32b(TestBlock__A_op94, TestBlock__B_op49);
  assign smul_76468 = smul32b_32b_x_32b(TestBlock__A_op95, TestBlock__B_op59);
  assign smul_76469 = smul32b_32b_x_32b(TestBlock__A_op96, TestBlock__B_op69);
  assign smul_76470 = smul32b_32b_x_32b(TestBlock__A_op97, TestBlock__B_op79);
  assign smul_76471 = smul32b_32b_x_32b(TestBlock__A_op98, TestBlock__B_op89);
  assign smul_76472 = smul32b_32b_x_32b(TestBlock__A_op99, TestBlock__B_op99);
  assign add_76473 = add_75673 + add_75674;
  assign add_76474 = smul_75675 + smul_75676;
  assign add_76475 = smul_75677 + smul_75678;
  assign add_76476 = smul_75679 + smul_75680;
  assign add_76477 = add_75681 + add_75682;
  assign add_76478 = smul_75683 + smul_75684;
  assign add_76479 = smul_75685 + smul_75686;
  assign add_76480 = smul_75687 + smul_75688;
  assign add_76481 = add_75689 + add_75690;
  assign add_76482 = smul_75691 + smul_75692;
  assign add_76483 = smul_75693 + smul_75694;
  assign add_76484 = smul_75695 + smul_75696;
  assign add_76485 = add_75697 + add_75698;
  assign add_76486 = smul_75699 + smul_75700;
  assign add_76487 = smul_75701 + smul_75702;
  assign add_76488 = smul_75703 + smul_75704;
  assign add_76489 = add_75705 + add_75706;
  assign add_76490 = smul_75707 + smul_75708;
  assign add_76491 = smul_75709 + smul_75710;
  assign add_76492 = smul_75711 + smul_75712;
  assign add_76493 = add_75713 + add_75714;
  assign add_76494 = smul_75715 + smul_75716;
  assign add_76495 = smul_75717 + smul_75718;
  assign add_76496 = smul_75719 + smul_75720;
  assign add_76497 = add_75721 + add_75722;
  assign add_76498 = smul_75723 + smul_75724;
  assign add_76499 = smul_75725 + smul_75726;
  assign add_76500 = smul_75727 + smul_75728;
  assign add_76501 = add_75729 + add_75730;
  assign add_76502 = smul_75731 + smul_75732;
  assign add_76503 = smul_75733 + smul_75734;
  assign add_76504 = smul_75735 + smul_75736;
  assign add_76505 = add_75737 + add_75738;
  assign add_76506 = smul_75739 + smul_75740;
  assign add_76507 = smul_75741 + smul_75742;
  assign add_76508 = smul_75743 + smul_75744;
  assign add_76509 = add_75745 + add_75746;
  assign add_76510 = smul_75747 + smul_75748;
  assign add_76511 = smul_75749 + smul_75750;
  assign add_76512 = smul_75751 + smul_75752;
  assign add_76513 = add_75753 + add_75754;
  assign add_76514 = smul_75755 + smul_75756;
  assign add_76515 = smul_75757 + smul_75758;
  assign add_76516 = smul_75759 + smul_75760;
  assign add_76517 = add_75761 + add_75762;
  assign add_76518 = smul_75763 + smul_75764;
  assign add_76519 = smul_75765 + smul_75766;
  assign add_76520 = smul_75767 + smul_75768;
  assign add_76521 = add_75769 + add_75770;
  assign add_76522 = smul_75771 + smul_75772;
  assign add_76523 = smul_75773 + smul_75774;
  assign add_76524 = smul_75775 + smul_75776;
  assign add_76525 = add_75777 + add_75778;
  assign add_76526 = smul_75779 + smul_75780;
  assign add_76527 = smul_75781 + smul_75782;
  assign add_76528 = smul_75783 + smul_75784;
  assign add_76529 = add_75785 + add_75786;
  assign add_76530 = smul_75787 + smul_75788;
  assign add_76531 = smul_75789 + smul_75790;
  assign add_76532 = smul_75791 + smul_75792;
  assign add_76533 = add_75793 + add_75794;
  assign add_76534 = smul_75795 + smul_75796;
  assign add_76535 = smul_75797 + smul_75798;
  assign add_76536 = smul_75799 + smul_75800;
  assign add_76537 = add_75801 + add_75802;
  assign add_76538 = smul_75803 + smul_75804;
  assign add_76539 = smul_75805 + smul_75806;
  assign add_76540 = smul_75807 + smul_75808;
  assign add_76541 = add_75809 + add_75810;
  assign add_76542 = smul_75811 + smul_75812;
  assign add_76543 = smul_75813 + smul_75814;
  assign add_76544 = smul_75815 + smul_75816;
  assign add_76545 = add_75817 + add_75818;
  assign add_76546 = smul_75819 + smul_75820;
  assign add_76547 = smul_75821 + smul_75822;
  assign add_76548 = smul_75823 + smul_75824;
  assign add_76549 = add_75825 + add_75826;
  assign add_76550 = smul_75827 + smul_75828;
  assign add_76551 = smul_75829 + smul_75830;
  assign add_76552 = smul_75831 + smul_75832;
  assign add_76553 = add_75833 + add_75834;
  assign add_76554 = smul_75835 + smul_75836;
  assign add_76555 = smul_75837 + smul_75838;
  assign add_76556 = smul_75839 + smul_75840;
  assign add_76557 = add_75841 + add_75842;
  assign add_76558 = smul_75843 + smul_75844;
  assign add_76559 = smul_75845 + smul_75846;
  assign add_76560 = smul_75847 + smul_75848;
  assign add_76561 = add_75849 + add_75850;
  assign add_76562 = smul_75851 + smul_75852;
  assign add_76563 = smul_75853 + smul_75854;
  assign add_76564 = smul_75855 + smul_75856;
  assign add_76565 = add_75857 + add_75858;
  assign add_76566 = smul_75859 + smul_75860;
  assign add_76567 = smul_75861 + smul_75862;
  assign add_76568 = smul_75863 + smul_75864;
  assign add_76569 = add_75865 + add_75866;
  assign add_76570 = smul_75867 + smul_75868;
  assign add_76571 = smul_75869 + smul_75870;
  assign add_76572 = smul_75871 + smul_75872;
  assign add_76573 = add_75873 + add_75874;
  assign add_76574 = smul_75875 + smul_75876;
  assign add_76575 = smul_75877 + smul_75878;
  assign add_76576 = smul_75879 + smul_75880;
  assign add_76577 = add_75881 + add_75882;
  assign add_76578 = smul_75883 + smul_75884;
  assign add_76579 = smul_75885 + smul_75886;
  assign add_76580 = smul_75887 + smul_75888;
  assign add_76581 = add_75889 + add_75890;
  assign add_76582 = smul_75891 + smul_75892;
  assign add_76583 = smul_75893 + smul_75894;
  assign add_76584 = smul_75895 + smul_75896;
  assign add_76585 = add_75897 + add_75898;
  assign add_76586 = smul_75899 + smul_75900;
  assign add_76587 = smul_75901 + smul_75902;
  assign add_76588 = smul_75903 + smul_75904;
  assign add_76589 = add_75905 + add_75906;
  assign add_76590 = smul_75907 + smul_75908;
  assign add_76591 = smul_75909 + smul_75910;
  assign add_76592 = smul_75911 + smul_75912;
  assign add_76593 = add_75913 + add_75914;
  assign add_76594 = smul_75915 + smul_75916;
  assign add_76595 = smul_75917 + smul_75918;
  assign add_76596 = smul_75919 + smul_75920;
  assign add_76597 = add_75921 + add_75922;
  assign add_76598 = smul_75923 + smul_75924;
  assign add_76599 = smul_75925 + smul_75926;
  assign add_76600 = smul_75927 + smul_75928;
  assign add_76601 = add_75929 + add_75930;
  assign add_76602 = smul_75931 + smul_75932;
  assign add_76603 = smul_75933 + smul_75934;
  assign add_76604 = smul_75935 + smul_75936;
  assign add_76605 = add_75937 + add_75938;
  assign add_76606 = smul_75939 + smul_75940;
  assign add_76607 = smul_75941 + smul_75942;
  assign add_76608 = smul_75943 + smul_75944;
  assign add_76609 = add_75945 + add_75946;
  assign add_76610 = smul_75947 + smul_75948;
  assign add_76611 = smul_75949 + smul_75950;
  assign add_76612 = smul_75951 + smul_75952;
  assign add_76613 = add_75953 + add_75954;
  assign add_76614 = smul_75955 + smul_75956;
  assign add_76615 = smul_75957 + smul_75958;
  assign add_76616 = smul_75959 + smul_75960;
  assign add_76617 = add_75961 + add_75962;
  assign add_76618 = smul_75963 + smul_75964;
  assign add_76619 = smul_75965 + smul_75966;
  assign add_76620 = smul_75967 + smul_75968;
  assign add_76621 = add_75969 + add_75970;
  assign add_76622 = smul_75971 + smul_75972;
  assign add_76623 = smul_75973 + smul_75974;
  assign add_76624 = smul_75975 + smul_75976;
  assign add_76625 = add_75977 + add_75978;
  assign add_76626 = smul_75979 + smul_75980;
  assign add_76627 = smul_75981 + smul_75982;
  assign add_76628 = smul_75983 + smul_75984;
  assign add_76629 = add_75985 + add_75986;
  assign add_76630 = smul_75987 + smul_75988;
  assign add_76631 = smul_75989 + smul_75990;
  assign add_76632 = smul_75991 + smul_75992;
  assign add_76633 = add_75993 + add_75994;
  assign add_76634 = smul_75995 + smul_75996;
  assign add_76635 = smul_75997 + smul_75998;
  assign add_76636 = smul_75999 + smul_76000;
  assign add_76637 = add_76001 + add_76002;
  assign add_76638 = smul_76003 + smul_76004;
  assign add_76639 = smul_76005 + smul_76006;
  assign add_76640 = smul_76007 + smul_76008;
  assign add_76641 = add_76009 + add_76010;
  assign add_76642 = smul_76011 + smul_76012;
  assign add_76643 = smul_76013 + smul_76014;
  assign add_76644 = smul_76015 + smul_76016;
  assign add_76645 = add_76017 + add_76018;
  assign add_76646 = smul_76019 + smul_76020;
  assign add_76647 = smul_76021 + smul_76022;
  assign add_76648 = smul_76023 + smul_76024;
  assign add_76649 = add_76025 + add_76026;
  assign add_76650 = smul_76027 + smul_76028;
  assign add_76651 = smul_76029 + smul_76030;
  assign add_76652 = smul_76031 + smul_76032;
  assign add_76653 = add_76033 + add_76034;
  assign add_76654 = smul_76035 + smul_76036;
  assign add_76655 = smul_76037 + smul_76038;
  assign add_76656 = smul_76039 + smul_76040;
  assign add_76657 = add_76041 + add_76042;
  assign add_76658 = smul_76043 + smul_76044;
  assign add_76659 = smul_76045 + smul_76046;
  assign add_76660 = smul_76047 + smul_76048;
  assign add_76661 = add_76049 + add_76050;
  assign add_76662 = smul_76051 + smul_76052;
  assign add_76663 = smul_76053 + smul_76054;
  assign add_76664 = smul_76055 + smul_76056;
  assign add_76665 = add_76057 + add_76058;
  assign add_76666 = smul_76059 + smul_76060;
  assign add_76667 = smul_76061 + smul_76062;
  assign add_76668 = smul_76063 + smul_76064;
  assign add_76669 = add_76065 + add_76066;
  assign add_76670 = smul_76067 + smul_76068;
  assign add_76671 = smul_76069 + smul_76070;
  assign add_76672 = smul_76071 + smul_76072;
  assign add_76673 = add_76073 + add_76074;
  assign add_76674 = smul_76075 + smul_76076;
  assign add_76675 = smul_76077 + smul_76078;
  assign add_76676 = smul_76079 + smul_76080;
  assign add_76677 = add_76081 + add_76082;
  assign add_76678 = smul_76083 + smul_76084;
  assign add_76679 = smul_76085 + smul_76086;
  assign add_76680 = smul_76087 + smul_76088;
  assign add_76681 = add_76089 + add_76090;
  assign add_76682 = smul_76091 + smul_76092;
  assign add_76683 = smul_76093 + smul_76094;
  assign add_76684 = smul_76095 + smul_76096;
  assign add_76685 = add_76097 + add_76098;
  assign add_76686 = smul_76099 + smul_76100;
  assign add_76687 = smul_76101 + smul_76102;
  assign add_76688 = smul_76103 + smul_76104;
  assign add_76689 = add_76105 + add_76106;
  assign add_76690 = smul_76107 + smul_76108;
  assign add_76691 = smul_76109 + smul_76110;
  assign add_76692 = smul_76111 + smul_76112;
  assign add_76693 = add_76113 + add_76114;
  assign add_76694 = smul_76115 + smul_76116;
  assign add_76695 = smul_76117 + smul_76118;
  assign add_76696 = smul_76119 + smul_76120;
  assign add_76697 = add_76121 + add_76122;
  assign add_76698 = smul_76123 + smul_76124;
  assign add_76699 = smul_76125 + smul_76126;
  assign add_76700 = smul_76127 + smul_76128;
  assign add_76701 = add_76129 + add_76130;
  assign add_76702 = smul_76131 + smul_76132;
  assign add_76703 = smul_76133 + smul_76134;
  assign add_76704 = smul_76135 + smul_76136;
  assign add_76705 = add_76137 + add_76138;
  assign add_76706 = smul_76139 + smul_76140;
  assign add_76707 = smul_76141 + smul_76142;
  assign add_76708 = smul_76143 + smul_76144;
  assign add_76709 = add_76145 + add_76146;
  assign add_76710 = smul_76147 + smul_76148;
  assign add_76711 = smul_76149 + smul_76150;
  assign add_76712 = smul_76151 + smul_76152;
  assign add_76713 = add_76153 + add_76154;
  assign add_76714 = smul_76155 + smul_76156;
  assign add_76715 = smul_76157 + smul_76158;
  assign add_76716 = smul_76159 + smul_76160;
  assign add_76717 = add_76161 + add_76162;
  assign add_76718 = smul_76163 + smul_76164;
  assign add_76719 = smul_76165 + smul_76166;
  assign add_76720 = smul_76167 + smul_76168;
  assign add_76721 = add_76169 + add_76170;
  assign add_76722 = smul_76171 + smul_76172;
  assign add_76723 = smul_76173 + smul_76174;
  assign add_76724 = smul_76175 + smul_76176;
  assign add_76725 = add_76177 + add_76178;
  assign add_76726 = smul_76179 + smul_76180;
  assign add_76727 = smul_76181 + smul_76182;
  assign add_76728 = smul_76183 + smul_76184;
  assign add_76729 = add_76185 + add_76186;
  assign add_76730 = smul_76187 + smul_76188;
  assign add_76731 = smul_76189 + smul_76190;
  assign add_76732 = smul_76191 + smul_76192;
  assign add_76733 = add_76193 + add_76194;
  assign add_76734 = smul_76195 + smul_76196;
  assign add_76735 = smul_76197 + smul_76198;
  assign add_76736 = smul_76199 + smul_76200;
  assign add_76737 = add_76201 + add_76202;
  assign add_76738 = smul_76203 + smul_76204;
  assign add_76739 = smul_76205 + smul_76206;
  assign add_76740 = smul_76207 + smul_76208;
  assign add_76741 = add_76209 + add_76210;
  assign add_76742 = smul_76211 + smul_76212;
  assign add_76743 = smul_76213 + smul_76214;
  assign add_76744 = smul_76215 + smul_76216;
  assign add_76745 = add_76217 + add_76218;
  assign add_76746 = smul_76219 + smul_76220;
  assign add_76747 = smul_76221 + smul_76222;
  assign add_76748 = smul_76223 + smul_76224;
  assign add_76749 = add_76225 + add_76226;
  assign add_76750 = smul_76227 + smul_76228;
  assign add_76751 = smul_76229 + smul_76230;
  assign add_76752 = smul_76231 + smul_76232;
  assign add_76753 = add_76233 + add_76234;
  assign add_76754 = smul_76235 + smul_76236;
  assign add_76755 = smul_76237 + smul_76238;
  assign add_76756 = smul_76239 + smul_76240;
  assign add_76757 = add_76241 + add_76242;
  assign add_76758 = smul_76243 + smul_76244;
  assign add_76759 = smul_76245 + smul_76246;
  assign add_76760 = smul_76247 + smul_76248;
  assign add_76761 = add_76249 + add_76250;
  assign add_76762 = smul_76251 + smul_76252;
  assign add_76763 = smul_76253 + smul_76254;
  assign add_76764 = smul_76255 + smul_76256;
  assign add_76765 = add_76257 + add_76258;
  assign add_76766 = smul_76259 + smul_76260;
  assign add_76767 = smul_76261 + smul_76262;
  assign add_76768 = smul_76263 + smul_76264;
  assign add_76769 = add_76265 + add_76266;
  assign add_76770 = smul_76267 + smul_76268;
  assign add_76771 = smul_76269 + smul_76270;
  assign add_76772 = smul_76271 + smul_76272;
  assign add_76773 = add_76273 + add_76274;
  assign add_76774 = smul_76275 + smul_76276;
  assign add_76775 = smul_76277 + smul_76278;
  assign add_76776 = smul_76279 + smul_76280;
  assign add_76777 = add_76281 + add_76282;
  assign add_76778 = smul_76283 + smul_76284;
  assign add_76779 = smul_76285 + smul_76286;
  assign add_76780 = smul_76287 + smul_76288;
  assign add_76781 = add_76289 + add_76290;
  assign add_76782 = smul_76291 + smul_76292;
  assign add_76783 = smul_76293 + smul_76294;
  assign add_76784 = smul_76295 + smul_76296;
  assign add_76785 = add_76297 + add_76298;
  assign add_76786 = smul_76299 + smul_76300;
  assign add_76787 = smul_76301 + smul_76302;
  assign add_76788 = smul_76303 + smul_76304;
  assign add_76789 = add_76305 + add_76306;
  assign add_76790 = smul_76307 + smul_76308;
  assign add_76791 = smul_76309 + smul_76310;
  assign add_76792 = smul_76311 + smul_76312;
  assign add_76793 = add_76313 + add_76314;
  assign add_76794 = smul_76315 + smul_76316;
  assign add_76795 = smul_76317 + smul_76318;
  assign add_76796 = smul_76319 + smul_76320;
  assign add_76797 = add_76321 + add_76322;
  assign add_76798 = smul_76323 + smul_76324;
  assign add_76799 = smul_76325 + smul_76326;
  assign add_76800 = smul_76327 + smul_76328;
  assign add_76801 = add_76329 + add_76330;
  assign add_76802 = smul_76331 + smul_76332;
  assign add_76803 = smul_76333 + smul_76334;
  assign add_76804 = smul_76335 + smul_76336;
  assign add_76805 = add_76337 + add_76338;
  assign add_76806 = smul_76339 + smul_76340;
  assign add_76807 = smul_76341 + smul_76342;
  assign add_76808 = smul_76343 + smul_76344;
  assign add_76809 = add_76345 + add_76346;
  assign add_76810 = smul_76347 + smul_76348;
  assign add_76811 = smul_76349 + smul_76350;
  assign add_76812 = smul_76351 + smul_76352;
  assign add_76813 = add_76353 + add_76354;
  assign add_76814 = smul_76355 + smul_76356;
  assign add_76815 = smul_76357 + smul_76358;
  assign add_76816 = smul_76359 + smul_76360;
  assign add_76817 = add_76361 + add_76362;
  assign add_76818 = smul_76363 + smul_76364;
  assign add_76819 = smul_76365 + smul_76366;
  assign add_76820 = smul_76367 + smul_76368;
  assign add_76821 = add_76369 + add_76370;
  assign add_76822 = smul_76371 + smul_76372;
  assign add_76823 = smul_76373 + smul_76374;
  assign add_76824 = smul_76375 + smul_76376;
  assign add_76825 = add_76377 + add_76378;
  assign add_76826 = smul_76379 + smul_76380;
  assign add_76827 = smul_76381 + smul_76382;
  assign add_76828 = smul_76383 + smul_76384;
  assign add_76829 = add_76385 + add_76386;
  assign add_76830 = smul_76387 + smul_76388;
  assign add_76831 = smul_76389 + smul_76390;
  assign add_76832 = smul_76391 + smul_76392;
  assign add_76833 = add_76393 + add_76394;
  assign add_76834 = smul_76395 + smul_76396;
  assign add_76835 = smul_76397 + smul_76398;
  assign add_76836 = smul_76399 + smul_76400;
  assign add_76837 = add_76401 + add_76402;
  assign add_76838 = smul_76403 + smul_76404;
  assign add_76839 = smul_76405 + smul_76406;
  assign add_76840 = smul_76407 + smul_76408;
  assign add_76841 = add_76409 + add_76410;
  assign add_76842 = smul_76411 + smul_76412;
  assign add_76843 = smul_76413 + smul_76414;
  assign add_76844 = smul_76415 + smul_76416;
  assign add_76845 = add_76417 + add_76418;
  assign add_76846 = smul_76419 + smul_76420;
  assign add_76847 = smul_76421 + smul_76422;
  assign add_76848 = smul_76423 + smul_76424;
  assign add_76849 = add_76425 + add_76426;
  assign add_76850 = smul_76427 + smul_76428;
  assign add_76851 = smul_76429 + smul_76430;
  assign add_76852 = smul_76431 + smul_76432;
  assign add_76853 = add_76433 + add_76434;
  assign add_76854 = smul_76435 + smul_76436;
  assign add_76855 = smul_76437 + smul_76438;
  assign add_76856 = smul_76439 + smul_76440;
  assign add_76857 = add_76441 + add_76442;
  assign add_76858 = smul_76443 + smul_76444;
  assign add_76859 = smul_76445 + smul_76446;
  assign add_76860 = smul_76447 + smul_76448;
  assign add_76861 = add_76449 + add_76450;
  assign add_76862 = smul_76451 + smul_76452;
  assign add_76863 = smul_76453 + smul_76454;
  assign add_76864 = smul_76455 + smul_76456;
  assign add_76865 = add_76457 + add_76458;
  assign add_76866 = smul_76459 + smul_76460;
  assign add_76867 = smul_76461 + smul_76462;
  assign add_76868 = smul_76463 + smul_76464;
  assign add_76869 = add_76465 + add_76466;
  assign add_76870 = smul_76467 + smul_76468;
  assign add_76871 = smul_76469 + smul_76470;
  assign add_76872 = smul_76471 + smul_76472;
  assign add_76873 = add_76473 + add_76474;
  assign add_76874 = add_76475 + add_76476;
  assign add_76875 = add_76477 + add_76478;
  assign add_76876 = add_76479 + add_76480;
  assign add_76877 = add_76481 + add_76482;
  assign add_76878 = add_76483 + add_76484;
  assign add_76879 = add_76485 + add_76486;
  assign add_76880 = add_76487 + add_76488;
  assign add_76881 = add_76489 + add_76490;
  assign add_76882 = add_76491 + add_76492;
  assign add_76883 = add_76493 + add_76494;
  assign add_76884 = add_76495 + add_76496;
  assign add_76885 = add_76497 + add_76498;
  assign add_76886 = add_76499 + add_76500;
  assign add_76887 = add_76501 + add_76502;
  assign add_76888 = add_76503 + add_76504;
  assign add_76889 = add_76505 + add_76506;
  assign add_76890 = add_76507 + add_76508;
  assign add_76891 = add_76509 + add_76510;
  assign add_76892 = add_76511 + add_76512;
  assign add_76893 = add_76513 + add_76514;
  assign add_76894 = add_76515 + add_76516;
  assign add_76895 = add_76517 + add_76518;
  assign add_76896 = add_76519 + add_76520;
  assign add_76897 = add_76521 + add_76522;
  assign add_76898 = add_76523 + add_76524;
  assign add_76899 = add_76525 + add_76526;
  assign add_76900 = add_76527 + add_76528;
  assign add_76901 = add_76529 + add_76530;
  assign add_76902 = add_76531 + add_76532;
  assign add_76903 = add_76533 + add_76534;
  assign add_76904 = add_76535 + add_76536;
  assign add_76905 = add_76537 + add_76538;
  assign add_76906 = add_76539 + add_76540;
  assign add_76907 = add_76541 + add_76542;
  assign add_76908 = add_76543 + add_76544;
  assign add_76909 = add_76545 + add_76546;
  assign add_76910 = add_76547 + add_76548;
  assign add_76911 = add_76549 + add_76550;
  assign add_76912 = add_76551 + add_76552;
  assign add_76913 = add_76553 + add_76554;
  assign add_76914 = add_76555 + add_76556;
  assign add_76915 = add_76557 + add_76558;
  assign add_76916 = add_76559 + add_76560;
  assign add_76917 = add_76561 + add_76562;
  assign add_76918 = add_76563 + add_76564;
  assign add_76919 = add_76565 + add_76566;
  assign add_76920 = add_76567 + add_76568;
  assign add_76921 = add_76569 + add_76570;
  assign add_76922 = add_76571 + add_76572;
  assign add_76923 = add_76573 + add_76574;
  assign add_76924 = add_76575 + add_76576;
  assign add_76925 = add_76577 + add_76578;
  assign add_76926 = add_76579 + add_76580;
  assign add_76927 = add_76581 + add_76582;
  assign add_76928 = add_76583 + add_76584;
  assign add_76929 = add_76585 + add_76586;
  assign add_76930 = add_76587 + add_76588;
  assign add_76931 = add_76589 + add_76590;
  assign add_76932 = add_76591 + add_76592;
  assign add_76933 = add_76593 + add_76594;
  assign add_76934 = add_76595 + add_76596;
  assign add_76935 = add_76597 + add_76598;
  assign add_76936 = add_76599 + add_76600;
  assign add_76937 = add_76601 + add_76602;
  assign add_76938 = add_76603 + add_76604;
  assign add_76939 = add_76605 + add_76606;
  assign add_76940 = add_76607 + add_76608;
  assign add_76941 = add_76609 + add_76610;
  assign add_76942 = add_76611 + add_76612;
  assign add_76943 = add_76613 + add_76614;
  assign add_76944 = add_76615 + add_76616;
  assign add_76945 = add_76617 + add_76618;
  assign add_76946 = add_76619 + add_76620;
  assign add_76947 = add_76621 + add_76622;
  assign add_76948 = add_76623 + add_76624;
  assign add_76949 = add_76625 + add_76626;
  assign add_76950 = add_76627 + add_76628;
  assign add_76951 = add_76629 + add_76630;
  assign add_76952 = add_76631 + add_76632;
  assign add_76953 = add_76633 + add_76634;
  assign add_76954 = add_76635 + add_76636;
  assign add_76955 = add_76637 + add_76638;
  assign add_76956 = add_76639 + add_76640;
  assign add_76957 = add_76641 + add_76642;
  assign add_76958 = add_76643 + add_76644;
  assign add_76959 = add_76645 + add_76646;
  assign add_76960 = add_76647 + add_76648;
  assign add_76961 = add_76649 + add_76650;
  assign add_76962 = add_76651 + add_76652;
  assign add_76963 = add_76653 + add_76654;
  assign add_76964 = add_76655 + add_76656;
  assign add_76965 = add_76657 + add_76658;
  assign add_76966 = add_76659 + add_76660;
  assign add_76967 = add_76661 + add_76662;
  assign add_76968 = add_76663 + add_76664;
  assign add_76969 = add_76665 + add_76666;
  assign add_76970 = add_76667 + add_76668;
  assign add_76971 = add_76669 + add_76670;
  assign add_76972 = add_76671 + add_76672;
  assign add_76973 = add_76673 + add_76674;
  assign add_76974 = add_76675 + add_76676;
  assign add_76975 = add_76677 + add_76678;
  assign add_76976 = add_76679 + add_76680;
  assign add_76977 = add_76681 + add_76682;
  assign add_76978 = add_76683 + add_76684;
  assign add_76979 = add_76685 + add_76686;
  assign add_76980 = add_76687 + add_76688;
  assign add_76981 = add_76689 + add_76690;
  assign add_76982 = add_76691 + add_76692;
  assign add_76983 = add_76693 + add_76694;
  assign add_76984 = add_76695 + add_76696;
  assign add_76985 = add_76697 + add_76698;
  assign add_76986 = add_76699 + add_76700;
  assign add_76987 = add_76701 + add_76702;
  assign add_76988 = add_76703 + add_76704;
  assign add_76989 = add_76705 + add_76706;
  assign add_76990 = add_76707 + add_76708;
  assign add_76991 = add_76709 + add_76710;
  assign add_76992 = add_76711 + add_76712;
  assign add_76993 = add_76713 + add_76714;
  assign add_76994 = add_76715 + add_76716;
  assign add_76995 = add_76717 + add_76718;
  assign add_76996 = add_76719 + add_76720;
  assign add_76997 = add_76721 + add_76722;
  assign add_76998 = add_76723 + add_76724;
  assign add_76999 = add_76725 + add_76726;
  assign add_77000 = add_76727 + add_76728;
  assign add_77001 = add_76729 + add_76730;
  assign add_77002 = add_76731 + add_76732;
  assign add_77003 = add_76733 + add_76734;
  assign add_77004 = add_76735 + add_76736;
  assign add_77005 = add_76737 + add_76738;
  assign add_77006 = add_76739 + add_76740;
  assign add_77007 = add_76741 + add_76742;
  assign add_77008 = add_76743 + add_76744;
  assign add_77009 = add_76745 + add_76746;
  assign add_77010 = add_76747 + add_76748;
  assign add_77011 = add_76749 + add_76750;
  assign add_77012 = add_76751 + add_76752;
  assign add_77013 = add_76753 + add_76754;
  assign add_77014 = add_76755 + add_76756;
  assign add_77015 = add_76757 + add_76758;
  assign add_77016 = add_76759 + add_76760;
  assign add_77017 = add_76761 + add_76762;
  assign add_77018 = add_76763 + add_76764;
  assign add_77019 = add_76765 + add_76766;
  assign add_77020 = add_76767 + add_76768;
  assign add_77021 = add_76769 + add_76770;
  assign add_77022 = add_76771 + add_76772;
  assign add_77023 = add_76773 + add_76774;
  assign add_77024 = add_76775 + add_76776;
  assign add_77025 = add_76777 + add_76778;
  assign add_77026 = add_76779 + add_76780;
  assign add_77027 = add_76781 + add_76782;
  assign add_77028 = add_76783 + add_76784;
  assign add_77029 = add_76785 + add_76786;
  assign add_77030 = add_76787 + add_76788;
  assign add_77031 = add_76789 + add_76790;
  assign add_77032 = add_76791 + add_76792;
  assign add_77033 = add_76793 + add_76794;
  assign add_77034 = add_76795 + add_76796;
  assign add_77035 = add_76797 + add_76798;
  assign add_77036 = add_76799 + add_76800;
  assign add_77037 = add_76801 + add_76802;
  assign add_77038 = add_76803 + add_76804;
  assign add_77039 = add_76805 + add_76806;
  assign add_77040 = add_76807 + add_76808;
  assign add_77041 = add_76809 + add_76810;
  assign add_77042 = add_76811 + add_76812;
  assign add_77043 = add_76813 + add_76814;
  assign add_77044 = add_76815 + add_76816;
  assign add_77045 = add_76817 + add_76818;
  assign add_77046 = add_76819 + add_76820;
  assign add_77047 = add_76821 + add_76822;
  assign add_77048 = add_76823 + add_76824;
  assign add_77049 = add_76825 + add_76826;
  assign add_77050 = add_76827 + add_76828;
  assign add_77051 = add_76829 + add_76830;
  assign add_77052 = add_76831 + add_76832;
  assign add_77053 = add_76833 + add_76834;
  assign add_77054 = add_76835 + add_76836;
  assign add_77055 = add_76837 + add_76838;
  assign add_77056 = add_76839 + add_76840;
  assign add_77057 = add_76841 + add_76842;
  assign add_77058 = add_76843 + add_76844;
  assign add_77059 = add_76845 + add_76846;
  assign add_77060 = add_76847 + add_76848;
  assign add_77061 = add_76849 + add_76850;
  assign add_77062 = add_76851 + add_76852;
  assign add_77063 = add_76853 + add_76854;
  assign add_77064 = add_76855 + add_76856;
  assign add_77065 = add_76857 + add_76858;
  assign add_77066 = add_76859 + add_76860;
  assign add_77067 = add_76861 + add_76862;
  assign add_77068 = add_76863 + add_76864;
  assign add_77069 = add_76865 + add_76866;
  assign add_77070 = add_76867 + add_76868;
  assign add_77071 = add_76869 + add_76870;
  assign add_77072 = add_76871 + add_76872;
  assign add_77073 = add_76873 + add_76874;
  assign literal_77074 = 1'h1;
  assign add_77075 = add_76875 + add_76876;
  assign add_77076 = add_76877 + add_76878;
  assign add_77077 = add_76879 + add_76880;
  assign add_77078 = add_76881 + add_76882;
  assign add_77079 = add_76883 + add_76884;
  assign add_77080 = add_76885 + add_76886;
  assign add_77081 = add_76887 + add_76888;
  assign add_77082 = add_76889 + add_76890;
  assign add_77083 = add_76891 + add_76892;
  assign add_77084 = add_76893 + add_76894;
  assign add_77085 = add_76895 + add_76896;
  assign add_77086 = add_76897 + add_76898;
  assign add_77087 = add_76899 + add_76900;
  assign add_77088 = add_76901 + add_76902;
  assign add_77089 = add_76903 + add_76904;
  assign add_77090 = add_76905 + add_76906;
  assign add_77091 = add_76907 + add_76908;
  assign add_77092 = add_76909 + add_76910;
  assign add_77093 = add_76911 + add_76912;
  assign add_77094 = add_76913 + add_76914;
  assign add_77095 = add_76915 + add_76916;
  assign add_77096 = add_76917 + add_76918;
  assign add_77097 = add_76919 + add_76920;
  assign add_77098 = add_76921 + add_76922;
  assign add_77099 = add_76923 + add_76924;
  assign add_77100 = add_76925 + add_76926;
  assign add_77101 = add_76927 + add_76928;
  assign add_77102 = add_76929 + add_76930;
  assign add_77103 = add_76931 + add_76932;
  assign add_77104 = add_76933 + add_76934;
  assign add_77105 = add_76935 + add_76936;
  assign add_77106 = add_76937 + add_76938;
  assign add_77107 = add_76939 + add_76940;
  assign add_77108 = add_76941 + add_76942;
  assign add_77109 = add_76943 + add_76944;
  assign add_77110 = add_76945 + add_76946;
  assign add_77111 = add_76947 + add_76948;
  assign add_77112 = add_76949 + add_76950;
  assign add_77113 = add_76951 + add_76952;
  assign add_77114 = add_76953 + add_76954;
  assign add_77115 = add_76955 + add_76956;
  assign add_77116 = add_76957 + add_76958;
  assign add_77117 = add_76959 + add_76960;
  assign add_77118 = add_76961 + add_76962;
  assign add_77119 = add_76963 + add_76964;
  assign add_77120 = add_76965 + add_76966;
  assign add_77121 = add_76967 + add_76968;
  assign add_77122 = add_76969 + add_76970;
  assign add_77123 = add_76971 + add_76972;
  assign add_77124 = add_76973 + add_76974;
  assign add_77125 = add_76975 + add_76976;
  assign add_77126 = add_76977 + add_76978;
  assign add_77127 = add_76979 + add_76980;
  assign add_77128 = add_76981 + add_76982;
  assign add_77129 = add_76983 + add_76984;
  assign add_77130 = add_76985 + add_76986;
  assign add_77131 = add_76987 + add_76988;
  assign add_77132 = add_76989 + add_76990;
  assign add_77133 = add_76991 + add_76992;
  assign add_77134 = add_76993 + add_76994;
  assign add_77135 = add_76995 + add_76996;
  assign add_77136 = add_76997 + add_76998;
  assign add_77137 = add_76999 + add_77000;
  assign add_77138 = add_77001 + add_77002;
  assign add_77139 = add_77003 + add_77004;
  assign add_77140 = add_77005 + add_77006;
  assign add_77141 = add_77007 + add_77008;
  assign add_77142 = add_77009 + add_77010;
  assign add_77143 = add_77011 + add_77012;
  assign add_77144 = add_77013 + add_77014;
  assign add_77145 = add_77015 + add_77016;
  assign add_77146 = add_77017 + add_77018;
  assign add_77147 = add_77019 + add_77020;
  assign add_77148 = add_77021 + add_77022;
  assign add_77149 = add_77023 + add_77024;
  assign add_77150 = add_77025 + add_77026;
  assign add_77151 = add_77027 + add_77028;
  assign add_77152 = add_77029 + add_77030;
  assign add_77153 = add_77031 + add_77032;
  assign add_77154 = add_77033 + add_77034;
  assign add_77155 = add_77035 + add_77036;
  assign add_77156 = add_77037 + add_77038;
  assign add_77157 = add_77039 + add_77040;
  assign add_77158 = add_77041 + add_77042;
  assign add_77159 = add_77043 + add_77044;
  assign add_77160 = add_77045 + add_77046;
  assign add_77161 = add_77047 + add_77048;
  assign add_77162 = add_77049 + add_77050;
  assign add_77163 = add_77051 + add_77052;
  assign add_77164 = add_77053 + add_77054;
  assign add_77165 = add_77055 + add_77056;
  assign add_77166 = add_77057 + add_77058;
  assign add_77167 = add_77059 + add_77060;
  assign add_77168 = add_77061 + add_77062;
  assign add_77169 = add_77063 + add_77064;
  assign add_77170 = add_77065 + add_77066;
  assign add_77171 = add_77067 + add_77068;
  assign add_77172 = add_77069 + add_77070;
  assign add_77173 = add_77071 + add_77072;
  assign out = {literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, literal_77074, {add_77073, literal_77074}, {add_77075, literal_77074}, {add_77076, literal_77074}, {add_77077, literal_77074}, {add_77078, literal_77074}, {add_77079, literal_77074}, {add_77080, literal_77074}, {add_77081, literal_77074}, {add_77082, literal_77074}, {add_77083, literal_77074}, {add_77084, literal_77074}, {add_77085, literal_77074}, {add_77086, literal_77074}, {add_77087, literal_77074}, {add_77088, literal_77074}, {add_77089, literal_77074}, {add_77090, literal_77074}, {add_77091, literal_77074}, {add_77092, literal_77074}, {add_77093, literal_77074}, {add_77094, literal_77074}, {add_77095, literal_77074}, {add_77096, literal_77074}, {add_77097, literal_77074}, {add_77098, literal_77074}, {add_77099, literal_77074}, {add_77100, literal_77074}, {add_77101, literal_77074}, {add_77102, literal_77074}, {add_77103, literal_77074}, {add_77104, literal_77074}, {add_77105, literal_77074}, {add_77106, literal_77074}, {add_77107, literal_77074}, {add_77108, literal_77074}, {add_77109, literal_77074}, {add_77110, literal_77074}, {add_77111, literal_77074}, {add_77112, literal_77074}, {add_77113, literal_77074}, {add_77114, literal_77074}, {add_77115, literal_77074}, {add_77116, literal_77074}, {add_77117, literal_77074}, {add_77118, literal_77074}, {add_77119, literal_77074}, {add_77120, literal_77074}, {add_77121, literal_77074}, {add_77122, literal_77074}, {add_77123, literal_77074}, {add_77124, literal_77074}, {add_77125, literal_77074}, {add_77126, literal_77074}, {add_77127, literal_77074}, {add_77128, literal_77074}, {add_77129, literal_77074}, {add_77130, literal_77074}, {add_77131, literal_77074}, {add_77132, literal_77074}, {add_77133, literal_77074}, {add_77134, literal_77074}, {add_77135, literal_77074}, {add_77136, literal_77074}, {add_77137, literal_77074}, {add_77138, literal_77074}, {add_77139, literal_77074}, {add_77140, literal_77074}, {add_77141, literal_77074}, {add_77142, literal_77074}, {add_77143, literal_77074}, {add_77144, literal_77074}, {add_77145, literal_77074}, {add_77146, literal_77074}, {add_77147, literal_77074}, {add_77148, literal_77074}, {add_77149, literal_77074}, {add_77150, literal_77074}, {add_77151, literal_77074}, {add_77152, literal_77074}, {add_77153, literal_77074}, {add_77154, literal_77074}, {add_77155, literal_77074}, {add_77156, literal_77074}, {add_77157, literal_77074}, {add_77158, literal_77074}, {add_77159, literal_77074}, {add_77160, literal_77074}, {add_77161, literal_77074}, {add_77162, literal_77074}, {add_77163, literal_77074}, {add_77164, literal_77074}, {add_77165, literal_77074}, {add_77166, literal_77074}, {add_77167, literal_77074}, {add_77168, literal_77074}, {add_77169, literal_77074}, {add_77170, literal_77074}, {add_77171, literal_77074}, {add_77172, literal_77074}, {add_77173, literal_77074}};
endmodule
